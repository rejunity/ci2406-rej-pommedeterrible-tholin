magic
tech sky130B
magscale 1 2
timestamp 1717680035
<< obsli1 >>
rect 1104 2159 438840 157777
<< obsm1 >>
rect 1104 76 439378 159724
<< metal2 >>
rect 8390 159200 8446 160000
rect 9402 159200 9458 160000
rect 10414 159200 10470 160000
rect 11426 159200 11482 160000
rect 12438 159200 12494 160000
rect 13450 159200 13506 160000
rect 14462 159200 14518 160000
rect 15474 159200 15530 160000
rect 16486 159200 16542 160000
rect 17498 159200 17554 160000
rect 18510 159200 18566 160000
rect 19522 159200 19578 160000
rect 20534 159200 20590 160000
rect 21546 159200 21602 160000
rect 22558 159200 22614 160000
rect 23570 159200 23626 160000
rect 24582 159200 24638 160000
rect 25594 159200 25650 160000
rect 26606 159200 26662 160000
rect 27618 159200 27674 160000
rect 28630 159200 28686 160000
rect 29642 159200 29698 160000
rect 30654 159200 30710 160000
rect 31666 159200 31722 160000
rect 32678 159200 32734 160000
rect 33690 159200 33746 160000
rect 34702 159200 34758 160000
rect 35714 159200 35770 160000
rect 36726 159200 36782 160000
rect 37738 159200 37794 160000
rect 38750 159200 38806 160000
rect 39762 159200 39818 160000
rect 40774 159200 40830 160000
rect 41786 159200 41842 160000
rect 42798 159200 42854 160000
rect 43810 159200 43866 160000
rect 44822 159200 44878 160000
rect 45834 159200 45890 160000
rect 46846 159200 46902 160000
rect 47858 159200 47914 160000
rect 48870 159200 48926 160000
rect 49882 159200 49938 160000
rect 50894 159200 50950 160000
rect 51906 159200 51962 160000
rect 52918 159200 52974 160000
rect 53930 159200 53986 160000
rect 54942 159200 54998 160000
rect 55954 159200 56010 160000
rect 56966 159200 57022 160000
rect 57978 159200 58034 160000
rect 58990 159200 59046 160000
rect 60002 159200 60058 160000
rect 61014 159200 61070 160000
rect 62026 159200 62082 160000
rect 63038 159200 63094 160000
rect 64050 159200 64106 160000
rect 65062 159200 65118 160000
rect 66074 159200 66130 160000
rect 67086 159200 67142 160000
rect 68098 159200 68154 160000
rect 69110 159200 69166 160000
rect 70122 159200 70178 160000
rect 71134 159200 71190 160000
rect 72146 159200 72202 160000
rect 73158 159200 73214 160000
rect 74170 159200 74226 160000
rect 75182 159200 75238 160000
rect 76194 159200 76250 160000
rect 77206 159200 77262 160000
rect 78218 159200 78274 160000
rect 79230 159200 79286 160000
rect 80242 159200 80298 160000
rect 81254 159200 81310 160000
rect 82266 159200 82322 160000
rect 83278 159200 83334 160000
rect 84290 159200 84346 160000
rect 85302 159200 85358 160000
rect 86314 159200 86370 160000
rect 87326 159200 87382 160000
rect 88338 159200 88394 160000
rect 89350 159200 89406 160000
rect 90362 159200 90418 160000
rect 91374 159200 91430 160000
rect 92386 159200 92442 160000
rect 93398 159200 93454 160000
rect 94410 159200 94466 160000
rect 95422 159200 95478 160000
rect 96434 159200 96490 160000
rect 97446 159200 97502 160000
rect 98458 159200 98514 160000
rect 99470 159200 99526 160000
rect 100482 159200 100538 160000
rect 101494 159200 101550 160000
rect 102506 159200 102562 160000
rect 103518 159200 103574 160000
rect 104530 159200 104586 160000
rect 105542 159200 105598 160000
rect 106554 159200 106610 160000
rect 107566 159200 107622 160000
rect 108578 159200 108634 160000
rect 109590 159200 109646 160000
rect 110602 159200 110658 160000
rect 111614 159200 111670 160000
rect 112626 159200 112682 160000
rect 113638 159200 113694 160000
rect 114650 159200 114706 160000
rect 115662 159200 115718 160000
rect 116674 159200 116730 160000
rect 117686 159200 117742 160000
rect 118698 159200 118754 160000
rect 119710 159200 119766 160000
rect 120722 159200 120778 160000
rect 121734 159200 121790 160000
rect 122746 159200 122802 160000
rect 123758 159200 123814 160000
rect 124770 159200 124826 160000
rect 125782 159200 125838 160000
rect 126794 159200 126850 160000
rect 127806 159200 127862 160000
rect 128818 159200 128874 160000
rect 129830 159200 129886 160000
rect 130842 159200 130898 160000
rect 131854 159200 131910 160000
rect 132866 159200 132922 160000
rect 133878 159200 133934 160000
rect 134890 159200 134946 160000
rect 135902 159200 135958 160000
rect 136914 159200 136970 160000
rect 137926 159200 137982 160000
rect 138938 159200 138994 160000
rect 139950 159200 140006 160000
rect 140962 159200 141018 160000
rect 141974 159200 142030 160000
rect 142986 159200 143042 160000
rect 143998 159200 144054 160000
rect 145010 159200 145066 160000
rect 146022 159200 146078 160000
rect 147034 159200 147090 160000
rect 148046 159200 148102 160000
rect 149058 159200 149114 160000
rect 150070 159200 150126 160000
rect 151082 159200 151138 160000
rect 152094 159200 152150 160000
rect 153106 159200 153162 160000
rect 154118 159200 154174 160000
rect 155130 159200 155186 160000
rect 156142 159200 156198 160000
rect 157154 159200 157210 160000
rect 158166 159200 158222 160000
rect 159178 159200 159234 160000
rect 160190 159200 160246 160000
rect 161202 159200 161258 160000
rect 162214 159200 162270 160000
rect 163226 159200 163282 160000
rect 164238 159200 164294 160000
rect 165250 159200 165306 160000
rect 166262 159200 166318 160000
rect 167274 159200 167330 160000
rect 168286 159200 168342 160000
rect 169298 159200 169354 160000
rect 170310 159200 170366 160000
rect 171322 159200 171378 160000
rect 172334 159200 172390 160000
rect 173346 159200 173402 160000
rect 174358 159200 174414 160000
rect 175370 159200 175426 160000
rect 176382 159200 176438 160000
rect 177394 159200 177450 160000
rect 178406 159200 178462 160000
rect 179418 159200 179474 160000
rect 180430 159200 180486 160000
rect 181442 159200 181498 160000
rect 182454 159200 182510 160000
rect 183466 159200 183522 160000
rect 184478 159200 184534 160000
rect 185490 159200 185546 160000
rect 186502 159200 186558 160000
rect 187514 159200 187570 160000
rect 188526 159200 188582 160000
rect 189538 159200 189594 160000
rect 190550 159200 190606 160000
rect 191562 159200 191618 160000
rect 192574 159200 192630 160000
rect 193586 159200 193642 160000
rect 194598 159200 194654 160000
rect 195610 159200 195666 160000
rect 196622 159200 196678 160000
rect 197634 159200 197690 160000
rect 198646 159200 198702 160000
rect 199658 159200 199714 160000
rect 200670 159200 200726 160000
rect 201682 159200 201738 160000
rect 202694 159200 202750 160000
rect 203706 159200 203762 160000
rect 204718 159200 204774 160000
rect 205730 159200 205786 160000
rect 206742 159200 206798 160000
rect 207754 159200 207810 160000
rect 208766 159200 208822 160000
rect 209778 159200 209834 160000
rect 210790 159200 210846 160000
rect 211802 159200 211858 160000
rect 212814 159200 212870 160000
rect 213826 159200 213882 160000
rect 214838 159200 214894 160000
rect 215850 159200 215906 160000
rect 216862 159200 216918 160000
rect 217874 159200 217930 160000
rect 218886 159200 218942 160000
rect 219898 159200 219954 160000
rect 220910 159200 220966 160000
rect 221922 159200 221978 160000
rect 222934 159200 222990 160000
rect 223946 159200 224002 160000
rect 224958 159200 225014 160000
rect 225970 159200 226026 160000
rect 226982 159200 227038 160000
rect 227994 159200 228050 160000
rect 229006 159200 229062 160000
rect 230018 159200 230074 160000
rect 231030 159200 231086 160000
rect 232042 159200 232098 160000
rect 233054 159200 233110 160000
rect 234066 159200 234122 160000
rect 235078 159200 235134 160000
rect 236090 159200 236146 160000
rect 237102 159200 237158 160000
rect 238114 159200 238170 160000
rect 239126 159200 239182 160000
rect 240138 159200 240194 160000
rect 241150 159200 241206 160000
rect 242162 159200 242218 160000
rect 243174 159200 243230 160000
rect 244186 159200 244242 160000
rect 245198 159200 245254 160000
rect 246210 159200 246266 160000
rect 247222 159200 247278 160000
rect 248234 159200 248290 160000
rect 249246 159200 249302 160000
rect 250258 159200 250314 160000
rect 251270 159200 251326 160000
rect 252282 159200 252338 160000
rect 253294 159200 253350 160000
rect 254306 159200 254362 160000
rect 255318 159200 255374 160000
rect 256330 159200 256386 160000
rect 257342 159200 257398 160000
rect 258354 159200 258410 160000
rect 259366 159200 259422 160000
rect 260378 159200 260434 160000
rect 261390 159200 261446 160000
rect 262402 159200 262458 160000
rect 263414 159200 263470 160000
rect 264426 159200 264482 160000
rect 265438 159200 265494 160000
rect 266450 159200 266506 160000
rect 267462 159200 267518 160000
rect 268474 159200 268530 160000
rect 269486 159200 269542 160000
rect 270498 159200 270554 160000
rect 271510 159200 271566 160000
rect 272522 159200 272578 160000
rect 273534 159200 273590 160000
rect 274546 159200 274602 160000
rect 275558 159200 275614 160000
rect 276570 159200 276626 160000
rect 277582 159200 277638 160000
rect 278594 159200 278650 160000
rect 279606 159200 279662 160000
rect 280618 159200 280674 160000
rect 281630 159200 281686 160000
rect 282642 159200 282698 160000
rect 283654 159200 283710 160000
rect 284666 159200 284722 160000
rect 285678 159200 285734 160000
rect 286690 159200 286746 160000
rect 287702 159200 287758 160000
rect 288714 159200 288770 160000
rect 289726 159200 289782 160000
rect 290738 159200 290794 160000
rect 291750 159200 291806 160000
rect 292762 159200 292818 160000
rect 293774 159200 293830 160000
rect 294786 159200 294842 160000
rect 295798 159200 295854 160000
rect 296810 159200 296866 160000
rect 297822 159200 297878 160000
rect 298834 159200 298890 160000
rect 299846 159200 299902 160000
rect 300858 159200 300914 160000
rect 301870 159200 301926 160000
rect 302882 159200 302938 160000
rect 303894 159200 303950 160000
rect 304906 159200 304962 160000
rect 305918 159200 305974 160000
rect 306930 159200 306986 160000
rect 307942 159200 307998 160000
rect 308954 159200 309010 160000
rect 309966 159200 310022 160000
rect 310978 159200 311034 160000
rect 311990 159200 312046 160000
rect 313002 159200 313058 160000
rect 314014 159200 314070 160000
rect 315026 159200 315082 160000
rect 316038 159200 316094 160000
rect 317050 159200 317106 160000
rect 318062 159200 318118 160000
rect 319074 159200 319130 160000
rect 320086 159200 320142 160000
rect 321098 159200 321154 160000
rect 322110 159200 322166 160000
rect 323122 159200 323178 160000
rect 324134 159200 324190 160000
rect 325146 159200 325202 160000
rect 326158 159200 326214 160000
rect 327170 159200 327226 160000
rect 328182 159200 328238 160000
rect 329194 159200 329250 160000
rect 330206 159200 330262 160000
rect 331218 159200 331274 160000
rect 332230 159200 332286 160000
rect 333242 159200 333298 160000
rect 334254 159200 334310 160000
rect 335266 159200 335322 160000
rect 336278 159200 336334 160000
rect 337290 159200 337346 160000
rect 338302 159200 338358 160000
rect 339314 159200 339370 160000
rect 340326 159200 340382 160000
rect 341338 159200 341394 160000
rect 342350 159200 342406 160000
rect 343362 159200 343418 160000
rect 344374 159200 344430 160000
rect 345386 159200 345442 160000
rect 346398 159200 346454 160000
rect 347410 159200 347466 160000
rect 348422 159200 348478 160000
rect 349434 159200 349490 160000
rect 350446 159200 350502 160000
rect 351458 159200 351514 160000
rect 352470 159200 352526 160000
rect 353482 159200 353538 160000
rect 354494 159200 354550 160000
rect 355506 159200 355562 160000
rect 356518 159200 356574 160000
rect 357530 159200 357586 160000
rect 358542 159200 358598 160000
rect 359554 159200 359610 160000
rect 360566 159200 360622 160000
rect 361578 159200 361634 160000
rect 362590 159200 362646 160000
rect 363602 159200 363658 160000
rect 364614 159200 364670 160000
rect 365626 159200 365682 160000
rect 366638 159200 366694 160000
rect 367650 159200 367706 160000
rect 368662 159200 368718 160000
rect 369674 159200 369730 160000
rect 370686 159200 370742 160000
rect 371698 159200 371754 160000
rect 372710 159200 372766 160000
rect 373722 159200 373778 160000
rect 374734 159200 374790 160000
rect 375746 159200 375802 160000
rect 376758 159200 376814 160000
rect 377770 159200 377826 160000
rect 378782 159200 378838 160000
rect 379794 159200 379850 160000
rect 380806 159200 380862 160000
rect 381818 159200 381874 160000
rect 382830 159200 382886 160000
rect 383842 159200 383898 160000
rect 384854 159200 384910 160000
rect 385866 159200 385922 160000
rect 386878 159200 386934 160000
rect 387890 159200 387946 160000
rect 388902 159200 388958 160000
rect 389914 159200 389970 160000
rect 390926 159200 390982 160000
rect 391938 159200 391994 160000
rect 392950 159200 393006 160000
rect 393962 159200 394018 160000
rect 394974 159200 395030 160000
rect 395986 159200 396042 160000
rect 396998 159200 397054 160000
rect 398010 159200 398066 160000
rect 399022 159200 399078 160000
rect 400034 159200 400090 160000
rect 401046 159200 401102 160000
rect 402058 159200 402114 160000
rect 403070 159200 403126 160000
rect 404082 159200 404138 160000
rect 405094 159200 405150 160000
rect 406106 159200 406162 160000
rect 407118 159200 407174 160000
rect 408130 159200 408186 160000
rect 409142 159200 409198 160000
rect 410154 159200 410210 160000
rect 411166 159200 411222 160000
rect 412178 159200 412234 160000
rect 413190 159200 413246 160000
rect 414202 159200 414258 160000
rect 415214 159200 415270 160000
rect 416226 159200 416282 160000
rect 417238 159200 417294 160000
rect 418250 159200 418306 160000
rect 419262 159200 419318 160000
rect 420274 159200 420330 160000
rect 421286 159200 421342 160000
rect 422298 159200 422354 160000
rect 423310 159200 423366 160000
rect 424322 159200 424378 160000
rect 425334 159200 425390 160000
rect 426346 159200 426402 160000
rect 427358 159200 427414 160000
rect 428370 159200 428426 160000
rect 429382 159200 429438 160000
rect 430394 159200 430450 160000
rect 431406 159200 431462 160000
rect 8390 0 8446 800
rect 10138 0 10194 800
rect 11886 0 11942 800
rect 13634 0 13690 800
rect 15382 0 15438 800
rect 17130 0 17186 800
rect 18878 0 18934 800
rect 20626 0 20682 800
rect 22374 0 22430 800
rect 24122 0 24178 800
rect 25870 0 25926 800
rect 27618 0 27674 800
rect 29366 0 29422 800
rect 31114 0 31170 800
rect 32862 0 32918 800
rect 34610 0 34666 800
rect 36358 0 36414 800
rect 38106 0 38162 800
rect 39854 0 39910 800
rect 41602 0 41658 800
rect 43350 0 43406 800
rect 45098 0 45154 800
rect 46846 0 46902 800
rect 48594 0 48650 800
rect 50342 0 50398 800
rect 52090 0 52146 800
rect 53838 0 53894 800
rect 55586 0 55642 800
rect 57334 0 57390 800
rect 59082 0 59138 800
rect 60830 0 60886 800
rect 62578 0 62634 800
rect 64326 0 64382 800
rect 66074 0 66130 800
rect 67822 0 67878 800
rect 69570 0 69626 800
rect 71318 0 71374 800
rect 73066 0 73122 800
rect 74814 0 74870 800
rect 76562 0 76618 800
rect 78310 0 78366 800
rect 80058 0 80114 800
rect 81806 0 81862 800
rect 83554 0 83610 800
rect 85302 0 85358 800
rect 87050 0 87106 800
rect 88798 0 88854 800
rect 90546 0 90602 800
rect 92294 0 92350 800
rect 94042 0 94098 800
rect 95790 0 95846 800
rect 97538 0 97594 800
rect 99286 0 99342 800
rect 101034 0 101090 800
rect 102782 0 102838 800
rect 104530 0 104586 800
rect 106278 0 106334 800
rect 108026 0 108082 800
rect 109774 0 109830 800
rect 111522 0 111578 800
rect 113270 0 113326 800
rect 115018 0 115074 800
rect 116766 0 116822 800
rect 118514 0 118570 800
rect 120262 0 120318 800
rect 122010 0 122066 800
rect 123758 0 123814 800
rect 125506 0 125562 800
rect 127254 0 127310 800
rect 129002 0 129058 800
rect 130750 0 130806 800
rect 132498 0 132554 800
rect 134246 0 134302 800
rect 135994 0 136050 800
rect 137742 0 137798 800
rect 139490 0 139546 800
rect 141238 0 141294 800
rect 142986 0 143042 800
rect 144734 0 144790 800
rect 146482 0 146538 800
rect 148230 0 148286 800
rect 149978 0 150034 800
rect 151726 0 151782 800
rect 153474 0 153530 800
rect 155222 0 155278 800
rect 156970 0 157026 800
rect 158718 0 158774 800
rect 160466 0 160522 800
rect 162214 0 162270 800
rect 163962 0 164018 800
rect 165710 0 165766 800
rect 167458 0 167514 800
rect 169206 0 169262 800
rect 170954 0 171010 800
rect 172702 0 172758 800
rect 174450 0 174506 800
rect 176198 0 176254 800
rect 177946 0 178002 800
rect 179694 0 179750 800
rect 181442 0 181498 800
rect 183190 0 183246 800
rect 184938 0 184994 800
rect 186686 0 186742 800
rect 188434 0 188490 800
rect 190182 0 190238 800
rect 191930 0 191986 800
rect 193678 0 193734 800
rect 195426 0 195482 800
rect 197174 0 197230 800
rect 198922 0 198978 800
rect 200670 0 200726 800
rect 202418 0 202474 800
rect 204166 0 204222 800
rect 205914 0 205970 800
rect 207662 0 207718 800
rect 209410 0 209466 800
rect 211158 0 211214 800
rect 212906 0 212962 800
rect 214654 0 214710 800
rect 216402 0 216458 800
rect 218150 0 218206 800
rect 219898 0 219954 800
rect 221646 0 221702 800
rect 223394 0 223450 800
rect 225142 0 225198 800
rect 226890 0 226946 800
rect 228638 0 228694 800
rect 230386 0 230442 800
rect 232134 0 232190 800
rect 233882 0 233938 800
rect 235630 0 235686 800
rect 237378 0 237434 800
rect 239126 0 239182 800
rect 240874 0 240930 800
rect 242622 0 242678 800
rect 244370 0 244426 800
rect 246118 0 246174 800
rect 247866 0 247922 800
rect 249614 0 249670 800
rect 251362 0 251418 800
rect 253110 0 253166 800
rect 254858 0 254914 800
rect 256606 0 256662 800
rect 258354 0 258410 800
rect 260102 0 260158 800
rect 261850 0 261906 800
rect 263598 0 263654 800
rect 265346 0 265402 800
rect 267094 0 267150 800
rect 268842 0 268898 800
rect 270590 0 270646 800
rect 272338 0 272394 800
rect 274086 0 274142 800
rect 275834 0 275890 800
rect 277582 0 277638 800
rect 279330 0 279386 800
rect 281078 0 281134 800
rect 282826 0 282882 800
rect 284574 0 284630 800
rect 286322 0 286378 800
rect 288070 0 288126 800
rect 289818 0 289874 800
rect 291566 0 291622 800
rect 293314 0 293370 800
rect 295062 0 295118 800
rect 296810 0 296866 800
rect 298558 0 298614 800
rect 300306 0 300362 800
rect 302054 0 302110 800
rect 303802 0 303858 800
rect 305550 0 305606 800
rect 307298 0 307354 800
rect 309046 0 309102 800
rect 310794 0 310850 800
rect 312542 0 312598 800
rect 314290 0 314346 800
rect 316038 0 316094 800
rect 317786 0 317842 800
rect 319534 0 319590 800
rect 321282 0 321338 800
rect 323030 0 323086 800
rect 324778 0 324834 800
rect 326526 0 326582 800
rect 328274 0 328330 800
rect 330022 0 330078 800
rect 331770 0 331826 800
rect 333518 0 333574 800
rect 335266 0 335322 800
rect 337014 0 337070 800
rect 338762 0 338818 800
rect 340510 0 340566 800
rect 342258 0 342314 800
rect 344006 0 344062 800
rect 345754 0 345810 800
rect 347502 0 347558 800
rect 349250 0 349306 800
rect 350998 0 351054 800
rect 352746 0 352802 800
rect 354494 0 354550 800
rect 356242 0 356298 800
rect 357990 0 358046 800
rect 359738 0 359794 800
rect 361486 0 361542 800
rect 363234 0 363290 800
rect 364982 0 365038 800
rect 366730 0 366786 800
rect 368478 0 368534 800
rect 370226 0 370282 800
rect 371974 0 372030 800
rect 373722 0 373778 800
rect 375470 0 375526 800
rect 377218 0 377274 800
rect 378966 0 379022 800
rect 380714 0 380770 800
rect 382462 0 382518 800
rect 384210 0 384266 800
rect 385958 0 386014 800
rect 387706 0 387762 800
rect 389454 0 389510 800
rect 391202 0 391258 800
rect 392950 0 393006 800
rect 394698 0 394754 800
rect 396446 0 396502 800
rect 398194 0 398250 800
rect 399942 0 399998 800
rect 401690 0 401746 800
rect 403438 0 403494 800
rect 405186 0 405242 800
rect 406934 0 406990 800
rect 408682 0 408738 800
rect 410430 0 410486 800
rect 412178 0 412234 800
rect 413926 0 413982 800
rect 415674 0 415730 800
rect 417422 0 417478 800
rect 419170 0 419226 800
rect 420918 0 420974 800
rect 422666 0 422722 800
rect 424414 0 424470 800
rect 426162 0 426218 800
rect 427910 0 427966 800
rect 429658 0 429714 800
rect 431406 0 431462 800
<< obsm2 >>
rect 1306 159144 8334 159730
rect 8502 159144 9346 159730
rect 9514 159144 10358 159730
rect 10526 159144 11370 159730
rect 11538 159144 12382 159730
rect 12550 159144 13394 159730
rect 13562 159144 14406 159730
rect 14574 159144 15418 159730
rect 15586 159144 16430 159730
rect 16598 159144 17442 159730
rect 17610 159144 18454 159730
rect 18622 159144 19466 159730
rect 19634 159144 20478 159730
rect 20646 159144 21490 159730
rect 21658 159144 22502 159730
rect 22670 159144 23514 159730
rect 23682 159144 24526 159730
rect 24694 159144 25538 159730
rect 25706 159144 26550 159730
rect 26718 159144 27562 159730
rect 27730 159144 28574 159730
rect 28742 159144 29586 159730
rect 29754 159144 30598 159730
rect 30766 159144 31610 159730
rect 31778 159144 32622 159730
rect 32790 159144 33634 159730
rect 33802 159144 34646 159730
rect 34814 159144 35658 159730
rect 35826 159144 36670 159730
rect 36838 159144 37682 159730
rect 37850 159144 38694 159730
rect 38862 159144 39706 159730
rect 39874 159144 40718 159730
rect 40886 159144 41730 159730
rect 41898 159144 42742 159730
rect 42910 159144 43754 159730
rect 43922 159144 44766 159730
rect 44934 159144 45778 159730
rect 45946 159144 46790 159730
rect 46958 159144 47802 159730
rect 47970 159144 48814 159730
rect 48982 159144 49826 159730
rect 49994 159144 50838 159730
rect 51006 159144 51850 159730
rect 52018 159144 52862 159730
rect 53030 159144 53874 159730
rect 54042 159144 54886 159730
rect 55054 159144 55898 159730
rect 56066 159144 56910 159730
rect 57078 159144 57922 159730
rect 58090 159144 58934 159730
rect 59102 159144 59946 159730
rect 60114 159144 60958 159730
rect 61126 159144 61970 159730
rect 62138 159144 62982 159730
rect 63150 159144 63994 159730
rect 64162 159144 65006 159730
rect 65174 159144 66018 159730
rect 66186 159144 67030 159730
rect 67198 159144 68042 159730
rect 68210 159144 69054 159730
rect 69222 159144 70066 159730
rect 70234 159144 71078 159730
rect 71246 159144 72090 159730
rect 72258 159144 73102 159730
rect 73270 159144 74114 159730
rect 74282 159144 75126 159730
rect 75294 159144 76138 159730
rect 76306 159144 77150 159730
rect 77318 159144 78162 159730
rect 78330 159144 79174 159730
rect 79342 159144 80186 159730
rect 80354 159144 81198 159730
rect 81366 159144 82210 159730
rect 82378 159144 83222 159730
rect 83390 159144 84234 159730
rect 84402 159144 85246 159730
rect 85414 159144 86258 159730
rect 86426 159144 87270 159730
rect 87438 159144 88282 159730
rect 88450 159144 89294 159730
rect 89462 159144 90306 159730
rect 90474 159144 91318 159730
rect 91486 159144 92330 159730
rect 92498 159144 93342 159730
rect 93510 159144 94354 159730
rect 94522 159144 95366 159730
rect 95534 159144 96378 159730
rect 96546 159144 97390 159730
rect 97558 159144 98402 159730
rect 98570 159144 99414 159730
rect 99582 159144 100426 159730
rect 100594 159144 101438 159730
rect 101606 159144 102450 159730
rect 102618 159144 103462 159730
rect 103630 159144 104474 159730
rect 104642 159144 105486 159730
rect 105654 159144 106498 159730
rect 106666 159144 107510 159730
rect 107678 159144 108522 159730
rect 108690 159144 109534 159730
rect 109702 159144 110546 159730
rect 110714 159144 111558 159730
rect 111726 159144 112570 159730
rect 112738 159144 113582 159730
rect 113750 159144 114594 159730
rect 114762 159144 115606 159730
rect 115774 159144 116618 159730
rect 116786 159144 117630 159730
rect 117798 159144 118642 159730
rect 118810 159144 119654 159730
rect 119822 159144 120666 159730
rect 120834 159144 121678 159730
rect 121846 159144 122690 159730
rect 122858 159144 123702 159730
rect 123870 159144 124714 159730
rect 124882 159144 125726 159730
rect 125894 159144 126738 159730
rect 126906 159144 127750 159730
rect 127918 159144 128762 159730
rect 128930 159144 129774 159730
rect 129942 159144 130786 159730
rect 130954 159144 131798 159730
rect 131966 159144 132810 159730
rect 132978 159144 133822 159730
rect 133990 159144 134834 159730
rect 135002 159144 135846 159730
rect 136014 159144 136858 159730
rect 137026 159144 137870 159730
rect 138038 159144 138882 159730
rect 139050 159144 139894 159730
rect 140062 159144 140906 159730
rect 141074 159144 141918 159730
rect 142086 159144 142930 159730
rect 143098 159144 143942 159730
rect 144110 159144 144954 159730
rect 145122 159144 145966 159730
rect 146134 159144 146978 159730
rect 147146 159144 147990 159730
rect 148158 159144 149002 159730
rect 149170 159144 150014 159730
rect 150182 159144 151026 159730
rect 151194 159144 152038 159730
rect 152206 159144 153050 159730
rect 153218 159144 154062 159730
rect 154230 159144 155074 159730
rect 155242 159144 156086 159730
rect 156254 159144 157098 159730
rect 157266 159144 158110 159730
rect 158278 159144 159122 159730
rect 159290 159144 160134 159730
rect 160302 159144 161146 159730
rect 161314 159144 162158 159730
rect 162326 159144 163170 159730
rect 163338 159144 164182 159730
rect 164350 159144 165194 159730
rect 165362 159144 166206 159730
rect 166374 159144 167218 159730
rect 167386 159144 168230 159730
rect 168398 159144 169242 159730
rect 169410 159144 170254 159730
rect 170422 159144 171266 159730
rect 171434 159144 172278 159730
rect 172446 159144 173290 159730
rect 173458 159144 174302 159730
rect 174470 159144 175314 159730
rect 175482 159144 176326 159730
rect 176494 159144 177338 159730
rect 177506 159144 178350 159730
rect 178518 159144 179362 159730
rect 179530 159144 180374 159730
rect 180542 159144 181386 159730
rect 181554 159144 182398 159730
rect 182566 159144 183410 159730
rect 183578 159144 184422 159730
rect 184590 159144 185434 159730
rect 185602 159144 186446 159730
rect 186614 159144 187458 159730
rect 187626 159144 188470 159730
rect 188638 159144 189482 159730
rect 189650 159144 190494 159730
rect 190662 159144 191506 159730
rect 191674 159144 192518 159730
rect 192686 159144 193530 159730
rect 193698 159144 194542 159730
rect 194710 159144 195554 159730
rect 195722 159144 196566 159730
rect 196734 159144 197578 159730
rect 197746 159144 198590 159730
rect 198758 159144 199602 159730
rect 199770 159144 200614 159730
rect 200782 159144 201626 159730
rect 201794 159144 202638 159730
rect 202806 159144 203650 159730
rect 203818 159144 204662 159730
rect 204830 159144 205674 159730
rect 205842 159144 206686 159730
rect 206854 159144 207698 159730
rect 207866 159144 208710 159730
rect 208878 159144 209722 159730
rect 209890 159144 210734 159730
rect 210902 159144 211746 159730
rect 211914 159144 212758 159730
rect 212926 159144 213770 159730
rect 213938 159144 214782 159730
rect 214950 159144 215794 159730
rect 215962 159144 216806 159730
rect 216974 159144 217818 159730
rect 217986 159144 218830 159730
rect 218998 159144 219842 159730
rect 220010 159144 220854 159730
rect 221022 159144 221866 159730
rect 222034 159144 222878 159730
rect 223046 159144 223890 159730
rect 224058 159144 224902 159730
rect 225070 159144 225914 159730
rect 226082 159144 226926 159730
rect 227094 159144 227938 159730
rect 228106 159144 228950 159730
rect 229118 159144 229962 159730
rect 230130 159144 230974 159730
rect 231142 159144 231986 159730
rect 232154 159144 232998 159730
rect 233166 159144 234010 159730
rect 234178 159144 235022 159730
rect 235190 159144 236034 159730
rect 236202 159144 237046 159730
rect 237214 159144 238058 159730
rect 238226 159144 239070 159730
rect 239238 159144 240082 159730
rect 240250 159144 241094 159730
rect 241262 159144 242106 159730
rect 242274 159144 243118 159730
rect 243286 159144 244130 159730
rect 244298 159144 245142 159730
rect 245310 159144 246154 159730
rect 246322 159144 247166 159730
rect 247334 159144 248178 159730
rect 248346 159144 249190 159730
rect 249358 159144 250202 159730
rect 250370 159144 251214 159730
rect 251382 159144 252226 159730
rect 252394 159144 253238 159730
rect 253406 159144 254250 159730
rect 254418 159144 255262 159730
rect 255430 159144 256274 159730
rect 256442 159144 257286 159730
rect 257454 159144 258298 159730
rect 258466 159144 259310 159730
rect 259478 159144 260322 159730
rect 260490 159144 261334 159730
rect 261502 159144 262346 159730
rect 262514 159144 263358 159730
rect 263526 159144 264370 159730
rect 264538 159144 265382 159730
rect 265550 159144 266394 159730
rect 266562 159144 267406 159730
rect 267574 159144 268418 159730
rect 268586 159144 269430 159730
rect 269598 159144 270442 159730
rect 270610 159144 271454 159730
rect 271622 159144 272466 159730
rect 272634 159144 273478 159730
rect 273646 159144 274490 159730
rect 274658 159144 275502 159730
rect 275670 159144 276514 159730
rect 276682 159144 277526 159730
rect 277694 159144 278538 159730
rect 278706 159144 279550 159730
rect 279718 159144 280562 159730
rect 280730 159144 281574 159730
rect 281742 159144 282586 159730
rect 282754 159144 283598 159730
rect 283766 159144 284610 159730
rect 284778 159144 285622 159730
rect 285790 159144 286634 159730
rect 286802 159144 287646 159730
rect 287814 159144 288658 159730
rect 288826 159144 289670 159730
rect 289838 159144 290682 159730
rect 290850 159144 291694 159730
rect 291862 159144 292706 159730
rect 292874 159144 293718 159730
rect 293886 159144 294730 159730
rect 294898 159144 295742 159730
rect 295910 159144 296754 159730
rect 296922 159144 297766 159730
rect 297934 159144 298778 159730
rect 298946 159144 299790 159730
rect 299958 159144 300802 159730
rect 300970 159144 301814 159730
rect 301982 159144 302826 159730
rect 302994 159144 303838 159730
rect 304006 159144 304850 159730
rect 305018 159144 305862 159730
rect 306030 159144 306874 159730
rect 307042 159144 307886 159730
rect 308054 159144 308898 159730
rect 309066 159144 309910 159730
rect 310078 159144 310922 159730
rect 311090 159144 311934 159730
rect 312102 159144 312946 159730
rect 313114 159144 313958 159730
rect 314126 159144 314970 159730
rect 315138 159144 315982 159730
rect 316150 159144 316994 159730
rect 317162 159144 318006 159730
rect 318174 159144 319018 159730
rect 319186 159144 320030 159730
rect 320198 159144 321042 159730
rect 321210 159144 322054 159730
rect 322222 159144 323066 159730
rect 323234 159144 324078 159730
rect 324246 159144 325090 159730
rect 325258 159144 326102 159730
rect 326270 159144 327114 159730
rect 327282 159144 328126 159730
rect 328294 159144 329138 159730
rect 329306 159144 330150 159730
rect 330318 159144 331162 159730
rect 331330 159144 332174 159730
rect 332342 159144 333186 159730
rect 333354 159144 334198 159730
rect 334366 159144 335210 159730
rect 335378 159144 336222 159730
rect 336390 159144 337234 159730
rect 337402 159144 338246 159730
rect 338414 159144 339258 159730
rect 339426 159144 340270 159730
rect 340438 159144 341282 159730
rect 341450 159144 342294 159730
rect 342462 159144 343306 159730
rect 343474 159144 344318 159730
rect 344486 159144 345330 159730
rect 345498 159144 346342 159730
rect 346510 159144 347354 159730
rect 347522 159144 348366 159730
rect 348534 159144 349378 159730
rect 349546 159144 350390 159730
rect 350558 159144 351402 159730
rect 351570 159144 352414 159730
rect 352582 159144 353426 159730
rect 353594 159144 354438 159730
rect 354606 159144 355450 159730
rect 355618 159144 356462 159730
rect 356630 159144 357474 159730
rect 357642 159144 358486 159730
rect 358654 159144 359498 159730
rect 359666 159144 360510 159730
rect 360678 159144 361522 159730
rect 361690 159144 362534 159730
rect 362702 159144 363546 159730
rect 363714 159144 364558 159730
rect 364726 159144 365570 159730
rect 365738 159144 366582 159730
rect 366750 159144 367594 159730
rect 367762 159144 368606 159730
rect 368774 159144 369618 159730
rect 369786 159144 370630 159730
rect 370798 159144 371642 159730
rect 371810 159144 372654 159730
rect 372822 159144 373666 159730
rect 373834 159144 374678 159730
rect 374846 159144 375690 159730
rect 375858 159144 376702 159730
rect 376870 159144 377714 159730
rect 377882 159144 378726 159730
rect 378894 159144 379738 159730
rect 379906 159144 380750 159730
rect 380918 159144 381762 159730
rect 381930 159144 382774 159730
rect 382942 159144 383786 159730
rect 383954 159144 384798 159730
rect 384966 159144 385810 159730
rect 385978 159144 386822 159730
rect 386990 159144 387834 159730
rect 388002 159144 388846 159730
rect 389014 159144 389858 159730
rect 390026 159144 390870 159730
rect 391038 159144 391882 159730
rect 392050 159144 392894 159730
rect 393062 159144 393906 159730
rect 394074 159144 394918 159730
rect 395086 159144 395930 159730
rect 396098 159144 396942 159730
rect 397110 159144 397954 159730
rect 398122 159144 398966 159730
rect 399134 159144 399978 159730
rect 400146 159144 400990 159730
rect 401158 159144 402002 159730
rect 402170 159144 403014 159730
rect 403182 159144 404026 159730
rect 404194 159144 405038 159730
rect 405206 159144 406050 159730
rect 406218 159144 407062 159730
rect 407230 159144 408074 159730
rect 408242 159144 409086 159730
rect 409254 159144 410098 159730
rect 410266 159144 411110 159730
rect 411278 159144 412122 159730
rect 412290 159144 413134 159730
rect 413302 159144 414146 159730
rect 414314 159144 415158 159730
rect 415326 159144 416170 159730
rect 416338 159144 417182 159730
rect 417350 159144 418194 159730
rect 418362 159144 419206 159730
rect 419374 159144 420218 159730
rect 420386 159144 421230 159730
rect 421398 159144 422242 159730
rect 422410 159144 423254 159730
rect 423422 159144 424266 159730
rect 424434 159144 425278 159730
rect 425446 159144 426290 159730
rect 426458 159144 427302 159730
rect 427470 159144 428314 159730
rect 428482 159144 429326 159730
rect 429494 159144 430338 159730
rect 430506 159144 431350 159730
rect 431518 159144 439372 159730
rect 1306 856 439372 159144
rect 1306 70 8334 856
rect 8502 70 10082 856
rect 10250 70 11830 856
rect 11998 70 13578 856
rect 13746 70 15326 856
rect 15494 70 17074 856
rect 17242 70 18822 856
rect 18990 70 20570 856
rect 20738 70 22318 856
rect 22486 70 24066 856
rect 24234 70 25814 856
rect 25982 70 27562 856
rect 27730 70 29310 856
rect 29478 70 31058 856
rect 31226 70 32806 856
rect 32974 70 34554 856
rect 34722 70 36302 856
rect 36470 70 38050 856
rect 38218 70 39798 856
rect 39966 70 41546 856
rect 41714 70 43294 856
rect 43462 70 45042 856
rect 45210 70 46790 856
rect 46958 70 48538 856
rect 48706 70 50286 856
rect 50454 70 52034 856
rect 52202 70 53782 856
rect 53950 70 55530 856
rect 55698 70 57278 856
rect 57446 70 59026 856
rect 59194 70 60774 856
rect 60942 70 62522 856
rect 62690 70 64270 856
rect 64438 70 66018 856
rect 66186 70 67766 856
rect 67934 70 69514 856
rect 69682 70 71262 856
rect 71430 70 73010 856
rect 73178 70 74758 856
rect 74926 70 76506 856
rect 76674 70 78254 856
rect 78422 70 80002 856
rect 80170 70 81750 856
rect 81918 70 83498 856
rect 83666 70 85246 856
rect 85414 70 86994 856
rect 87162 70 88742 856
rect 88910 70 90490 856
rect 90658 70 92238 856
rect 92406 70 93986 856
rect 94154 70 95734 856
rect 95902 70 97482 856
rect 97650 70 99230 856
rect 99398 70 100978 856
rect 101146 70 102726 856
rect 102894 70 104474 856
rect 104642 70 106222 856
rect 106390 70 107970 856
rect 108138 70 109718 856
rect 109886 70 111466 856
rect 111634 70 113214 856
rect 113382 70 114962 856
rect 115130 70 116710 856
rect 116878 70 118458 856
rect 118626 70 120206 856
rect 120374 70 121954 856
rect 122122 70 123702 856
rect 123870 70 125450 856
rect 125618 70 127198 856
rect 127366 70 128946 856
rect 129114 70 130694 856
rect 130862 70 132442 856
rect 132610 70 134190 856
rect 134358 70 135938 856
rect 136106 70 137686 856
rect 137854 70 139434 856
rect 139602 70 141182 856
rect 141350 70 142930 856
rect 143098 70 144678 856
rect 144846 70 146426 856
rect 146594 70 148174 856
rect 148342 70 149922 856
rect 150090 70 151670 856
rect 151838 70 153418 856
rect 153586 70 155166 856
rect 155334 70 156914 856
rect 157082 70 158662 856
rect 158830 70 160410 856
rect 160578 70 162158 856
rect 162326 70 163906 856
rect 164074 70 165654 856
rect 165822 70 167402 856
rect 167570 70 169150 856
rect 169318 70 170898 856
rect 171066 70 172646 856
rect 172814 70 174394 856
rect 174562 70 176142 856
rect 176310 70 177890 856
rect 178058 70 179638 856
rect 179806 70 181386 856
rect 181554 70 183134 856
rect 183302 70 184882 856
rect 185050 70 186630 856
rect 186798 70 188378 856
rect 188546 70 190126 856
rect 190294 70 191874 856
rect 192042 70 193622 856
rect 193790 70 195370 856
rect 195538 70 197118 856
rect 197286 70 198866 856
rect 199034 70 200614 856
rect 200782 70 202362 856
rect 202530 70 204110 856
rect 204278 70 205858 856
rect 206026 70 207606 856
rect 207774 70 209354 856
rect 209522 70 211102 856
rect 211270 70 212850 856
rect 213018 70 214598 856
rect 214766 70 216346 856
rect 216514 70 218094 856
rect 218262 70 219842 856
rect 220010 70 221590 856
rect 221758 70 223338 856
rect 223506 70 225086 856
rect 225254 70 226834 856
rect 227002 70 228582 856
rect 228750 70 230330 856
rect 230498 70 232078 856
rect 232246 70 233826 856
rect 233994 70 235574 856
rect 235742 70 237322 856
rect 237490 70 239070 856
rect 239238 70 240818 856
rect 240986 70 242566 856
rect 242734 70 244314 856
rect 244482 70 246062 856
rect 246230 70 247810 856
rect 247978 70 249558 856
rect 249726 70 251306 856
rect 251474 70 253054 856
rect 253222 70 254802 856
rect 254970 70 256550 856
rect 256718 70 258298 856
rect 258466 70 260046 856
rect 260214 70 261794 856
rect 261962 70 263542 856
rect 263710 70 265290 856
rect 265458 70 267038 856
rect 267206 70 268786 856
rect 268954 70 270534 856
rect 270702 70 272282 856
rect 272450 70 274030 856
rect 274198 70 275778 856
rect 275946 70 277526 856
rect 277694 70 279274 856
rect 279442 70 281022 856
rect 281190 70 282770 856
rect 282938 70 284518 856
rect 284686 70 286266 856
rect 286434 70 288014 856
rect 288182 70 289762 856
rect 289930 70 291510 856
rect 291678 70 293258 856
rect 293426 70 295006 856
rect 295174 70 296754 856
rect 296922 70 298502 856
rect 298670 70 300250 856
rect 300418 70 301998 856
rect 302166 70 303746 856
rect 303914 70 305494 856
rect 305662 70 307242 856
rect 307410 70 308990 856
rect 309158 70 310738 856
rect 310906 70 312486 856
rect 312654 70 314234 856
rect 314402 70 315982 856
rect 316150 70 317730 856
rect 317898 70 319478 856
rect 319646 70 321226 856
rect 321394 70 322974 856
rect 323142 70 324722 856
rect 324890 70 326470 856
rect 326638 70 328218 856
rect 328386 70 329966 856
rect 330134 70 331714 856
rect 331882 70 333462 856
rect 333630 70 335210 856
rect 335378 70 336958 856
rect 337126 70 338706 856
rect 338874 70 340454 856
rect 340622 70 342202 856
rect 342370 70 343950 856
rect 344118 70 345698 856
rect 345866 70 347446 856
rect 347614 70 349194 856
rect 349362 70 350942 856
rect 351110 70 352690 856
rect 352858 70 354438 856
rect 354606 70 356186 856
rect 356354 70 357934 856
rect 358102 70 359682 856
rect 359850 70 361430 856
rect 361598 70 363178 856
rect 363346 70 364926 856
rect 365094 70 366674 856
rect 366842 70 368422 856
rect 368590 70 370170 856
rect 370338 70 371918 856
rect 372086 70 373666 856
rect 373834 70 375414 856
rect 375582 70 377162 856
rect 377330 70 378910 856
rect 379078 70 380658 856
rect 380826 70 382406 856
rect 382574 70 384154 856
rect 384322 70 385902 856
rect 386070 70 387650 856
rect 387818 70 389398 856
rect 389566 70 391146 856
rect 391314 70 392894 856
rect 393062 70 394642 856
rect 394810 70 396390 856
rect 396558 70 398138 856
rect 398306 70 399886 856
rect 400054 70 401634 856
rect 401802 70 403382 856
rect 403550 70 405130 856
rect 405298 70 406878 856
rect 407046 70 408626 856
rect 408794 70 410374 856
rect 410542 70 412122 856
rect 412290 70 413870 856
rect 414038 70 415618 856
rect 415786 70 417366 856
rect 417534 70 419114 856
rect 419282 70 420862 856
rect 421030 70 422610 856
rect 422778 70 424358 856
rect 424526 70 426106 856
rect 426274 70 427854 856
rect 428022 70 429602 856
rect 429770 70 431350 856
rect 431518 70 439372 856
<< metal3 >>
rect 439200 144168 440000 144288
rect 439200 143624 440000 143744
rect 0 143080 800 143200
rect 439200 143080 440000 143200
rect 0 142536 800 142656
rect 439200 142536 440000 142656
rect 0 141992 800 142112
rect 439200 141992 440000 142112
rect 0 141448 800 141568
rect 439200 141448 440000 141568
rect 0 140904 800 141024
rect 439200 140904 440000 141024
rect 0 140360 800 140480
rect 439200 140360 440000 140480
rect 0 139816 800 139936
rect 439200 139816 440000 139936
rect 0 139272 800 139392
rect 439200 139272 440000 139392
rect 0 138728 800 138848
rect 439200 138728 440000 138848
rect 0 138184 800 138304
rect 439200 138184 440000 138304
rect 0 137640 800 137760
rect 439200 137640 440000 137760
rect 0 137096 800 137216
rect 439200 137096 440000 137216
rect 0 136552 800 136672
rect 439200 136552 440000 136672
rect 0 136008 800 136128
rect 439200 136008 440000 136128
rect 0 135464 800 135584
rect 439200 135464 440000 135584
rect 0 134920 800 135040
rect 439200 134920 440000 135040
rect 0 134376 800 134496
rect 439200 134376 440000 134496
rect 0 133832 800 133952
rect 439200 133832 440000 133952
rect 0 133288 800 133408
rect 439200 133288 440000 133408
rect 0 132744 800 132864
rect 439200 132744 440000 132864
rect 0 132200 800 132320
rect 439200 132200 440000 132320
rect 0 131656 800 131776
rect 439200 131656 440000 131776
rect 0 131112 800 131232
rect 439200 131112 440000 131232
rect 0 130568 800 130688
rect 439200 130568 440000 130688
rect 0 130024 800 130144
rect 439200 130024 440000 130144
rect 0 129480 800 129600
rect 439200 129480 440000 129600
rect 0 128936 800 129056
rect 439200 128936 440000 129056
rect 0 128392 800 128512
rect 439200 128392 440000 128512
rect 0 127848 800 127968
rect 439200 127848 440000 127968
rect 0 127304 800 127424
rect 439200 127304 440000 127424
rect 0 126760 800 126880
rect 439200 126760 440000 126880
rect 0 126216 800 126336
rect 439200 126216 440000 126336
rect 0 125672 800 125792
rect 439200 125672 440000 125792
rect 0 125128 800 125248
rect 439200 125128 440000 125248
rect 0 124584 800 124704
rect 439200 124584 440000 124704
rect 0 124040 800 124160
rect 439200 124040 440000 124160
rect 0 123496 800 123616
rect 439200 123496 440000 123616
rect 0 122952 800 123072
rect 439200 122952 440000 123072
rect 0 122408 800 122528
rect 439200 122408 440000 122528
rect 0 121864 800 121984
rect 439200 121864 440000 121984
rect 0 121320 800 121440
rect 439200 121320 440000 121440
rect 0 120776 800 120896
rect 439200 120776 440000 120896
rect 0 120232 800 120352
rect 439200 120232 440000 120352
rect 0 119688 800 119808
rect 439200 119688 440000 119808
rect 0 119144 800 119264
rect 439200 119144 440000 119264
rect 0 118600 800 118720
rect 439200 118600 440000 118720
rect 0 118056 800 118176
rect 439200 118056 440000 118176
rect 0 117512 800 117632
rect 439200 117512 440000 117632
rect 0 116968 800 117088
rect 439200 116968 440000 117088
rect 0 116424 800 116544
rect 439200 116424 440000 116544
rect 0 115880 800 116000
rect 439200 115880 440000 116000
rect 0 115336 800 115456
rect 439200 115336 440000 115456
rect 0 114792 800 114912
rect 439200 114792 440000 114912
rect 0 114248 800 114368
rect 439200 114248 440000 114368
rect 0 113704 800 113824
rect 439200 113704 440000 113824
rect 0 113160 800 113280
rect 439200 113160 440000 113280
rect 0 112616 800 112736
rect 439200 112616 440000 112736
rect 0 112072 800 112192
rect 439200 112072 440000 112192
rect 0 111528 800 111648
rect 439200 111528 440000 111648
rect 0 110984 800 111104
rect 439200 110984 440000 111104
rect 0 110440 800 110560
rect 439200 110440 440000 110560
rect 0 109896 800 110016
rect 439200 109896 440000 110016
rect 0 109352 800 109472
rect 439200 109352 440000 109472
rect 0 108808 800 108928
rect 439200 108808 440000 108928
rect 0 108264 800 108384
rect 439200 108264 440000 108384
rect 0 107720 800 107840
rect 439200 107720 440000 107840
rect 0 107176 800 107296
rect 439200 107176 440000 107296
rect 0 106632 800 106752
rect 439200 106632 440000 106752
rect 0 106088 800 106208
rect 439200 106088 440000 106208
rect 0 105544 800 105664
rect 439200 105544 440000 105664
rect 0 105000 800 105120
rect 439200 105000 440000 105120
rect 0 104456 800 104576
rect 439200 104456 440000 104576
rect 0 103912 800 104032
rect 439200 103912 440000 104032
rect 0 103368 800 103488
rect 439200 103368 440000 103488
rect 0 102824 800 102944
rect 439200 102824 440000 102944
rect 0 102280 800 102400
rect 439200 102280 440000 102400
rect 0 101736 800 101856
rect 439200 101736 440000 101856
rect 0 101192 800 101312
rect 439200 101192 440000 101312
rect 0 100648 800 100768
rect 439200 100648 440000 100768
rect 0 100104 800 100224
rect 439200 100104 440000 100224
rect 0 99560 800 99680
rect 439200 99560 440000 99680
rect 0 99016 800 99136
rect 439200 99016 440000 99136
rect 0 98472 800 98592
rect 439200 98472 440000 98592
rect 0 97928 800 98048
rect 439200 97928 440000 98048
rect 0 97384 800 97504
rect 439200 97384 440000 97504
rect 0 96840 800 96960
rect 439200 96840 440000 96960
rect 0 96296 800 96416
rect 439200 96296 440000 96416
rect 0 95752 800 95872
rect 439200 95752 440000 95872
rect 0 95208 800 95328
rect 439200 95208 440000 95328
rect 0 94664 800 94784
rect 439200 94664 440000 94784
rect 0 94120 800 94240
rect 439200 94120 440000 94240
rect 0 93576 800 93696
rect 439200 93576 440000 93696
rect 0 93032 800 93152
rect 439200 93032 440000 93152
rect 0 92488 800 92608
rect 439200 92488 440000 92608
rect 0 91944 800 92064
rect 439200 91944 440000 92064
rect 0 91400 800 91520
rect 439200 91400 440000 91520
rect 0 90856 800 90976
rect 439200 90856 440000 90976
rect 0 90312 800 90432
rect 439200 90312 440000 90432
rect 0 89768 800 89888
rect 439200 89768 440000 89888
rect 0 89224 800 89344
rect 439200 89224 440000 89344
rect 0 88680 800 88800
rect 439200 88680 440000 88800
rect 0 88136 800 88256
rect 439200 88136 440000 88256
rect 0 87592 800 87712
rect 439200 87592 440000 87712
rect 0 87048 800 87168
rect 439200 87048 440000 87168
rect 0 86504 800 86624
rect 439200 86504 440000 86624
rect 0 85960 800 86080
rect 439200 85960 440000 86080
rect 0 85416 800 85536
rect 439200 85416 440000 85536
rect 0 84872 800 84992
rect 439200 84872 440000 84992
rect 0 84328 800 84448
rect 439200 84328 440000 84448
rect 0 83784 800 83904
rect 439200 83784 440000 83904
rect 0 83240 800 83360
rect 439200 83240 440000 83360
rect 0 82696 800 82816
rect 439200 82696 440000 82816
rect 0 82152 800 82272
rect 439200 82152 440000 82272
rect 0 81608 800 81728
rect 439200 81608 440000 81728
rect 0 81064 800 81184
rect 439200 81064 440000 81184
rect 0 80520 800 80640
rect 439200 80520 440000 80640
rect 0 79976 800 80096
rect 439200 79976 440000 80096
rect 0 79432 800 79552
rect 439200 79432 440000 79552
rect 0 78888 800 79008
rect 439200 78888 440000 79008
rect 0 78344 800 78464
rect 439200 78344 440000 78464
rect 0 77800 800 77920
rect 439200 77800 440000 77920
rect 0 77256 800 77376
rect 439200 77256 440000 77376
rect 0 76712 800 76832
rect 439200 76712 440000 76832
rect 0 76168 800 76288
rect 439200 76168 440000 76288
rect 0 75624 800 75744
rect 439200 75624 440000 75744
rect 0 75080 800 75200
rect 439200 75080 440000 75200
rect 0 74536 800 74656
rect 439200 74536 440000 74656
rect 0 73992 800 74112
rect 439200 73992 440000 74112
rect 0 73448 800 73568
rect 439200 73448 440000 73568
rect 0 72904 800 73024
rect 439200 72904 440000 73024
rect 0 72360 800 72480
rect 439200 72360 440000 72480
rect 0 71816 800 71936
rect 439200 71816 440000 71936
rect 0 71272 800 71392
rect 439200 71272 440000 71392
rect 0 70728 800 70848
rect 439200 70728 440000 70848
rect 0 70184 800 70304
rect 439200 70184 440000 70304
rect 0 69640 800 69760
rect 439200 69640 440000 69760
rect 0 69096 800 69216
rect 439200 69096 440000 69216
rect 0 68552 800 68672
rect 439200 68552 440000 68672
rect 0 68008 800 68128
rect 439200 68008 440000 68128
rect 0 67464 800 67584
rect 439200 67464 440000 67584
rect 0 66920 800 67040
rect 439200 66920 440000 67040
rect 0 66376 800 66496
rect 439200 66376 440000 66496
rect 0 65832 800 65952
rect 439200 65832 440000 65952
rect 0 65288 800 65408
rect 439200 65288 440000 65408
rect 0 64744 800 64864
rect 439200 64744 440000 64864
rect 0 64200 800 64320
rect 439200 64200 440000 64320
rect 0 63656 800 63776
rect 439200 63656 440000 63776
rect 0 63112 800 63232
rect 439200 63112 440000 63232
rect 0 62568 800 62688
rect 439200 62568 440000 62688
rect 0 62024 800 62144
rect 439200 62024 440000 62144
rect 0 61480 800 61600
rect 439200 61480 440000 61600
rect 0 60936 800 61056
rect 439200 60936 440000 61056
rect 0 60392 800 60512
rect 439200 60392 440000 60512
rect 0 59848 800 59968
rect 439200 59848 440000 59968
rect 0 59304 800 59424
rect 439200 59304 440000 59424
rect 0 58760 800 58880
rect 439200 58760 440000 58880
rect 0 58216 800 58336
rect 439200 58216 440000 58336
rect 0 57672 800 57792
rect 439200 57672 440000 57792
rect 0 57128 800 57248
rect 439200 57128 440000 57248
rect 0 56584 800 56704
rect 439200 56584 440000 56704
rect 0 56040 800 56160
rect 439200 56040 440000 56160
rect 0 55496 800 55616
rect 439200 55496 440000 55616
rect 0 54952 800 55072
rect 439200 54952 440000 55072
rect 0 54408 800 54528
rect 439200 54408 440000 54528
rect 0 53864 800 53984
rect 439200 53864 440000 53984
rect 0 53320 800 53440
rect 439200 53320 440000 53440
rect 0 52776 800 52896
rect 439200 52776 440000 52896
rect 0 52232 800 52352
rect 439200 52232 440000 52352
rect 0 51688 800 51808
rect 439200 51688 440000 51808
rect 0 51144 800 51264
rect 439200 51144 440000 51264
rect 0 50600 800 50720
rect 439200 50600 440000 50720
rect 0 50056 800 50176
rect 439200 50056 440000 50176
rect 0 49512 800 49632
rect 439200 49512 440000 49632
rect 0 48968 800 49088
rect 439200 48968 440000 49088
rect 0 48424 800 48544
rect 439200 48424 440000 48544
rect 0 47880 800 48000
rect 439200 47880 440000 48000
rect 0 47336 800 47456
rect 439200 47336 440000 47456
rect 0 46792 800 46912
rect 439200 46792 440000 46912
rect 0 46248 800 46368
rect 439200 46248 440000 46368
rect 0 45704 800 45824
rect 439200 45704 440000 45824
rect 0 45160 800 45280
rect 439200 45160 440000 45280
rect 0 44616 800 44736
rect 439200 44616 440000 44736
rect 0 44072 800 44192
rect 439200 44072 440000 44192
rect 0 43528 800 43648
rect 439200 43528 440000 43648
rect 0 42984 800 43104
rect 439200 42984 440000 43104
rect 0 42440 800 42560
rect 439200 42440 440000 42560
rect 0 41896 800 42016
rect 439200 41896 440000 42016
rect 0 41352 800 41472
rect 439200 41352 440000 41472
rect 0 40808 800 40928
rect 439200 40808 440000 40928
rect 0 40264 800 40384
rect 439200 40264 440000 40384
rect 0 39720 800 39840
rect 439200 39720 440000 39840
rect 0 39176 800 39296
rect 439200 39176 440000 39296
rect 0 38632 800 38752
rect 439200 38632 440000 38752
rect 0 38088 800 38208
rect 439200 38088 440000 38208
rect 0 37544 800 37664
rect 439200 37544 440000 37664
rect 0 37000 800 37120
rect 439200 37000 440000 37120
rect 0 36456 800 36576
rect 439200 36456 440000 36576
rect 0 35912 800 36032
rect 439200 35912 440000 36032
rect 0 35368 800 35488
rect 439200 35368 440000 35488
rect 0 34824 800 34944
rect 439200 34824 440000 34944
rect 0 34280 800 34400
rect 439200 34280 440000 34400
rect 0 33736 800 33856
rect 439200 33736 440000 33856
rect 0 33192 800 33312
rect 439200 33192 440000 33312
rect 0 32648 800 32768
rect 439200 32648 440000 32768
rect 0 32104 800 32224
rect 439200 32104 440000 32224
rect 0 31560 800 31680
rect 439200 31560 440000 31680
rect 0 31016 800 31136
rect 439200 31016 440000 31136
rect 0 30472 800 30592
rect 439200 30472 440000 30592
rect 0 29928 800 30048
rect 439200 29928 440000 30048
rect 0 29384 800 29504
rect 439200 29384 440000 29504
rect 0 28840 800 28960
rect 439200 28840 440000 28960
rect 0 28296 800 28416
rect 439200 28296 440000 28416
rect 0 27752 800 27872
rect 439200 27752 440000 27872
rect 0 27208 800 27328
rect 439200 27208 440000 27328
rect 0 26664 800 26784
rect 439200 26664 440000 26784
rect 0 26120 800 26240
rect 439200 26120 440000 26240
rect 0 25576 800 25696
rect 439200 25576 440000 25696
rect 0 25032 800 25152
rect 439200 25032 440000 25152
rect 0 24488 800 24608
rect 439200 24488 440000 24608
rect 0 23944 800 24064
rect 439200 23944 440000 24064
rect 0 23400 800 23520
rect 439200 23400 440000 23520
rect 0 22856 800 22976
rect 439200 22856 440000 22976
rect 0 22312 800 22432
rect 439200 22312 440000 22432
rect 0 21768 800 21888
rect 439200 21768 440000 21888
rect 0 21224 800 21344
rect 439200 21224 440000 21344
rect 0 20680 800 20800
rect 439200 20680 440000 20800
rect 0 20136 800 20256
rect 439200 20136 440000 20256
rect 0 19592 800 19712
rect 439200 19592 440000 19712
rect 0 19048 800 19168
rect 439200 19048 440000 19168
rect 0 18504 800 18624
rect 439200 18504 440000 18624
rect 0 17960 800 18080
rect 439200 17960 440000 18080
rect 0 17416 800 17536
rect 439200 17416 440000 17536
rect 0 16872 800 16992
rect 439200 16872 440000 16992
rect 0 16328 800 16448
rect 439200 16328 440000 16448
rect 439200 15784 440000 15904
rect 439200 15240 440000 15360
<< obsm3 >>
rect 800 144368 439200 159357
rect 800 144088 439120 144368
rect 800 143824 439200 144088
rect 800 143544 439120 143824
rect 800 143280 439200 143544
rect 880 143000 439120 143280
rect 800 142736 439200 143000
rect 880 142456 439120 142736
rect 800 142192 439200 142456
rect 880 141912 439120 142192
rect 800 141648 439200 141912
rect 880 141368 439120 141648
rect 800 141104 439200 141368
rect 880 140824 439120 141104
rect 800 140560 439200 140824
rect 880 140280 439120 140560
rect 800 140016 439200 140280
rect 880 139736 439120 140016
rect 800 139472 439200 139736
rect 880 139192 439120 139472
rect 800 138928 439200 139192
rect 880 138648 439120 138928
rect 800 138384 439200 138648
rect 880 138104 439120 138384
rect 800 137840 439200 138104
rect 880 137560 439120 137840
rect 800 137296 439200 137560
rect 880 137016 439120 137296
rect 800 136752 439200 137016
rect 880 136472 439120 136752
rect 800 136208 439200 136472
rect 880 135928 439120 136208
rect 800 135664 439200 135928
rect 880 135384 439120 135664
rect 800 135120 439200 135384
rect 880 134840 439120 135120
rect 800 134576 439200 134840
rect 880 134296 439120 134576
rect 800 134032 439200 134296
rect 880 133752 439120 134032
rect 800 133488 439200 133752
rect 880 133208 439120 133488
rect 800 132944 439200 133208
rect 880 132664 439120 132944
rect 800 132400 439200 132664
rect 880 132120 439120 132400
rect 800 131856 439200 132120
rect 880 131576 439120 131856
rect 800 131312 439200 131576
rect 880 131032 439120 131312
rect 800 130768 439200 131032
rect 880 130488 439120 130768
rect 800 130224 439200 130488
rect 880 129944 439120 130224
rect 800 129680 439200 129944
rect 880 129400 439120 129680
rect 800 129136 439200 129400
rect 880 128856 439120 129136
rect 800 128592 439200 128856
rect 880 128312 439120 128592
rect 800 128048 439200 128312
rect 880 127768 439120 128048
rect 800 127504 439200 127768
rect 880 127224 439120 127504
rect 800 126960 439200 127224
rect 880 126680 439120 126960
rect 800 126416 439200 126680
rect 880 126136 439120 126416
rect 800 125872 439200 126136
rect 880 125592 439120 125872
rect 800 125328 439200 125592
rect 880 125048 439120 125328
rect 800 124784 439200 125048
rect 880 124504 439120 124784
rect 800 124240 439200 124504
rect 880 123960 439120 124240
rect 800 123696 439200 123960
rect 880 123416 439120 123696
rect 800 123152 439200 123416
rect 880 122872 439120 123152
rect 800 122608 439200 122872
rect 880 122328 439120 122608
rect 800 122064 439200 122328
rect 880 121784 439120 122064
rect 800 121520 439200 121784
rect 880 121240 439120 121520
rect 800 120976 439200 121240
rect 880 120696 439120 120976
rect 800 120432 439200 120696
rect 880 120152 439120 120432
rect 800 119888 439200 120152
rect 880 119608 439120 119888
rect 800 119344 439200 119608
rect 880 119064 439120 119344
rect 800 118800 439200 119064
rect 880 118520 439120 118800
rect 800 118256 439200 118520
rect 880 117976 439120 118256
rect 800 117712 439200 117976
rect 880 117432 439120 117712
rect 800 117168 439200 117432
rect 880 116888 439120 117168
rect 800 116624 439200 116888
rect 880 116344 439120 116624
rect 800 116080 439200 116344
rect 880 115800 439120 116080
rect 800 115536 439200 115800
rect 880 115256 439120 115536
rect 800 114992 439200 115256
rect 880 114712 439120 114992
rect 800 114448 439200 114712
rect 880 114168 439120 114448
rect 800 113904 439200 114168
rect 880 113624 439120 113904
rect 800 113360 439200 113624
rect 880 113080 439120 113360
rect 800 112816 439200 113080
rect 880 112536 439120 112816
rect 800 112272 439200 112536
rect 880 111992 439120 112272
rect 800 111728 439200 111992
rect 880 111448 439120 111728
rect 800 111184 439200 111448
rect 880 110904 439120 111184
rect 800 110640 439200 110904
rect 880 110360 439120 110640
rect 800 110096 439200 110360
rect 880 109816 439120 110096
rect 800 109552 439200 109816
rect 880 109272 439120 109552
rect 800 109008 439200 109272
rect 880 108728 439120 109008
rect 800 108464 439200 108728
rect 880 108184 439120 108464
rect 800 107920 439200 108184
rect 880 107640 439120 107920
rect 800 107376 439200 107640
rect 880 107096 439120 107376
rect 800 106832 439200 107096
rect 880 106552 439120 106832
rect 800 106288 439200 106552
rect 880 106008 439120 106288
rect 800 105744 439200 106008
rect 880 105464 439120 105744
rect 800 105200 439200 105464
rect 880 104920 439120 105200
rect 800 104656 439200 104920
rect 880 104376 439120 104656
rect 800 104112 439200 104376
rect 880 103832 439120 104112
rect 800 103568 439200 103832
rect 880 103288 439120 103568
rect 800 103024 439200 103288
rect 880 102744 439120 103024
rect 800 102480 439200 102744
rect 880 102200 439120 102480
rect 800 101936 439200 102200
rect 880 101656 439120 101936
rect 800 101392 439200 101656
rect 880 101112 439120 101392
rect 800 100848 439200 101112
rect 880 100568 439120 100848
rect 800 100304 439200 100568
rect 880 100024 439120 100304
rect 800 99760 439200 100024
rect 880 99480 439120 99760
rect 800 99216 439200 99480
rect 880 98936 439120 99216
rect 800 98672 439200 98936
rect 880 98392 439120 98672
rect 800 98128 439200 98392
rect 880 97848 439120 98128
rect 800 97584 439200 97848
rect 880 97304 439120 97584
rect 800 97040 439200 97304
rect 880 96760 439120 97040
rect 800 96496 439200 96760
rect 880 96216 439120 96496
rect 800 95952 439200 96216
rect 880 95672 439120 95952
rect 800 95408 439200 95672
rect 880 95128 439120 95408
rect 800 94864 439200 95128
rect 880 94584 439120 94864
rect 800 94320 439200 94584
rect 880 94040 439120 94320
rect 800 93776 439200 94040
rect 880 93496 439120 93776
rect 800 93232 439200 93496
rect 880 92952 439120 93232
rect 800 92688 439200 92952
rect 880 92408 439120 92688
rect 800 92144 439200 92408
rect 880 91864 439120 92144
rect 800 91600 439200 91864
rect 880 91320 439120 91600
rect 800 91056 439200 91320
rect 880 90776 439120 91056
rect 800 90512 439200 90776
rect 880 90232 439120 90512
rect 800 89968 439200 90232
rect 880 89688 439120 89968
rect 800 89424 439200 89688
rect 880 89144 439120 89424
rect 800 88880 439200 89144
rect 880 88600 439120 88880
rect 800 88336 439200 88600
rect 880 88056 439120 88336
rect 800 87792 439200 88056
rect 880 87512 439120 87792
rect 800 87248 439200 87512
rect 880 86968 439120 87248
rect 800 86704 439200 86968
rect 880 86424 439120 86704
rect 800 86160 439200 86424
rect 880 85880 439120 86160
rect 800 85616 439200 85880
rect 880 85336 439120 85616
rect 800 85072 439200 85336
rect 880 84792 439120 85072
rect 800 84528 439200 84792
rect 880 84248 439120 84528
rect 800 83984 439200 84248
rect 880 83704 439120 83984
rect 800 83440 439200 83704
rect 880 83160 439120 83440
rect 800 82896 439200 83160
rect 880 82616 439120 82896
rect 800 82352 439200 82616
rect 880 82072 439120 82352
rect 800 81808 439200 82072
rect 880 81528 439120 81808
rect 800 81264 439200 81528
rect 880 80984 439120 81264
rect 800 80720 439200 80984
rect 880 80440 439120 80720
rect 800 80176 439200 80440
rect 880 79896 439120 80176
rect 800 79632 439200 79896
rect 880 79352 439120 79632
rect 800 79088 439200 79352
rect 880 78808 439120 79088
rect 800 78544 439200 78808
rect 880 78264 439120 78544
rect 800 78000 439200 78264
rect 880 77720 439120 78000
rect 800 77456 439200 77720
rect 880 77176 439120 77456
rect 800 76912 439200 77176
rect 880 76632 439120 76912
rect 800 76368 439200 76632
rect 880 76088 439120 76368
rect 800 75824 439200 76088
rect 880 75544 439120 75824
rect 800 75280 439200 75544
rect 880 75000 439120 75280
rect 800 74736 439200 75000
rect 880 74456 439120 74736
rect 800 74192 439200 74456
rect 880 73912 439120 74192
rect 800 73648 439200 73912
rect 880 73368 439120 73648
rect 800 73104 439200 73368
rect 880 72824 439120 73104
rect 800 72560 439200 72824
rect 880 72280 439120 72560
rect 800 72016 439200 72280
rect 880 71736 439120 72016
rect 800 71472 439200 71736
rect 880 71192 439120 71472
rect 800 70928 439200 71192
rect 880 70648 439120 70928
rect 800 70384 439200 70648
rect 880 70104 439120 70384
rect 800 69840 439200 70104
rect 880 69560 439120 69840
rect 800 69296 439200 69560
rect 880 69016 439120 69296
rect 800 68752 439200 69016
rect 880 68472 439120 68752
rect 800 68208 439200 68472
rect 880 67928 439120 68208
rect 800 67664 439200 67928
rect 880 67384 439120 67664
rect 800 67120 439200 67384
rect 880 66840 439120 67120
rect 800 66576 439200 66840
rect 880 66296 439120 66576
rect 800 66032 439200 66296
rect 880 65752 439120 66032
rect 800 65488 439200 65752
rect 880 65208 439120 65488
rect 800 64944 439200 65208
rect 880 64664 439120 64944
rect 800 64400 439200 64664
rect 880 64120 439120 64400
rect 800 63856 439200 64120
rect 880 63576 439120 63856
rect 800 63312 439200 63576
rect 880 63032 439120 63312
rect 800 62768 439200 63032
rect 880 62488 439120 62768
rect 800 62224 439200 62488
rect 880 61944 439120 62224
rect 800 61680 439200 61944
rect 880 61400 439120 61680
rect 800 61136 439200 61400
rect 880 60856 439120 61136
rect 800 60592 439200 60856
rect 880 60312 439120 60592
rect 800 60048 439200 60312
rect 880 59768 439120 60048
rect 800 59504 439200 59768
rect 880 59224 439120 59504
rect 800 58960 439200 59224
rect 880 58680 439120 58960
rect 800 58416 439200 58680
rect 880 58136 439120 58416
rect 800 57872 439200 58136
rect 880 57592 439120 57872
rect 800 57328 439200 57592
rect 880 57048 439120 57328
rect 800 56784 439200 57048
rect 880 56504 439120 56784
rect 800 56240 439200 56504
rect 880 55960 439120 56240
rect 800 55696 439200 55960
rect 880 55416 439120 55696
rect 800 55152 439200 55416
rect 880 54872 439120 55152
rect 800 54608 439200 54872
rect 880 54328 439120 54608
rect 800 54064 439200 54328
rect 880 53784 439120 54064
rect 800 53520 439200 53784
rect 880 53240 439120 53520
rect 800 52976 439200 53240
rect 880 52696 439120 52976
rect 800 52432 439200 52696
rect 880 52152 439120 52432
rect 800 51888 439200 52152
rect 880 51608 439120 51888
rect 800 51344 439200 51608
rect 880 51064 439120 51344
rect 800 50800 439200 51064
rect 880 50520 439120 50800
rect 800 50256 439200 50520
rect 880 49976 439120 50256
rect 800 49712 439200 49976
rect 880 49432 439120 49712
rect 800 49168 439200 49432
rect 880 48888 439120 49168
rect 800 48624 439200 48888
rect 880 48344 439120 48624
rect 800 48080 439200 48344
rect 880 47800 439120 48080
rect 800 47536 439200 47800
rect 880 47256 439120 47536
rect 800 46992 439200 47256
rect 880 46712 439120 46992
rect 800 46448 439200 46712
rect 880 46168 439120 46448
rect 800 45904 439200 46168
rect 880 45624 439120 45904
rect 800 45360 439200 45624
rect 880 45080 439120 45360
rect 800 44816 439200 45080
rect 880 44536 439120 44816
rect 800 44272 439200 44536
rect 880 43992 439120 44272
rect 800 43728 439200 43992
rect 880 43448 439120 43728
rect 800 43184 439200 43448
rect 880 42904 439120 43184
rect 800 42640 439200 42904
rect 880 42360 439120 42640
rect 800 42096 439200 42360
rect 880 41816 439120 42096
rect 800 41552 439200 41816
rect 880 41272 439120 41552
rect 800 41008 439200 41272
rect 880 40728 439120 41008
rect 800 40464 439200 40728
rect 880 40184 439120 40464
rect 800 39920 439200 40184
rect 880 39640 439120 39920
rect 800 39376 439200 39640
rect 880 39096 439120 39376
rect 800 38832 439200 39096
rect 880 38552 439120 38832
rect 800 38288 439200 38552
rect 880 38008 439120 38288
rect 800 37744 439200 38008
rect 880 37464 439120 37744
rect 800 37200 439200 37464
rect 880 36920 439120 37200
rect 800 36656 439200 36920
rect 880 36376 439120 36656
rect 800 36112 439200 36376
rect 880 35832 439120 36112
rect 800 35568 439200 35832
rect 880 35288 439120 35568
rect 800 35024 439200 35288
rect 880 34744 439120 35024
rect 800 34480 439200 34744
rect 880 34200 439120 34480
rect 800 33936 439200 34200
rect 880 33656 439120 33936
rect 800 33392 439200 33656
rect 880 33112 439120 33392
rect 800 32848 439200 33112
rect 880 32568 439120 32848
rect 800 32304 439200 32568
rect 880 32024 439120 32304
rect 800 31760 439200 32024
rect 880 31480 439120 31760
rect 800 31216 439200 31480
rect 880 30936 439120 31216
rect 800 30672 439200 30936
rect 880 30392 439120 30672
rect 800 30128 439200 30392
rect 880 29848 439120 30128
rect 800 29584 439200 29848
rect 880 29304 439120 29584
rect 800 29040 439200 29304
rect 880 28760 439120 29040
rect 800 28496 439200 28760
rect 880 28216 439120 28496
rect 800 27952 439200 28216
rect 880 27672 439120 27952
rect 800 27408 439200 27672
rect 880 27128 439120 27408
rect 800 26864 439200 27128
rect 880 26584 439120 26864
rect 800 26320 439200 26584
rect 880 26040 439120 26320
rect 800 25776 439200 26040
rect 880 25496 439120 25776
rect 800 25232 439200 25496
rect 880 24952 439120 25232
rect 800 24688 439200 24952
rect 880 24408 439120 24688
rect 800 24144 439200 24408
rect 880 23864 439120 24144
rect 800 23600 439200 23864
rect 880 23320 439120 23600
rect 800 23056 439200 23320
rect 880 22776 439120 23056
rect 800 22512 439200 22776
rect 880 22232 439120 22512
rect 800 21968 439200 22232
rect 880 21688 439120 21968
rect 800 21424 439200 21688
rect 880 21144 439120 21424
rect 800 20880 439200 21144
rect 880 20600 439120 20880
rect 800 20336 439200 20600
rect 880 20056 439120 20336
rect 800 19792 439200 20056
rect 880 19512 439120 19792
rect 800 19248 439200 19512
rect 880 18968 439120 19248
rect 800 18704 439200 18968
rect 880 18424 439120 18704
rect 800 18160 439200 18424
rect 880 17880 439120 18160
rect 800 17616 439200 17880
rect 880 17336 439120 17616
rect 800 17072 439200 17336
rect 880 16792 439120 17072
rect 800 16528 439200 16792
rect 880 16248 439120 16528
rect 800 15984 439200 16248
rect 800 15704 439120 15984
rect 800 15440 439200 15704
rect 800 15160 439120 15440
rect 800 1939 439200 15160
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
rect 127088 2128 127408 157808
rect 142448 2128 142768 157808
rect 157808 2128 158128 157808
rect 173168 2128 173488 157808
rect 188528 2128 188848 157808
rect 203888 2128 204208 157808
rect 219248 2128 219568 157808
rect 234608 2128 234928 157808
rect 249968 2128 250288 157808
rect 265328 2128 265648 157808
rect 280688 2128 281008 157808
rect 296048 2128 296368 157808
rect 311408 2128 311728 157808
rect 326768 2128 327088 157808
rect 342128 2128 342448 157808
rect 357488 2128 357808 157808
rect 372848 2128 373168 157808
rect 388208 2128 388528 157808
rect 403568 2128 403888 157808
rect 418928 2128 419248 157808
rect 434288 2128 434608 157808
<< obsm4 >>
rect 3371 157888 437309 159357
rect 3371 3027 4128 157888
rect 4608 3027 19488 157888
rect 19968 3027 34848 157888
rect 35328 3027 50208 157888
rect 50688 3027 65568 157888
rect 66048 3027 80928 157888
rect 81408 3027 96288 157888
rect 96768 3027 111648 157888
rect 112128 3027 127008 157888
rect 127488 3027 142368 157888
rect 142848 3027 157728 157888
rect 158208 3027 173088 157888
rect 173568 3027 188448 157888
rect 188928 3027 203808 157888
rect 204288 3027 219168 157888
rect 219648 3027 234528 157888
rect 235008 3027 249888 157888
rect 250368 3027 265248 157888
rect 265728 3027 280608 157888
rect 281088 3027 295968 157888
rect 296448 3027 311328 157888
rect 311808 3027 326688 157888
rect 327168 3027 342048 157888
rect 342528 3027 357408 157888
rect 357888 3027 372768 157888
rect 373248 3027 388128 157888
rect 388608 3027 403488 157888
rect 403968 3027 418848 157888
rect 419328 3027 434208 157888
rect 434688 3027 437309 157888
<< labels >>
rlabel metal2 s 8390 159200 8446 160000 6 cache_PC[0]
port 1 nsew signal output
rlabel metal2 s 18510 159200 18566 160000 6 cache_PC[10]
port 2 nsew signal output
rlabel metal2 s 19522 159200 19578 160000 6 cache_PC[11]
port 3 nsew signal output
rlabel metal2 s 20534 159200 20590 160000 6 cache_PC[12]
port 4 nsew signal output
rlabel metal2 s 21546 159200 21602 160000 6 cache_PC[13]
port 5 nsew signal output
rlabel metal2 s 22558 159200 22614 160000 6 cache_PC[14]
port 6 nsew signal output
rlabel metal2 s 23570 159200 23626 160000 6 cache_PC[15]
port 7 nsew signal output
rlabel metal2 s 24582 159200 24638 160000 6 cache_PC[16]
port 8 nsew signal output
rlabel metal2 s 25594 159200 25650 160000 6 cache_PC[17]
port 9 nsew signal output
rlabel metal2 s 26606 159200 26662 160000 6 cache_PC[18]
port 10 nsew signal output
rlabel metal2 s 27618 159200 27674 160000 6 cache_PC[19]
port 11 nsew signal output
rlabel metal2 s 9402 159200 9458 160000 6 cache_PC[1]
port 12 nsew signal output
rlabel metal2 s 28630 159200 28686 160000 6 cache_PC[20]
port 13 nsew signal output
rlabel metal2 s 29642 159200 29698 160000 6 cache_PC[21]
port 14 nsew signal output
rlabel metal2 s 30654 159200 30710 160000 6 cache_PC[22]
port 15 nsew signal output
rlabel metal2 s 31666 159200 31722 160000 6 cache_PC[23]
port 16 nsew signal output
rlabel metal2 s 32678 159200 32734 160000 6 cache_PC[24]
port 17 nsew signal output
rlabel metal2 s 33690 159200 33746 160000 6 cache_PC[25]
port 18 nsew signal output
rlabel metal2 s 34702 159200 34758 160000 6 cache_PC[26]
port 19 nsew signal output
rlabel metal2 s 35714 159200 35770 160000 6 cache_PC[27]
port 20 nsew signal output
rlabel metal2 s 10414 159200 10470 160000 6 cache_PC[2]
port 21 nsew signal output
rlabel metal2 s 11426 159200 11482 160000 6 cache_PC[3]
port 22 nsew signal output
rlabel metal2 s 12438 159200 12494 160000 6 cache_PC[4]
port 23 nsew signal output
rlabel metal2 s 13450 159200 13506 160000 6 cache_PC[5]
port 24 nsew signal output
rlabel metal2 s 14462 159200 14518 160000 6 cache_PC[6]
port 25 nsew signal output
rlabel metal2 s 15474 159200 15530 160000 6 cache_PC[7]
port 26 nsew signal output
rlabel metal2 s 16486 159200 16542 160000 6 cache_PC[8]
port 27 nsew signal output
rlabel metal2 s 17498 159200 17554 160000 6 cache_PC[9]
port 28 nsew signal output
rlabel metal2 s 36726 159200 36782 160000 6 cache_entry[0]
port 29 nsew signal input
rlabel metal2 s 137926 159200 137982 160000 6 cache_entry[100]
port 30 nsew signal input
rlabel metal2 s 138938 159200 138994 160000 6 cache_entry[101]
port 31 nsew signal input
rlabel metal2 s 139950 159200 140006 160000 6 cache_entry[102]
port 32 nsew signal input
rlabel metal2 s 140962 159200 141018 160000 6 cache_entry[103]
port 33 nsew signal input
rlabel metal2 s 141974 159200 142030 160000 6 cache_entry[104]
port 34 nsew signal input
rlabel metal2 s 142986 159200 143042 160000 6 cache_entry[105]
port 35 nsew signal input
rlabel metal2 s 143998 159200 144054 160000 6 cache_entry[106]
port 36 nsew signal input
rlabel metal2 s 145010 159200 145066 160000 6 cache_entry[107]
port 37 nsew signal input
rlabel metal2 s 146022 159200 146078 160000 6 cache_entry[108]
port 38 nsew signal input
rlabel metal2 s 147034 159200 147090 160000 6 cache_entry[109]
port 39 nsew signal input
rlabel metal2 s 46846 159200 46902 160000 6 cache_entry[10]
port 40 nsew signal input
rlabel metal2 s 148046 159200 148102 160000 6 cache_entry[110]
port 41 nsew signal input
rlabel metal2 s 149058 159200 149114 160000 6 cache_entry[111]
port 42 nsew signal input
rlabel metal2 s 150070 159200 150126 160000 6 cache_entry[112]
port 43 nsew signal input
rlabel metal2 s 151082 159200 151138 160000 6 cache_entry[113]
port 44 nsew signal input
rlabel metal2 s 152094 159200 152150 160000 6 cache_entry[114]
port 45 nsew signal input
rlabel metal2 s 153106 159200 153162 160000 6 cache_entry[115]
port 46 nsew signal input
rlabel metal2 s 154118 159200 154174 160000 6 cache_entry[116]
port 47 nsew signal input
rlabel metal2 s 155130 159200 155186 160000 6 cache_entry[117]
port 48 nsew signal input
rlabel metal2 s 156142 159200 156198 160000 6 cache_entry[118]
port 49 nsew signal input
rlabel metal2 s 157154 159200 157210 160000 6 cache_entry[119]
port 50 nsew signal input
rlabel metal2 s 47858 159200 47914 160000 6 cache_entry[11]
port 51 nsew signal input
rlabel metal2 s 158166 159200 158222 160000 6 cache_entry[120]
port 52 nsew signal input
rlabel metal2 s 159178 159200 159234 160000 6 cache_entry[121]
port 53 nsew signal input
rlabel metal2 s 160190 159200 160246 160000 6 cache_entry[122]
port 54 nsew signal input
rlabel metal2 s 161202 159200 161258 160000 6 cache_entry[123]
port 55 nsew signal input
rlabel metal2 s 162214 159200 162270 160000 6 cache_entry[124]
port 56 nsew signal input
rlabel metal2 s 163226 159200 163282 160000 6 cache_entry[125]
port 57 nsew signal input
rlabel metal2 s 164238 159200 164294 160000 6 cache_entry[126]
port 58 nsew signal input
rlabel metal2 s 165250 159200 165306 160000 6 cache_entry[127]
port 59 nsew signal input
rlabel metal2 s 48870 159200 48926 160000 6 cache_entry[12]
port 60 nsew signal input
rlabel metal2 s 49882 159200 49938 160000 6 cache_entry[13]
port 61 nsew signal input
rlabel metal2 s 50894 159200 50950 160000 6 cache_entry[14]
port 62 nsew signal input
rlabel metal2 s 51906 159200 51962 160000 6 cache_entry[15]
port 63 nsew signal input
rlabel metal2 s 52918 159200 52974 160000 6 cache_entry[16]
port 64 nsew signal input
rlabel metal2 s 53930 159200 53986 160000 6 cache_entry[17]
port 65 nsew signal input
rlabel metal2 s 54942 159200 54998 160000 6 cache_entry[18]
port 66 nsew signal input
rlabel metal2 s 55954 159200 56010 160000 6 cache_entry[19]
port 67 nsew signal input
rlabel metal2 s 37738 159200 37794 160000 6 cache_entry[1]
port 68 nsew signal input
rlabel metal2 s 56966 159200 57022 160000 6 cache_entry[20]
port 69 nsew signal input
rlabel metal2 s 57978 159200 58034 160000 6 cache_entry[21]
port 70 nsew signal input
rlabel metal2 s 58990 159200 59046 160000 6 cache_entry[22]
port 71 nsew signal input
rlabel metal2 s 60002 159200 60058 160000 6 cache_entry[23]
port 72 nsew signal input
rlabel metal2 s 61014 159200 61070 160000 6 cache_entry[24]
port 73 nsew signal input
rlabel metal2 s 62026 159200 62082 160000 6 cache_entry[25]
port 74 nsew signal input
rlabel metal2 s 63038 159200 63094 160000 6 cache_entry[26]
port 75 nsew signal input
rlabel metal2 s 64050 159200 64106 160000 6 cache_entry[27]
port 76 nsew signal input
rlabel metal2 s 65062 159200 65118 160000 6 cache_entry[28]
port 77 nsew signal input
rlabel metal2 s 66074 159200 66130 160000 6 cache_entry[29]
port 78 nsew signal input
rlabel metal2 s 38750 159200 38806 160000 6 cache_entry[2]
port 79 nsew signal input
rlabel metal2 s 67086 159200 67142 160000 6 cache_entry[30]
port 80 nsew signal input
rlabel metal2 s 68098 159200 68154 160000 6 cache_entry[31]
port 81 nsew signal input
rlabel metal2 s 69110 159200 69166 160000 6 cache_entry[32]
port 82 nsew signal input
rlabel metal2 s 70122 159200 70178 160000 6 cache_entry[33]
port 83 nsew signal input
rlabel metal2 s 71134 159200 71190 160000 6 cache_entry[34]
port 84 nsew signal input
rlabel metal2 s 72146 159200 72202 160000 6 cache_entry[35]
port 85 nsew signal input
rlabel metal2 s 73158 159200 73214 160000 6 cache_entry[36]
port 86 nsew signal input
rlabel metal2 s 74170 159200 74226 160000 6 cache_entry[37]
port 87 nsew signal input
rlabel metal2 s 75182 159200 75238 160000 6 cache_entry[38]
port 88 nsew signal input
rlabel metal2 s 76194 159200 76250 160000 6 cache_entry[39]
port 89 nsew signal input
rlabel metal2 s 39762 159200 39818 160000 6 cache_entry[3]
port 90 nsew signal input
rlabel metal2 s 77206 159200 77262 160000 6 cache_entry[40]
port 91 nsew signal input
rlabel metal2 s 78218 159200 78274 160000 6 cache_entry[41]
port 92 nsew signal input
rlabel metal2 s 79230 159200 79286 160000 6 cache_entry[42]
port 93 nsew signal input
rlabel metal2 s 80242 159200 80298 160000 6 cache_entry[43]
port 94 nsew signal input
rlabel metal2 s 81254 159200 81310 160000 6 cache_entry[44]
port 95 nsew signal input
rlabel metal2 s 82266 159200 82322 160000 6 cache_entry[45]
port 96 nsew signal input
rlabel metal2 s 83278 159200 83334 160000 6 cache_entry[46]
port 97 nsew signal input
rlabel metal2 s 84290 159200 84346 160000 6 cache_entry[47]
port 98 nsew signal input
rlabel metal2 s 85302 159200 85358 160000 6 cache_entry[48]
port 99 nsew signal input
rlabel metal2 s 86314 159200 86370 160000 6 cache_entry[49]
port 100 nsew signal input
rlabel metal2 s 40774 159200 40830 160000 6 cache_entry[4]
port 101 nsew signal input
rlabel metal2 s 87326 159200 87382 160000 6 cache_entry[50]
port 102 nsew signal input
rlabel metal2 s 88338 159200 88394 160000 6 cache_entry[51]
port 103 nsew signal input
rlabel metal2 s 89350 159200 89406 160000 6 cache_entry[52]
port 104 nsew signal input
rlabel metal2 s 90362 159200 90418 160000 6 cache_entry[53]
port 105 nsew signal input
rlabel metal2 s 91374 159200 91430 160000 6 cache_entry[54]
port 106 nsew signal input
rlabel metal2 s 92386 159200 92442 160000 6 cache_entry[55]
port 107 nsew signal input
rlabel metal2 s 93398 159200 93454 160000 6 cache_entry[56]
port 108 nsew signal input
rlabel metal2 s 94410 159200 94466 160000 6 cache_entry[57]
port 109 nsew signal input
rlabel metal2 s 95422 159200 95478 160000 6 cache_entry[58]
port 110 nsew signal input
rlabel metal2 s 96434 159200 96490 160000 6 cache_entry[59]
port 111 nsew signal input
rlabel metal2 s 41786 159200 41842 160000 6 cache_entry[5]
port 112 nsew signal input
rlabel metal2 s 97446 159200 97502 160000 6 cache_entry[60]
port 113 nsew signal input
rlabel metal2 s 98458 159200 98514 160000 6 cache_entry[61]
port 114 nsew signal input
rlabel metal2 s 99470 159200 99526 160000 6 cache_entry[62]
port 115 nsew signal input
rlabel metal2 s 100482 159200 100538 160000 6 cache_entry[63]
port 116 nsew signal input
rlabel metal2 s 101494 159200 101550 160000 6 cache_entry[64]
port 117 nsew signal input
rlabel metal2 s 102506 159200 102562 160000 6 cache_entry[65]
port 118 nsew signal input
rlabel metal2 s 103518 159200 103574 160000 6 cache_entry[66]
port 119 nsew signal input
rlabel metal2 s 104530 159200 104586 160000 6 cache_entry[67]
port 120 nsew signal input
rlabel metal2 s 105542 159200 105598 160000 6 cache_entry[68]
port 121 nsew signal input
rlabel metal2 s 106554 159200 106610 160000 6 cache_entry[69]
port 122 nsew signal input
rlabel metal2 s 42798 159200 42854 160000 6 cache_entry[6]
port 123 nsew signal input
rlabel metal2 s 107566 159200 107622 160000 6 cache_entry[70]
port 124 nsew signal input
rlabel metal2 s 108578 159200 108634 160000 6 cache_entry[71]
port 125 nsew signal input
rlabel metal2 s 109590 159200 109646 160000 6 cache_entry[72]
port 126 nsew signal input
rlabel metal2 s 110602 159200 110658 160000 6 cache_entry[73]
port 127 nsew signal input
rlabel metal2 s 111614 159200 111670 160000 6 cache_entry[74]
port 128 nsew signal input
rlabel metal2 s 112626 159200 112682 160000 6 cache_entry[75]
port 129 nsew signal input
rlabel metal2 s 113638 159200 113694 160000 6 cache_entry[76]
port 130 nsew signal input
rlabel metal2 s 114650 159200 114706 160000 6 cache_entry[77]
port 131 nsew signal input
rlabel metal2 s 115662 159200 115718 160000 6 cache_entry[78]
port 132 nsew signal input
rlabel metal2 s 116674 159200 116730 160000 6 cache_entry[79]
port 133 nsew signal input
rlabel metal2 s 43810 159200 43866 160000 6 cache_entry[7]
port 134 nsew signal input
rlabel metal2 s 117686 159200 117742 160000 6 cache_entry[80]
port 135 nsew signal input
rlabel metal2 s 118698 159200 118754 160000 6 cache_entry[81]
port 136 nsew signal input
rlabel metal2 s 119710 159200 119766 160000 6 cache_entry[82]
port 137 nsew signal input
rlabel metal2 s 120722 159200 120778 160000 6 cache_entry[83]
port 138 nsew signal input
rlabel metal2 s 121734 159200 121790 160000 6 cache_entry[84]
port 139 nsew signal input
rlabel metal2 s 122746 159200 122802 160000 6 cache_entry[85]
port 140 nsew signal input
rlabel metal2 s 123758 159200 123814 160000 6 cache_entry[86]
port 141 nsew signal input
rlabel metal2 s 124770 159200 124826 160000 6 cache_entry[87]
port 142 nsew signal input
rlabel metal2 s 125782 159200 125838 160000 6 cache_entry[88]
port 143 nsew signal input
rlabel metal2 s 126794 159200 126850 160000 6 cache_entry[89]
port 144 nsew signal input
rlabel metal2 s 44822 159200 44878 160000 6 cache_entry[8]
port 145 nsew signal input
rlabel metal2 s 127806 159200 127862 160000 6 cache_entry[90]
port 146 nsew signal input
rlabel metal2 s 128818 159200 128874 160000 6 cache_entry[91]
port 147 nsew signal input
rlabel metal2 s 129830 159200 129886 160000 6 cache_entry[92]
port 148 nsew signal input
rlabel metal2 s 130842 159200 130898 160000 6 cache_entry[93]
port 149 nsew signal input
rlabel metal2 s 131854 159200 131910 160000 6 cache_entry[94]
port 150 nsew signal input
rlabel metal2 s 132866 159200 132922 160000 6 cache_entry[95]
port 151 nsew signal input
rlabel metal2 s 133878 159200 133934 160000 6 cache_entry[96]
port 152 nsew signal input
rlabel metal2 s 134890 159200 134946 160000 6 cache_entry[97]
port 153 nsew signal input
rlabel metal2 s 135902 159200 135958 160000 6 cache_entry[98]
port 154 nsew signal input
rlabel metal2 s 136914 159200 136970 160000 6 cache_entry[99]
port 155 nsew signal input
rlabel metal2 s 45834 159200 45890 160000 6 cache_entry[9]
port 156 nsew signal input
rlabel metal3 s 439200 16872 440000 16992 6 cache_entry_valid
port 157 nsew signal output
rlabel metal3 s 439200 15240 440000 15360 6 cache_hit
port 158 nsew signal input
rlabel metal3 s 439200 15784 440000 15904 6 cache_invalidate
port 159 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 cache_new_entry[0]
port 160 nsew signal output
rlabel metal2 s 183190 0 183246 800 6 cache_new_entry[100]
port 161 nsew signal output
rlabel metal2 s 184938 0 184994 800 6 cache_new_entry[101]
port 162 nsew signal output
rlabel metal2 s 186686 0 186742 800 6 cache_new_entry[102]
port 163 nsew signal output
rlabel metal2 s 188434 0 188490 800 6 cache_new_entry[103]
port 164 nsew signal output
rlabel metal2 s 190182 0 190238 800 6 cache_new_entry[104]
port 165 nsew signal output
rlabel metal2 s 191930 0 191986 800 6 cache_new_entry[105]
port 166 nsew signal output
rlabel metal2 s 193678 0 193734 800 6 cache_new_entry[106]
port 167 nsew signal output
rlabel metal2 s 195426 0 195482 800 6 cache_new_entry[107]
port 168 nsew signal output
rlabel metal2 s 197174 0 197230 800 6 cache_new_entry[108]
port 169 nsew signal output
rlabel metal2 s 198922 0 198978 800 6 cache_new_entry[109]
port 170 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 cache_new_entry[10]
port 171 nsew signal output
rlabel metal2 s 200670 0 200726 800 6 cache_new_entry[110]
port 172 nsew signal output
rlabel metal2 s 202418 0 202474 800 6 cache_new_entry[111]
port 173 nsew signal output
rlabel metal2 s 204166 0 204222 800 6 cache_new_entry[112]
port 174 nsew signal output
rlabel metal2 s 205914 0 205970 800 6 cache_new_entry[113]
port 175 nsew signal output
rlabel metal2 s 207662 0 207718 800 6 cache_new_entry[114]
port 176 nsew signal output
rlabel metal2 s 209410 0 209466 800 6 cache_new_entry[115]
port 177 nsew signal output
rlabel metal2 s 211158 0 211214 800 6 cache_new_entry[116]
port 178 nsew signal output
rlabel metal2 s 212906 0 212962 800 6 cache_new_entry[117]
port 179 nsew signal output
rlabel metal2 s 214654 0 214710 800 6 cache_new_entry[118]
port 180 nsew signal output
rlabel metal2 s 216402 0 216458 800 6 cache_new_entry[119]
port 181 nsew signal output
rlabel metal2 s 27618 0 27674 800 6 cache_new_entry[11]
port 182 nsew signal output
rlabel metal2 s 218150 0 218206 800 6 cache_new_entry[120]
port 183 nsew signal output
rlabel metal2 s 219898 0 219954 800 6 cache_new_entry[121]
port 184 nsew signal output
rlabel metal2 s 221646 0 221702 800 6 cache_new_entry[122]
port 185 nsew signal output
rlabel metal2 s 223394 0 223450 800 6 cache_new_entry[123]
port 186 nsew signal output
rlabel metal2 s 225142 0 225198 800 6 cache_new_entry[124]
port 187 nsew signal output
rlabel metal2 s 226890 0 226946 800 6 cache_new_entry[125]
port 188 nsew signal output
rlabel metal2 s 228638 0 228694 800 6 cache_new_entry[126]
port 189 nsew signal output
rlabel metal2 s 230386 0 230442 800 6 cache_new_entry[127]
port 190 nsew signal output
rlabel metal2 s 29366 0 29422 800 6 cache_new_entry[12]
port 191 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 cache_new_entry[13]
port 192 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 cache_new_entry[14]
port 193 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 cache_new_entry[15]
port 194 nsew signal output
rlabel metal2 s 36358 0 36414 800 6 cache_new_entry[16]
port 195 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 cache_new_entry[17]
port 196 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 cache_new_entry[18]
port 197 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 cache_new_entry[19]
port 198 nsew signal output
rlabel metal2 s 10138 0 10194 800 6 cache_new_entry[1]
port 199 nsew signal output
rlabel metal2 s 43350 0 43406 800 6 cache_new_entry[20]
port 200 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 cache_new_entry[21]
port 201 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 cache_new_entry[22]
port 202 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 cache_new_entry[23]
port 203 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 cache_new_entry[24]
port 204 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 cache_new_entry[25]
port 205 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 cache_new_entry[26]
port 206 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 cache_new_entry[27]
port 207 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 cache_new_entry[28]
port 208 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 cache_new_entry[29]
port 209 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 cache_new_entry[2]
port 210 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 cache_new_entry[30]
port 211 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 cache_new_entry[31]
port 212 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 cache_new_entry[32]
port 213 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 cache_new_entry[33]
port 214 nsew signal output
rlabel metal2 s 67822 0 67878 800 6 cache_new_entry[34]
port 215 nsew signal output
rlabel metal2 s 69570 0 69626 800 6 cache_new_entry[35]
port 216 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 cache_new_entry[36]
port 217 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 cache_new_entry[37]
port 218 nsew signal output
rlabel metal2 s 74814 0 74870 800 6 cache_new_entry[38]
port 219 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 cache_new_entry[39]
port 220 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 cache_new_entry[3]
port 221 nsew signal output
rlabel metal2 s 78310 0 78366 800 6 cache_new_entry[40]
port 222 nsew signal output
rlabel metal2 s 80058 0 80114 800 6 cache_new_entry[41]
port 223 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 cache_new_entry[42]
port 224 nsew signal output
rlabel metal2 s 83554 0 83610 800 6 cache_new_entry[43]
port 225 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 cache_new_entry[44]
port 226 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 cache_new_entry[45]
port 227 nsew signal output
rlabel metal2 s 88798 0 88854 800 6 cache_new_entry[46]
port 228 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 cache_new_entry[47]
port 229 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 cache_new_entry[48]
port 230 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 cache_new_entry[49]
port 231 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 cache_new_entry[4]
port 232 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 cache_new_entry[50]
port 233 nsew signal output
rlabel metal2 s 97538 0 97594 800 6 cache_new_entry[51]
port 234 nsew signal output
rlabel metal2 s 99286 0 99342 800 6 cache_new_entry[52]
port 235 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 cache_new_entry[53]
port 236 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 cache_new_entry[54]
port 237 nsew signal output
rlabel metal2 s 104530 0 104586 800 6 cache_new_entry[55]
port 238 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 cache_new_entry[56]
port 239 nsew signal output
rlabel metal2 s 108026 0 108082 800 6 cache_new_entry[57]
port 240 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 cache_new_entry[58]
port 241 nsew signal output
rlabel metal2 s 111522 0 111578 800 6 cache_new_entry[59]
port 242 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 cache_new_entry[5]
port 243 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 cache_new_entry[60]
port 244 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 cache_new_entry[61]
port 245 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 cache_new_entry[62]
port 246 nsew signal output
rlabel metal2 s 118514 0 118570 800 6 cache_new_entry[63]
port 247 nsew signal output
rlabel metal2 s 120262 0 120318 800 6 cache_new_entry[64]
port 248 nsew signal output
rlabel metal2 s 122010 0 122066 800 6 cache_new_entry[65]
port 249 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 cache_new_entry[66]
port 250 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 cache_new_entry[67]
port 251 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 cache_new_entry[68]
port 252 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 cache_new_entry[69]
port 253 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 cache_new_entry[6]
port 254 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 cache_new_entry[70]
port 255 nsew signal output
rlabel metal2 s 132498 0 132554 800 6 cache_new_entry[71]
port 256 nsew signal output
rlabel metal2 s 134246 0 134302 800 6 cache_new_entry[72]
port 257 nsew signal output
rlabel metal2 s 135994 0 136050 800 6 cache_new_entry[73]
port 258 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 cache_new_entry[74]
port 259 nsew signal output
rlabel metal2 s 139490 0 139546 800 6 cache_new_entry[75]
port 260 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 cache_new_entry[76]
port 261 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 cache_new_entry[77]
port 262 nsew signal output
rlabel metal2 s 144734 0 144790 800 6 cache_new_entry[78]
port 263 nsew signal output
rlabel metal2 s 146482 0 146538 800 6 cache_new_entry[79]
port 264 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 cache_new_entry[7]
port 265 nsew signal output
rlabel metal2 s 148230 0 148286 800 6 cache_new_entry[80]
port 266 nsew signal output
rlabel metal2 s 149978 0 150034 800 6 cache_new_entry[81]
port 267 nsew signal output
rlabel metal2 s 151726 0 151782 800 6 cache_new_entry[82]
port 268 nsew signal output
rlabel metal2 s 153474 0 153530 800 6 cache_new_entry[83]
port 269 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 cache_new_entry[84]
port 270 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 cache_new_entry[85]
port 271 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 cache_new_entry[86]
port 272 nsew signal output
rlabel metal2 s 160466 0 160522 800 6 cache_new_entry[87]
port 273 nsew signal output
rlabel metal2 s 162214 0 162270 800 6 cache_new_entry[88]
port 274 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 cache_new_entry[89]
port 275 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 cache_new_entry[8]
port 276 nsew signal output
rlabel metal2 s 165710 0 165766 800 6 cache_new_entry[90]
port 277 nsew signal output
rlabel metal2 s 167458 0 167514 800 6 cache_new_entry[91]
port 278 nsew signal output
rlabel metal2 s 169206 0 169262 800 6 cache_new_entry[92]
port 279 nsew signal output
rlabel metal2 s 170954 0 171010 800 6 cache_new_entry[93]
port 280 nsew signal output
rlabel metal2 s 172702 0 172758 800 6 cache_new_entry[94]
port 281 nsew signal output
rlabel metal2 s 174450 0 174506 800 6 cache_new_entry[95]
port 282 nsew signal output
rlabel metal2 s 176198 0 176254 800 6 cache_new_entry[96]
port 283 nsew signal output
rlabel metal2 s 177946 0 178002 800 6 cache_new_entry[97]
port 284 nsew signal output
rlabel metal2 s 179694 0 179750 800 6 cache_new_entry[98]
port 285 nsew signal output
rlabel metal2 s 181442 0 181498 800 6 cache_new_entry[99]
port 286 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 cache_new_entry[9]
port 287 nsew signal output
rlabel metal3 s 439200 16328 440000 16448 6 cache_rst
port 288 nsew signal output
rlabel metal2 s 167274 159200 167330 160000 6 curr_PC[0]
port 289 nsew signal output
rlabel metal2 s 177394 159200 177450 160000 6 curr_PC[10]
port 290 nsew signal output
rlabel metal2 s 178406 159200 178462 160000 6 curr_PC[11]
port 291 nsew signal output
rlabel metal2 s 179418 159200 179474 160000 6 curr_PC[12]
port 292 nsew signal output
rlabel metal2 s 180430 159200 180486 160000 6 curr_PC[13]
port 293 nsew signal output
rlabel metal2 s 181442 159200 181498 160000 6 curr_PC[14]
port 294 nsew signal output
rlabel metal2 s 182454 159200 182510 160000 6 curr_PC[15]
port 295 nsew signal output
rlabel metal2 s 183466 159200 183522 160000 6 curr_PC[16]
port 296 nsew signal output
rlabel metal2 s 184478 159200 184534 160000 6 curr_PC[17]
port 297 nsew signal output
rlabel metal2 s 185490 159200 185546 160000 6 curr_PC[18]
port 298 nsew signal output
rlabel metal2 s 186502 159200 186558 160000 6 curr_PC[19]
port 299 nsew signal output
rlabel metal2 s 168286 159200 168342 160000 6 curr_PC[1]
port 300 nsew signal output
rlabel metal2 s 187514 159200 187570 160000 6 curr_PC[20]
port 301 nsew signal output
rlabel metal2 s 188526 159200 188582 160000 6 curr_PC[21]
port 302 nsew signal output
rlabel metal2 s 189538 159200 189594 160000 6 curr_PC[22]
port 303 nsew signal output
rlabel metal2 s 190550 159200 190606 160000 6 curr_PC[23]
port 304 nsew signal output
rlabel metal2 s 191562 159200 191618 160000 6 curr_PC[24]
port 305 nsew signal output
rlabel metal2 s 192574 159200 192630 160000 6 curr_PC[25]
port 306 nsew signal output
rlabel metal2 s 193586 159200 193642 160000 6 curr_PC[26]
port 307 nsew signal output
rlabel metal2 s 194598 159200 194654 160000 6 curr_PC[27]
port 308 nsew signal output
rlabel metal2 s 169298 159200 169354 160000 6 curr_PC[2]
port 309 nsew signal output
rlabel metal2 s 170310 159200 170366 160000 6 curr_PC[3]
port 310 nsew signal output
rlabel metal2 s 171322 159200 171378 160000 6 curr_PC[4]
port 311 nsew signal output
rlabel metal2 s 172334 159200 172390 160000 6 curr_PC[5]
port 312 nsew signal output
rlabel metal2 s 173346 159200 173402 160000 6 curr_PC[6]
port 313 nsew signal output
rlabel metal2 s 174358 159200 174414 160000 6 curr_PC[7]
port 314 nsew signal output
rlabel metal2 s 175370 159200 175426 160000 6 curr_PC[8]
port 315 nsew signal output
rlabel metal2 s 176382 159200 176438 160000 6 curr_PC[9]
port 316 nsew signal output
rlabel metal2 s 424414 0 424470 800 6 custom_settings[0]
port 317 nsew signal input
rlabel metal2 s 426162 0 426218 800 6 custom_settings[1]
port 318 nsew signal input
rlabel metal2 s 427910 0 427966 800 6 custom_settings[2]
port 319 nsew signal input
rlabel metal2 s 429658 0 429714 800 6 custom_settings[3]
port 320 nsew signal input
rlabel metal2 s 431406 0 431462 800 6 custom_settings[4]
port 321 nsew signal input
rlabel metal2 s 242162 159200 242218 160000 6 dest_idx0[0]
port 322 nsew signal input
rlabel metal2 s 243174 159200 243230 160000 6 dest_idx0[1]
port 323 nsew signal input
rlabel metal2 s 244186 159200 244242 160000 6 dest_idx0[2]
port 324 nsew signal input
rlabel metal2 s 245198 159200 245254 160000 6 dest_idx0[3]
port 325 nsew signal input
rlabel metal2 s 246210 159200 246266 160000 6 dest_idx0[4]
port 326 nsew signal input
rlabel metal2 s 247222 159200 247278 160000 6 dest_idx0[5]
port 327 nsew signal input
rlabel metal3 s 439200 42440 440000 42560 6 dest_idx1[0]
port 328 nsew signal input
rlabel metal3 s 439200 42984 440000 43104 6 dest_idx1[1]
port 329 nsew signal input
rlabel metal3 s 439200 43528 440000 43648 6 dest_idx1[2]
port 330 nsew signal input
rlabel metal3 s 439200 44072 440000 44192 6 dest_idx1[3]
port 331 nsew signal input
rlabel metal3 s 439200 44616 440000 44736 6 dest_idx1[4]
port 332 nsew signal input
rlabel metal3 s 439200 45160 440000 45280 6 dest_idx1[5]
port 333 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 dest_idx2[0]
port 334 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 dest_idx2[1]
port 335 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 dest_idx2[2]
port 336 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 dest_idx2[3]
port 337 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 dest_idx2[4]
port 338 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 dest_idx2[5]
port 339 nsew signal input
rlabel metal2 s 240138 159200 240194 160000 6 dest_mask0[0]
port 340 nsew signal input
rlabel metal2 s 241150 159200 241206 160000 6 dest_mask0[1]
port 341 nsew signal input
rlabel metal3 s 439200 41352 440000 41472 6 dest_mask1[0]
port 342 nsew signal input
rlabel metal3 s 439200 41896 440000 42016 6 dest_mask1[1]
port 343 nsew signal input
rlabel metal3 s 0 40264 800 40384 6 dest_mask2[0]
port 344 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 dest_mask2[1]
port 345 nsew signal input
rlabel metal2 s 251270 159200 251326 160000 6 dest_pred0[0]
port 346 nsew signal input
rlabel metal2 s 252282 159200 252338 160000 6 dest_pred0[1]
port 347 nsew signal input
rlabel metal2 s 253294 159200 253350 160000 6 dest_pred0[2]
port 348 nsew signal input
rlabel metal3 s 439200 47336 440000 47456 6 dest_pred1[0]
port 349 nsew signal input
rlabel metal3 s 439200 47880 440000 48000 6 dest_pred1[1]
port 350 nsew signal input
rlabel metal3 s 439200 48424 440000 48544 6 dest_pred1[2]
port 351 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 dest_pred2[0]
port 352 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 dest_pred2[1]
port 353 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 dest_pred2[2]
port 354 nsew signal input
rlabel metal2 s 254306 159200 254362 160000 6 dest_pred_val0
port 355 nsew signal input
rlabel metal3 s 439200 48968 440000 49088 6 dest_pred_val1
port 356 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 dest_pred_val2
port 357 nsew signal input
rlabel metal2 s 207754 159200 207810 160000 6 dest_val0[0]
port 358 nsew signal input
rlabel metal2 s 217874 159200 217930 160000 6 dest_val0[10]
port 359 nsew signal input
rlabel metal2 s 218886 159200 218942 160000 6 dest_val0[11]
port 360 nsew signal input
rlabel metal2 s 219898 159200 219954 160000 6 dest_val0[12]
port 361 nsew signal input
rlabel metal2 s 220910 159200 220966 160000 6 dest_val0[13]
port 362 nsew signal input
rlabel metal2 s 221922 159200 221978 160000 6 dest_val0[14]
port 363 nsew signal input
rlabel metal2 s 222934 159200 222990 160000 6 dest_val0[15]
port 364 nsew signal input
rlabel metal2 s 223946 159200 224002 160000 6 dest_val0[16]
port 365 nsew signal input
rlabel metal2 s 224958 159200 225014 160000 6 dest_val0[17]
port 366 nsew signal input
rlabel metal2 s 225970 159200 226026 160000 6 dest_val0[18]
port 367 nsew signal input
rlabel metal2 s 226982 159200 227038 160000 6 dest_val0[19]
port 368 nsew signal input
rlabel metal2 s 208766 159200 208822 160000 6 dest_val0[1]
port 369 nsew signal input
rlabel metal2 s 227994 159200 228050 160000 6 dest_val0[20]
port 370 nsew signal input
rlabel metal2 s 229006 159200 229062 160000 6 dest_val0[21]
port 371 nsew signal input
rlabel metal2 s 230018 159200 230074 160000 6 dest_val0[22]
port 372 nsew signal input
rlabel metal2 s 231030 159200 231086 160000 6 dest_val0[23]
port 373 nsew signal input
rlabel metal2 s 232042 159200 232098 160000 6 dest_val0[24]
port 374 nsew signal input
rlabel metal2 s 233054 159200 233110 160000 6 dest_val0[25]
port 375 nsew signal input
rlabel metal2 s 234066 159200 234122 160000 6 dest_val0[26]
port 376 nsew signal input
rlabel metal2 s 235078 159200 235134 160000 6 dest_val0[27]
port 377 nsew signal input
rlabel metal2 s 236090 159200 236146 160000 6 dest_val0[28]
port 378 nsew signal input
rlabel metal2 s 237102 159200 237158 160000 6 dest_val0[29]
port 379 nsew signal input
rlabel metal2 s 209778 159200 209834 160000 6 dest_val0[2]
port 380 nsew signal input
rlabel metal2 s 238114 159200 238170 160000 6 dest_val0[30]
port 381 nsew signal input
rlabel metal2 s 239126 159200 239182 160000 6 dest_val0[31]
port 382 nsew signal input
rlabel metal2 s 210790 159200 210846 160000 6 dest_val0[3]
port 383 nsew signal input
rlabel metal2 s 211802 159200 211858 160000 6 dest_val0[4]
port 384 nsew signal input
rlabel metal2 s 212814 159200 212870 160000 6 dest_val0[5]
port 385 nsew signal input
rlabel metal2 s 213826 159200 213882 160000 6 dest_val0[6]
port 386 nsew signal input
rlabel metal2 s 214838 159200 214894 160000 6 dest_val0[7]
port 387 nsew signal input
rlabel metal2 s 215850 159200 215906 160000 6 dest_val0[8]
port 388 nsew signal input
rlabel metal2 s 216862 159200 216918 160000 6 dest_val0[9]
port 389 nsew signal input
rlabel metal3 s 439200 23944 440000 24064 6 dest_val1[0]
port 390 nsew signal input
rlabel metal3 s 439200 29384 440000 29504 6 dest_val1[10]
port 391 nsew signal input
rlabel metal3 s 439200 29928 440000 30048 6 dest_val1[11]
port 392 nsew signal input
rlabel metal3 s 439200 30472 440000 30592 6 dest_val1[12]
port 393 nsew signal input
rlabel metal3 s 439200 31016 440000 31136 6 dest_val1[13]
port 394 nsew signal input
rlabel metal3 s 439200 31560 440000 31680 6 dest_val1[14]
port 395 nsew signal input
rlabel metal3 s 439200 32104 440000 32224 6 dest_val1[15]
port 396 nsew signal input
rlabel metal3 s 439200 32648 440000 32768 6 dest_val1[16]
port 397 nsew signal input
rlabel metal3 s 439200 33192 440000 33312 6 dest_val1[17]
port 398 nsew signal input
rlabel metal3 s 439200 33736 440000 33856 6 dest_val1[18]
port 399 nsew signal input
rlabel metal3 s 439200 34280 440000 34400 6 dest_val1[19]
port 400 nsew signal input
rlabel metal3 s 439200 24488 440000 24608 6 dest_val1[1]
port 401 nsew signal input
rlabel metal3 s 439200 34824 440000 34944 6 dest_val1[20]
port 402 nsew signal input
rlabel metal3 s 439200 35368 440000 35488 6 dest_val1[21]
port 403 nsew signal input
rlabel metal3 s 439200 35912 440000 36032 6 dest_val1[22]
port 404 nsew signal input
rlabel metal3 s 439200 36456 440000 36576 6 dest_val1[23]
port 405 nsew signal input
rlabel metal3 s 439200 37000 440000 37120 6 dest_val1[24]
port 406 nsew signal input
rlabel metal3 s 439200 37544 440000 37664 6 dest_val1[25]
port 407 nsew signal input
rlabel metal3 s 439200 38088 440000 38208 6 dest_val1[26]
port 408 nsew signal input
rlabel metal3 s 439200 38632 440000 38752 6 dest_val1[27]
port 409 nsew signal input
rlabel metal3 s 439200 39176 440000 39296 6 dest_val1[28]
port 410 nsew signal input
rlabel metal3 s 439200 39720 440000 39840 6 dest_val1[29]
port 411 nsew signal input
rlabel metal3 s 439200 25032 440000 25152 6 dest_val1[2]
port 412 nsew signal input
rlabel metal3 s 439200 40264 440000 40384 6 dest_val1[30]
port 413 nsew signal input
rlabel metal3 s 439200 40808 440000 40928 6 dest_val1[31]
port 414 nsew signal input
rlabel metal3 s 439200 25576 440000 25696 6 dest_val1[3]
port 415 nsew signal input
rlabel metal3 s 439200 26120 440000 26240 6 dest_val1[4]
port 416 nsew signal input
rlabel metal3 s 439200 26664 440000 26784 6 dest_val1[5]
port 417 nsew signal input
rlabel metal3 s 439200 27208 440000 27328 6 dest_val1[6]
port 418 nsew signal input
rlabel metal3 s 439200 27752 440000 27872 6 dest_val1[7]
port 419 nsew signal input
rlabel metal3 s 439200 28296 440000 28416 6 dest_val1[8]
port 420 nsew signal input
rlabel metal3 s 439200 28840 440000 28960 6 dest_val1[9]
port 421 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 dest_val2[0]
port 422 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 dest_val2[10]
port 423 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 dest_val2[11]
port 424 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 dest_val2[12]
port 425 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 dest_val2[13]
port 426 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 dest_val2[14]
port 427 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 dest_val2[15]
port 428 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 dest_val2[16]
port 429 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 dest_val2[17]
port 430 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 dest_val2[18]
port 431 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 dest_val2[19]
port 432 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 dest_val2[1]
port 433 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 dest_val2[20]
port 434 nsew signal input
rlabel metal3 s 0 34280 800 34400 6 dest_val2[21]
port 435 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 dest_val2[22]
port 436 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 dest_val2[23]
port 437 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 dest_val2[24]
port 438 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 dest_val2[25]
port 439 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 dest_val2[26]
port 440 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 dest_val2[27]
port 441 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 dest_val2[28]
port 442 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 dest_val2[29]
port 443 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 dest_val2[2]
port 444 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 dest_val2[30]
port 445 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 dest_val2[31]
port 446 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 dest_val2[3]
port 447 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 dest_val2[4]
port 448 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 dest_val2[5]
port 449 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 dest_val2[6]
port 450 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 dest_val2[7]
port 451 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 dest_val2[8]
port 452 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 dest_val2[9]
port 453 nsew signal input
rlabel metal2 s 322110 159200 322166 160000 6 eu0_busy
port 454 nsew signal input
rlabel metal2 s 323122 159200 323178 160000 6 eu0_instruction[0]
port 455 nsew signal output
rlabel metal2 s 333242 159200 333298 160000 6 eu0_instruction[10]
port 456 nsew signal output
rlabel metal2 s 334254 159200 334310 160000 6 eu0_instruction[11]
port 457 nsew signal output
rlabel metal2 s 335266 159200 335322 160000 6 eu0_instruction[12]
port 458 nsew signal output
rlabel metal2 s 336278 159200 336334 160000 6 eu0_instruction[13]
port 459 nsew signal output
rlabel metal2 s 337290 159200 337346 160000 6 eu0_instruction[14]
port 460 nsew signal output
rlabel metal2 s 338302 159200 338358 160000 6 eu0_instruction[15]
port 461 nsew signal output
rlabel metal2 s 339314 159200 339370 160000 6 eu0_instruction[16]
port 462 nsew signal output
rlabel metal2 s 340326 159200 340382 160000 6 eu0_instruction[17]
port 463 nsew signal output
rlabel metal2 s 341338 159200 341394 160000 6 eu0_instruction[18]
port 464 nsew signal output
rlabel metal2 s 342350 159200 342406 160000 6 eu0_instruction[19]
port 465 nsew signal output
rlabel metal2 s 324134 159200 324190 160000 6 eu0_instruction[1]
port 466 nsew signal output
rlabel metal2 s 343362 159200 343418 160000 6 eu0_instruction[20]
port 467 nsew signal output
rlabel metal2 s 344374 159200 344430 160000 6 eu0_instruction[21]
port 468 nsew signal output
rlabel metal2 s 345386 159200 345442 160000 6 eu0_instruction[22]
port 469 nsew signal output
rlabel metal2 s 346398 159200 346454 160000 6 eu0_instruction[23]
port 470 nsew signal output
rlabel metal2 s 347410 159200 347466 160000 6 eu0_instruction[24]
port 471 nsew signal output
rlabel metal2 s 348422 159200 348478 160000 6 eu0_instruction[25]
port 472 nsew signal output
rlabel metal2 s 349434 159200 349490 160000 6 eu0_instruction[26]
port 473 nsew signal output
rlabel metal2 s 350446 159200 350502 160000 6 eu0_instruction[27]
port 474 nsew signal output
rlabel metal2 s 351458 159200 351514 160000 6 eu0_instruction[28]
port 475 nsew signal output
rlabel metal2 s 352470 159200 352526 160000 6 eu0_instruction[29]
port 476 nsew signal output
rlabel metal2 s 325146 159200 325202 160000 6 eu0_instruction[2]
port 477 nsew signal output
rlabel metal2 s 353482 159200 353538 160000 6 eu0_instruction[30]
port 478 nsew signal output
rlabel metal2 s 354494 159200 354550 160000 6 eu0_instruction[31]
port 479 nsew signal output
rlabel metal2 s 355506 159200 355562 160000 6 eu0_instruction[32]
port 480 nsew signal output
rlabel metal2 s 356518 159200 356574 160000 6 eu0_instruction[33]
port 481 nsew signal output
rlabel metal2 s 357530 159200 357586 160000 6 eu0_instruction[34]
port 482 nsew signal output
rlabel metal2 s 358542 159200 358598 160000 6 eu0_instruction[35]
port 483 nsew signal output
rlabel metal2 s 359554 159200 359610 160000 6 eu0_instruction[36]
port 484 nsew signal output
rlabel metal2 s 360566 159200 360622 160000 6 eu0_instruction[37]
port 485 nsew signal output
rlabel metal2 s 361578 159200 361634 160000 6 eu0_instruction[38]
port 486 nsew signal output
rlabel metal2 s 362590 159200 362646 160000 6 eu0_instruction[39]
port 487 nsew signal output
rlabel metal2 s 326158 159200 326214 160000 6 eu0_instruction[3]
port 488 nsew signal output
rlabel metal2 s 363602 159200 363658 160000 6 eu0_instruction[40]
port 489 nsew signal output
rlabel metal2 s 364614 159200 364670 160000 6 eu0_instruction[41]
port 490 nsew signal output
rlabel metal2 s 327170 159200 327226 160000 6 eu0_instruction[4]
port 491 nsew signal output
rlabel metal2 s 328182 159200 328238 160000 6 eu0_instruction[5]
port 492 nsew signal output
rlabel metal2 s 329194 159200 329250 160000 6 eu0_instruction[6]
port 493 nsew signal output
rlabel metal2 s 330206 159200 330262 160000 6 eu0_instruction[7]
port 494 nsew signal output
rlabel metal2 s 331218 159200 331274 160000 6 eu0_instruction[8]
port 495 nsew signal output
rlabel metal2 s 332230 159200 332286 160000 6 eu0_instruction[9]
port 496 nsew signal output
rlabel metal3 s 439200 85416 440000 85536 6 eu1_busy
port 497 nsew signal input
rlabel metal3 s 439200 85960 440000 86080 6 eu1_instruction[0]
port 498 nsew signal output
rlabel metal3 s 439200 91400 440000 91520 6 eu1_instruction[10]
port 499 nsew signal output
rlabel metal3 s 439200 91944 440000 92064 6 eu1_instruction[11]
port 500 nsew signal output
rlabel metal3 s 439200 92488 440000 92608 6 eu1_instruction[12]
port 501 nsew signal output
rlabel metal3 s 439200 93032 440000 93152 6 eu1_instruction[13]
port 502 nsew signal output
rlabel metal3 s 439200 93576 440000 93696 6 eu1_instruction[14]
port 503 nsew signal output
rlabel metal3 s 439200 94120 440000 94240 6 eu1_instruction[15]
port 504 nsew signal output
rlabel metal3 s 439200 94664 440000 94784 6 eu1_instruction[16]
port 505 nsew signal output
rlabel metal3 s 439200 95208 440000 95328 6 eu1_instruction[17]
port 506 nsew signal output
rlabel metal3 s 439200 95752 440000 95872 6 eu1_instruction[18]
port 507 nsew signal output
rlabel metal3 s 439200 96296 440000 96416 6 eu1_instruction[19]
port 508 nsew signal output
rlabel metal3 s 439200 86504 440000 86624 6 eu1_instruction[1]
port 509 nsew signal output
rlabel metal3 s 439200 96840 440000 96960 6 eu1_instruction[20]
port 510 nsew signal output
rlabel metal3 s 439200 97384 440000 97504 6 eu1_instruction[21]
port 511 nsew signal output
rlabel metal3 s 439200 97928 440000 98048 6 eu1_instruction[22]
port 512 nsew signal output
rlabel metal3 s 439200 98472 440000 98592 6 eu1_instruction[23]
port 513 nsew signal output
rlabel metal3 s 439200 99016 440000 99136 6 eu1_instruction[24]
port 514 nsew signal output
rlabel metal3 s 439200 99560 440000 99680 6 eu1_instruction[25]
port 515 nsew signal output
rlabel metal3 s 439200 100104 440000 100224 6 eu1_instruction[26]
port 516 nsew signal output
rlabel metal3 s 439200 100648 440000 100768 6 eu1_instruction[27]
port 517 nsew signal output
rlabel metal3 s 439200 101192 440000 101312 6 eu1_instruction[28]
port 518 nsew signal output
rlabel metal3 s 439200 101736 440000 101856 6 eu1_instruction[29]
port 519 nsew signal output
rlabel metal3 s 439200 87048 440000 87168 6 eu1_instruction[2]
port 520 nsew signal output
rlabel metal3 s 439200 102280 440000 102400 6 eu1_instruction[30]
port 521 nsew signal output
rlabel metal3 s 439200 102824 440000 102944 6 eu1_instruction[31]
port 522 nsew signal output
rlabel metal3 s 439200 103368 440000 103488 6 eu1_instruction[32]
port 523 nsew signal output
rlabel metal3 s 439200 103912 440000 104032 6 eu1_instruction[33]
port 524 nsew signal output
rlabel metal3 s 439200 104456 440000 104576 6 eu1_instruction[34]
port 525 nsew signal output
rlabel metal3 s 439200 105000 440000 105120 6 eu1_instruction[35]
port 526 nsew signal output
rlabel metal3 s 439200 105544 440000 105664 6 eu1_instruction[36]
port 527 nsew signal output
rlabel metal3 s 439200 106088 440000 106208 6 eu1_instruction[37]
port 528 nsew signal output
rlabel metal3 s 439200 106632 440000 106752 6 eu1_instruction[38]
port 529 nsew signal output
rlabel metal3 s 439200 107176 440000 107296 6 eu1_instruction[39]
port 530 nsew signal output
rlabel metal3 s 439200 87592 440000 87712 6 eu1_instruction[3]
port 531 nsew signal output
rlabel metal3 s 439200 107720 440000 107840 6 eu1_instruction[40]
port 532 nsew signal output
rlabel metal3 s 439200 108264 440000 108384 6 eu1_instruction[41]
port 533 nsew signal output
rlabel metal3 s 439200 88136 440000 88256 6 eu1_instruction[4]
port 534 nsew signal output
rlabel metal3 s 439200 88680 440000 88800 6 eu1_instruction[5]
port 535 nsew signal output
rlabel metal3 s 439200 89224 440000 89344 6 eu1_instruction[6]
port 536 nsew signal output
rlabel metal3 s 439200 89768 440000 89888 6 eu1_instruction[7]
port 537 nsew signal output
rlabel metal3 s 439200 90312 440000 90432 6 eu1_instruction[8]
port 538 nsew signal output
rlabel metal3 s 439200 90856 440000 90976 6 eu1_instruction[9]
port 539 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 eu2_busy
port 540 nsew signal input
rlabel metal3 s 0 84872 800 84992 6 eu2_instruction[0]
port 541 nsew signal output
rlabel metal3 s 0 90312 800 90432 6 eu2_instruction[10]
port 542 nsew signal output
rlabel metal3 s 0 90856 800 90976 6 eu2_instruction[11]
port 543 nsew signal output
rlabel metal3 s 0 91400 800 91520 6 eu2_instruction[12]
port 544 nsew signal output
rlabel metal3 s 0 91944 800 92064 6 eu2_instruction[13]
port 545 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 eu2_instruction[14]
port 546 nsew signal output
rlabel metal3 s 0 93032 800 93152 6 eu2_instruction[15]
port 547 nsew signal output
rlabel metal3 s 0 93576 800 93696 6 eu2_instruction[16]
port 548 nsew signal output
rlabel metal3 s 0 94120 800 94240 6 eu2_instruction[17]
port 549 nsew signal output
rlabel metal3 s 0 94664 800 94784 6 eu2_instruction[18]
port 550 nsew signal output
rlabel metal3 s 0 95208 800 95328 6 eu2_instruction[19]
port 551 nsew signal output
rlabel metal3 s 0 85416 800 85536 6 eu2_instruction[1]
port 552 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 eu2_instruction[20]
port 553 nsew signal output
rlabel metal3 s 0 96296 800 96416 6 eu2_instruction[21]
port 554 nsew signal output
rlabel metal3 s 0 96840 800 96960 6 eu2_instruction[22]
port 555 nsew signal output
rlabel metal3 s 0 97384 800 97504 6 eu2_instruction[23]
port 556 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 eu2_instruction[24]
port 557 nsew signal output
rlabel metal3 s 0 98472 800 98592 6 eu2_instruction[25]
port 558 nsew signal output
rlabel metal3 s 0 99016 800 99136 6 eu2_instruction[26]
port 559 nsew signal output
rlabel metal3 s 0 99560 800 99680 6 eu2_instruction[27]
port 560 nsew signal output
rlabel metal3 s 0 100104 800 100224 6 eu2_instruction[28]
port 561 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 eu2_instruction[29]
port 562 nsew signal output
rlabel metal3 s 0 85960 800 86080 6 eu2_instruction[2]
port 563 nsew signal output
rlabel metal3 s 0 101192 800 101312 6 eu2_instruction[30]
port 564 nsew signal output
rlabel metal3 s 0 101736 800 101856 6 eu2_instruction[31]
port 565 nsew signal output
rlabel metal3 s 0 102280 800 102400 6 eu2_instruction[32]
port 566 nsew signal output
rlabel metal3 s 0 102824 800 102944 6 eu2_instruction[33]
port 567 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 eu2_instruction[34]
port 568 nsew signal output
rlabel metal3 s 0 103912 800 104032 6 eu2_instruction[35]
port 569 nsew signal output
rlabel metal3 s 0 104456 800 104576 6 eu2_instruction[36]
port 570 nsew signal output
rlabel metal3 s 0 105000 800 105120 6 eu2_instruction[37]
port 571 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 eu2_instruction[38]
port 572 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 eu2_instruction[39]
port 573 nsew signal output
rlabel metal3 s 0 86504 800 86624 6 eu2_instruction[3]
port 574 nsew signal output
rlabel metal3 s 0 106632 800 106752 6 eu2_instruction[40]
port 575 nsew signal output
rlabel metal3 s 0 107176 800 107296 6 eu2_instruction[41]
port 576 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 eu2_instruction[4]
port 577 nsew signal output
rlabel metal3 s 0 87592 800 87712 6 eu2_instruction[5]
port 578 nsew signal output
rlabel metal3 s 0 88136 800 88256 6 eu2_instruction[6]
port 579 nsew signal output
rlabel metal3 s 0 88680 800 88800 6 eu2_instruction[7]
port 580 nsew signal output
rlabel metal3 s 0 89224 800 89344 6 eu2_instruction[8]
port 581 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 eu2_instruction[9]
port 582 nsew signal output
rlabel metal2 s 431406 159200 431462 160000 6 int_return0
port 583 nsew signal input
rlabel metal3 s 439200 144168 440000 144288 6 int_return1
port 584 nsew signal input
rlabel metal3 s 0 143080 800 143200 6 int_return2
port 585 nsew signal input
rlabel metal2 s 232134 0 232190 800 6 io_in[0]
port 586 nsew signal input
rlabel metal2 s 249614 0 249670 800 6 io_in[10]
port 587 nsew signal input
rlabel metal2 s 251362 0 251418 800 6 io_in[11]
port 588 nsew signal input
rlabel metal2 s 253110 0 253166 800 6 io_in[12]
port 589 nsew signal input
rlabel metal2 s 254858 0 254914 800 6 io_in[13]
port 590 nsew signal input
rlabel metal2 s 256606 0 256662 800 6 io_in[14]
port 591 nsew signal input
rlabel metal2 s 258354 0 258410 800 6 io_in[15]
port 592 nsew signal input
rlabel metal2 s 260102 0 260158 800 6 io_in[16]
port 593 nsew signal input
rlabel metal2 s 261850 0 261906 800 6 io_in[17]
port 594 nsew signal input
rlabel metal2 s 263598 0 263654 800 6 io_in[18]
port 595 nsew signal input
rlabel metal2 s 265346 0 265402 800 6 io_in[19]
port 596 nsew signal input
rlabel metal2 s 233882 0 233938 800 6 io_in[1]
port 597 nsew signal input
rlabel metal2 s 267094 0 267150 800 6 io_in[20]
port 598 nsew signal input
rlabel metal2 s 268842 0 268898 800 6 io_in[21]
port 599 nsew signal input
rlabel metal2 s 270590 0 270646 800 6 io_in[22]
port 600 nsew signal input
rlabel metal2 s 272338 0 272394 800 6 io_in[23]
port 601 nsew signal input
rlabel metal2 s 274086 0 274142 800 6 io_in[24]
port 602 nsew signal input
rlabel metal2 s 275834 0 275890 800 6 io_in[25]
port 603 nsew signal input
rlabel metal2 s 277582 0 277638 800 6 io_in[26]
port 604 nsew signal input
rlabel metal2 s 279330 0 279386 800 6 io_in[27]
port 605 nsew signal input
rlabel metal2 s 281078 0 281134 800 6 io_in[28]
port 606 nsew signal input
rlabel metal2 s 282826 0 282882 800 6 io_in[29]
port 607 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 io_in[2]
port 608 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 io_in[30]
port 609 nsew signal input
rlabel metal2 s 286322 0 286378 800 6 io_in[31]
port 610 nsew signal input
rlabel metal2 s 288070 0 288126 800 6 io_in[32]
port 611 nsew signal input
rlabel metal2 s 289818 0 289874 800 6 io_in[33]
port 612 nsew signal input
rlabel metal2 s 291566 0 291622 800 6 io_in[34]
port 613 nsew signal input
rlabel metal2 s 293314 0 293370 800 6 io_in[35]
port 614 nsew signal input
rlabel metal2 s 237378 0 237434 800 6 io_in[3]
port 615 nsew signal input
rlabel metal2 s 239126 0 239182 800 6 io_in[4]
port 616 nsew signal input
rlabel metal2 s 240874 0 240930 800 6 io_in[5]
port 617 nsew signal input
rlabel metal2 s 242622 0 242678 800 6 io_in[6]
port 618 nsew signal input
rlabel metal2 s 244370 0 244426 800 6 io_in[7]
port 619 nsew signal input
rlabel metal2 s 246118 0 246174 800 6 io_in[8]
port 620 nsew signal input
rlabel metal2 s 247866 0 247922 800 6 io_in[9]
port 621 nsew signal input
rlabel metal2 s 295062 0 295118 800 6 io_oeb[0]
port 622 nsew signal output
rlabel metal2 s 312542 0 312598 800 6 io_oeb[10]
port 623 nsew signal output
rlabel metal2 s 314290 0 314346 800 6 io_oeb[11]
port 624 nsew signal output
rlabel metal2 s 316038 0 316094 800 6 io_oeb[12]
port 625 nsew signal output
rlabel metal2 s 317786 0 317842 800 6 io_oeb[13]
port 626 nsew signal output
rlabel metal2 s 319534 0 319590 800 6 io_oeb[14]
port 627 nsew signal output
rlabel metal2 s 321282 0 321338 800 6 io_oeb[15]
port 628 nsew signal output
rlabel metal2 s 323030 0 323086 800 6 io_oeb[16]
port 629 nsew signal output
rlabel metal2 s 324778 0 324834 800 6 io_oeb[17]
port 630 nsew signal output
rlabel metal2 s 326526 0 326582 800 6 io_oeb[18]
port 631 nsew signal output
rlabel metal2 s 328274 0 328330 800 6 io_oeb[19]
port 632 nsew signal output
rlabel metal2 s 296810 0 296866 800 6 io_oeb[1]
port 633 nsew signal output
rlabel metal2 s 330022 0 330078 800 6 io_oeb[20]
port 634 nsew signal output
rlabel metal2 s 331770 0 331826 800 6 io_oeb[21]
port 635 nsew signal output
rlabel metal2 s 333518 0 333574 800 6 io_oeb[22]
port 636 nsew signal output
rlabel metal2 s 335266 0 335322 800 6 io_oeb[23]
port 637 nsew signal output
rlabel metal2 s 337014 0 337070 800 6 io_oeb[24]
port 638 nsew signal output
rlabel metal2 s 338762 0 338818 800 6 io_oeb[25]
port 639 nsew signal output
rlabel metal2 s 340510 0 340566 800 6 io_oeb[26]
port 640 nsew signal output
rlabel metal2 s 342258 0 342314 800 6 io_oeb[27]
port 641 nsew signal output
rlabel metal2 s 344006 0 344062 800 6 io_oeb[28]
port 642 nsew signal output
rlabel metal2 s 345754 0 345810 800 6 io_oeb[29]
port 643 nsew signal output
rlabel metal2 s 298558 0 298614 800 6 io_oeb[2]
port 644 nsew signal output
rlabel metal2 s 347502 0 347558 800 6 io_oeb[30]
port 645 nsew signal output
rlabel metal2 s 349250 0 349306 800 6 io_oeb[31]
port 646 nsew signal output
rlabel metal2 s 350998 0 351054 800 6 io_oeb[32]
port 647 nsew signal output
rlabel metal2 s 352746 0 352802 800 6 io_oeb[33]
port 648 nsew signal output
rlabel metal2 s 354494 0 354550 800 6 io_oeb[34]
port 649 nsew signal output
rlabel metal2 s 356242 0 356298 800 6 io_oeb[35]
port 650 nsew signal output
rlabel metal2 s 300306 0 300362 800 6 io_oeb[3]
port 651 nsew signal output
rlabel metal2 s 302054 0 302110 800 6 io_oeb[4]
port 652 nsew signal output
rlabel metal2 s 303802 0 303858 800 6 io_oeb[5]
port 653 nsew signal output
rlabel metal2 s 305550 0 305606 800 6 io_oeb[6]
port 654 nsew signal output
rlabel metal2 s 307298 0 307354 800 6 io_oeb[7]
port 655 nsew signal output
rlabel metal2 s 309046 0 309102 800 6 io_oeb[8]
port 656 nsew signal output
rlabel metal2 s 310794 0 310850 800 6 io_oeb[9]
port 657 nsew signal output
rlabel metal2 s 357990 0 358046 800 6 io_out[0]
port 658 nsew signal output
rlabel metal2 s 375470 0 375526 800 6 io_out[10]
port 659 nsew signal output
rlabel metal2 s 377218 0 377274 800 6 io_out[11]
port 660 nsew signal output
rlabel metal2 s 378966 0 379022 800 6 io_out[12]
port 661 nsew signal output
rlabel metal2 s 380714 0 380770 800 6 io_out[13]
port 662 nsew signal output
rlabel metal2 s 382462 0 382518 800 6 io_out[14]
port 663 nsew signal output
rlabel metal2 s 384210 0 384266 800 6 io_out[15]
port 664 nsew signal output
rlabel metal2 s 385958 0 386014 800 6 io_out[16]
port 665 nsew signal output
rlabel metal2 s 387706 0 387762 800 6 io_out[17]
port 666 nsew signal output
rlabel metal2 s 389454 0 389510 800 6 io_out[18]
port 667 nsew signal output
rlabel metal2 s 391202 0 391258 800 6 io_out[19]
port 668 nsew signal output
rlabel metal2 s 359738 0 359794 800 6 io_out[1]
port 669 nsew signal output
rlabel metal2 s 392950 0 393006 800 6 io_out[20]
port 670 nsew signal output
rlabel metal2 s 394698 0 394754 800 6 io_out[21]
port 671 nsew signal output
rlabel metal2 s 396446 0 396502 800 6 io_out[22]
port 672 nsew signal output
rlabel metal2 s 398194 0 398250 800 6 io_out[23]
port 673 nsew signal output
rlabel metal2 s 399942 0 399998 800 6 io_out[24]
port 674 nsew signal output
rlabel metal2 s 401690 0 401746 800 6 io_out[25]
port 675 nsew signal output
rlabel metal2 s 403438 0 403494 800 6 io_out[26]
port 676 nsew signal output
rlabel metal2 s 405186 0 405242 800 6 io_out[27]
port 677 nsew signal output
rlabel metal2 s 406934 0 406990 800 6 io_out[28]
port 678 nsew signal output
rlabel metal2 s 408682 0 408738 800 6 io_out[29]
port 679 nsew signal output
rlabel metal2 s 361486 0 361542 800 6 io_out[2]
port 680 nsew signal output
rlabel metal2 s 410430 0 410486 800 6 io_out[30]
port 681 nsew signal output
rlabel metal2 s 412178 0 412234 800 6 io_out[31]
port 682 nsew signal output
rlabel metal2 s 413926 0 413982 800 6 io_out[32]
port 683 nsew signal output
rlabel metal2 s 415674 0 415730 800 6 io_out[33]
port 684 nsew signal output
rlabel metal2 s 417422 0 417478 800 6 io_out[34]
port 685 nsew signal output
rlabel metal2 s 419170 0 419226 800 6 io_out[35]
port 686 nsew signal output
rlabel metal2 s 363234 0 363290 800 6 io_out[3]
port 687 nsew signal output
rlabel metal2 s 364982 0 365038 800 6 io_out[4]
port 688 nsew signal output
rlabel metal2 s 366730 0 366786 800 6 io_out[5]
port 689 nsew signal output
rlabel metal2 s 368478 0 368534 800 6 io_out[6]
port 690 nsew signal output
rlabel metal2 s 370226 0 370282 800 6 io_out[7]
port 691 nsew signal output
rlabel metal2 s 371974 0 372030 800 6 io_out[8]
port 692 nsew signal output
rlabel metal2 s 373722 0 373778 800 6 io_out[9]
port 693 nsew signal output
rlabel metal2 s 287702 159200 287758 160000 6 is_load0
port 694 nsew signal input
rlabel metal3 s 439200 66920 440000 67040 6 is_load1
port 695 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 is_load2
port 696 nsew signal input
rlabel metal2 s 288714 159200 288770 160000 6 is_store0
port 697 nsew signal input
rlabel metal3 s 439200 67464 440000 67584 6 is_store1
port 698 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 is_store2
port 699 nsew signal input
rlabel metal2 s 255318 159200 255374 160000 6 loadstore_address0[0]
port 700 nsew signal input
rlabel metal2 s 265438 159200 265494 160000 6 loadstore_address0[10]
port 701 nsew signal input
rlabel metal2 s 266450 159200 266506 160000 6 loadstore_address0[11]
port 702 nsew signal input
rlabel metal2 s 267462 159200 267518 160000 6 loadstore_address0[12]
port 703 nsew signal input
rlabel metal2 s 268474 159200 268530 160000 6 loadstore_address0[13]
port 704 nsew signal input
rlabel metal2 s 269486 159200 269542 160000 6 loadstore_address0[14]
port 705 nsew signal input
rlabel metal2 s 270498 159200 270554 160000 6 loadstore_address0[15]
port 706 nsew signal input
rlabel metal2 s 271510 159200 271566 160000 6 loadstore_address0[16]
port 707 nsew signal input
rlabel metal2 s 272522 159200 272578 160000 6 loadstore_address0[17]
port 708 nsew signal input
rlabel metal2 s 273534 159200 273590 160000 6 loadstore_address0[18]
port 709 nsew signal input
rlabel metal2 s 274546 159200 274602 160000 6 loadstore_address0[19]
port 710 nsew signal input
rlabel metal2 s 256330 159200 256386 160000 6 loadstore_address0[1]
port 711 nsew signal input
rlabel metal2 s 275558 159200 275614 160000 6 loadstore_address0[20]
port 712 nsew signal input
rlabel metal2 s 276570 159200 276626 160000 6 loadstore_address0[21]
port 713 nsew signal input
rlabel metal2 s 277582 159200 277638 160000 6 loadstore_address0[22]
port 714 nsew signal input
rlabel metal2 s 278594 159200 278650 160000 6 loadstore_address0[23]
port 715 nsew signal input
rlabel metal2 s 279606 159200 279662 160000 6 loadstore_address0[24]
port 716 nsew signal input
rlabel metal2 s 280618 159200 280674 160000 6 loadstore_address0[25]
port 717 nsew signal input
rlabel metal2 s 281630 159200 281686 160000 6 loadstore_address0[26]
port 718 nsew signal input
rlabel metal2 s 282642 159200 282698 160000 6 loadstore_address0[27]
port 719 nsew signal input
rlabel metal2 s 283654 159200 283710 160000 6 loadstore_address0[28]
port 720 nsew signal input
rlabel metal2 s 284666 159200 284722 160000 6 loadstore_address0[29]
port 721 nsew signal input
rlabel metal2 s 257342 159200 257398 160000 6 loadstore_address0[2]
port 722 nsew signal input
rlabel metal2 s 285678 159200 285734 160000 6 loadstore_address0[30]
port 723 nsew signal input
rlabel metal2 s 286690 159200 286746 160000 6 loadstore_address0[31]
port 724 nsew signal input
rlabel metal2 s 258354 159200 258410 160000 6 loadstore_address0[3]
port 725 nsew signal input
rlabel metal2 s 259366 159200 259422 160000 6 loadstore_address0[4]
port 726 nsew signal input
rlabel metal2 s 260378 159200 260434 160000 6 loadstore_address0[5]
port 727 nsew signal input
rlabel metal2 s 261390 159200 261446 160000 6 loadstore_address0[6]
port 728 nsew signal input
rlabel metal2 s 262402 159200 262458 160000 6 loadstore_address0[7]
port 729 nsew signal input
rlabel metal2 s 263414 159200 263470 160000 6 loadstore_address0[8]
port 730 nsew signal input
rlabel metal2 s 264426 159200 264482 160000 6 loadstore_address0[9]
port 731 nsew signal input
rlabel metal3 s 439200 49512 440000 49632 6 loadstore_address1[0]
port 732 nsew signal input
rlabel metal3 s 439200 54952 440000 55072 6 loadstore_address1[10]
port 733 nsew signal input
rlabel metal3 s 439200 55496 440000 55616 6 loadstore_address1[11]
port 734 nsew signal input
rlabel metal3 s 439200 56040 440000 56160 6 loadstore_address1[12]
port 735 nsew signal input
rlabel metal3 s 439200 56584 440000 56704 6 loadstore_address1[13]
port 736 nsew signal input
rlabel metal3 s 439200 57128 440000 57248 6 loadstore_address1[14]
port 737 nsew signal input
rlabel metal3 s 439200 57672 440000 57792 6 loadstore_address1[15]
port 738 nsew signal input
rlabel metal3 s 439200 58216 440000 58336 6 loadstore_address1[16]
port 739 nsew signal input
rlabel metal3 s 439200 58760 440000 58880 6 loadstore_address1[17]
port 740 nsew signal input
rlabel metal3 s 439200 59304 440000 59424 6 loadstore_address1[18]
port 741 nsew signal input
rlabel metal3 s 439200 59848 440000 59968 6 loadstore_address1[19]
port 742 nsew signal input
rlabel metal3 s 439200 50056 440000 50176 6 loadstore_address1[1]
port 743 nsew signal input
rlabel metal3 s 439200 60392 440000 60512 6 loadstore_address1[20]
port 744 nsew signal input
rlabel metal3 s 439200 60936 440000 61056 6 loadstore_address1[21]
port 745 nsew signal input
rlabel metal3 s 439200 61480 440000 61600 6 loadstore_address1[22]
port 746 nsew signal input
rlabel metal3 s 439200 62024 440000 62144 6 loadstore_address1[23]
port 747 nsew signal input
rlabel metal3 s 439200 62568 440000 62688 6 loadstore_address1[24]
port 748 nsew signal input
rlabel metal3 s 439200 63112 440000 63232 6 loadstore_address1[25]
port 749 nsew signal input
rlabel metal3 s 439200 63656 440000 63776 6 loadstore_address1[26]
port 750 nsew signal input
rlabel metal3 s 439200 64200 440000 64320 6 loadstore_address1[27]
port 751 nsew signal input
rlabel metal3 s 439200 64744 440000 64864 6 loadstore_address1[28]
port 752 nsew signal input
rlabel metal3 s 439200 65288 440000 65408 6 loadstore_address1[29]
port 753 nsew signal input
rlabel metal3 s 439200 50600 440000 50720 6 loadstore_address1[2]
port 754 nsew signal input
rlabel metal3 s 439200 65832 440000 65952 6 loadstore_address1[30]
port 755 nsew signal input
rlabel metal3 s 439200 66376 440000 66496 6 loadstore_address1[31]
port 756 nsew signal input
rlabel metal3 s 439200 51144 440000 51264 6 loadstore_address1[3]
port 757 nsew signal input
rlabel metal3 s 439200 51688 440000 51808 6 loadstore_address1[4]
port 758 nsew signal input
rlabel metal3 s 439200 52232 440000 52352 6 loadstore_address1[5]
port 759 nsew signal input
rlabel metal3 s 439200 52776 440000 52896 6 loadstore_address1[6]
port 760 nsew signal input
rlabel metal3 s 439200 53320 440000 53440 6 loadstore_address1[7]
port 761 nsew signal input
rlabel metal3 s 439200 53864 440000 53984 6 loadstore_address1[8]
port 762 nsew signal input
rlabel metal3 s 439200 54408 440000 54528 6 loadstore_address1[9]
port 763 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 loadstore_address2[0]
port 764 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 loadstore_address2[10]
port 765 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 loadstore_address2[11]
port 766 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 loadstore_address2[12]
port 767 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 loadstore_address2[13]
port 768 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 loadstore_address2[14]
port 769 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 loadstore_address2[15]
port 770 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 loadstore_address2[16]
port 771 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 loadstore_address2[17]
port 772 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 loadstore_address2[18]
port 773 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 loadstore_address2[19]
port 774 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 loadstore_address2[1]
port 775 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 loadstore_address2[20]
port 776 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 loadstore_address2[21]
port 777 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 loadstore_address2[22]
port 778 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 loadstore_address2[23]
port 779 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 loadstore_address2[24]
port 780 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 loadstore_address2[25]
port 781 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 loadstore_address2[26]
port 782 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 loadstore_address2[27]
port 783 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 loadstore_address2[28]
port 784 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 loadstore_address2[29]
port 785 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 loadstore_address2[2]
port 786 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 loadstore_address2[30]
port 787 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 loadstore_address2[31]
port 788 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 loadstore_address2[3]
port 789 nsew signal input
rlabel metal3 s 0 50600 800 50720 6 loadstore_address2[4]
port 790 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 loadstore_address2[5]
port 791 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 loadstore_address2[6]
port 792 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 loadstore_address2[7]
port 793 nsew signal input
rlabel metal3 s 0 52776 800 52896 6 loadstore_address2[8]
port 794 nsew signal input
rlabel metal3 s 0 53320 800 53440 6 loadstore_address2[9]
port 795 nsew signal input
rlabel metal2 s 290738 159200 290794 160000 6 loadstore_size0[0]
port 796 nsew signal input
rlabel metal2 s 291750 159200 291806 160000 6 loadstore_size0[1]
port 797 nsew signal input
rlabel metal3 s 439200 68552 440000 68672 6 loadstore_size1[0]
port 798 nsew signal input
rlabel metal3 s 439200 69096 440000 69216 6 loadstore_size1[1]
port 799 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 loadstore_size2[0]
port 800 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 loadstore_size2[1]
port 801 nsew signal input
rlabel metal2 s 293774 159200 293830 160000 6 new_PC0[0]
port 802 nsew signal input
rlabel metal2 s 303894 159200 303950 160000 6 new_PC0[10]
port 803 nsew signal input
rlabel metal2 s 304906 159200 304962 160000 6 new_PC0[11]
port 804 nsew signal input
rlabel metal2 s 305918 159200 305974 160000 6 new_PC0[12]
port 805 nsew signal input
rlabel metal2 s 306930 159200 306986 160000 6 new_PC0[13]
port 806 nsew signal input
rlabel metal2 s 307942 159200 307998 160000 6 new_PC0[14]
port 807 nsew signal input
rlabel metal2 s 308954 159200 309010 160000 6 new_PC0[15]
port 808 nsew signal input
rlabel metal2 s 309966 159200 310022 160000 6 new_PC0[16]
port 809 nsew signal input
rlabel metal2 s 310978 159200 311034 160000 6 new_PC0[17]
port 810 nsew signal input
rlabel metal2 s 311990 159200 312046 160000 6 new_PC0[18]
port 811 nsew signal input
rlabel metal2 s 313002 159200 313058 160000 6 new_PC0[19]
port 812 nsew signal input
rlabel metal2 s 294786 159200 294842 160000 6 new_PC0[1]
port 813 nsew signal input
rlabel metal2 s 314014 159200 314070 160000 6 new_PC0[20]
port 814 nsew signal input
rlabel metal2 s 315026 159200 315082 160000 6 new_PC0[21]
port 815 nsew signal input
rlabel metal2 s 316038 159200 316094 160000 6 new_PC0[22]
port 816 nsew signal input
rlabel metal2 s 317050 159200 317106 160000 6 new_PC0[23]
port 817 nsew signal input
rlabel metal2 s 318062 159200 318118 160000 6 new_PC0[24]
port 818 nsew signal input
rlabel metal2 s 319074 159200 319130 160000 6 new_PC0[25]
port 819 nsew signal input
rlabel metal2 s 320086 159200 320142 160000 6 new_PC0[26]
port 820 nsew signal input
rlabel metal2 s 321098 159200 321154 160000 6 new_PC0[27]
port 821 nsew signal input
rlabel metal2 s 295798 159200 295854 160000 6 new_PC0[2]
port 822 nsew signal input
rlabel metal2 s 296810 159200 296866 160000 6 new_PC0[3]
port 823 nsew signal input
rlabel metal2 s 297822 159200 297878 160000 6 new_PC0[4]
port 824 nsew signal input
rlabel metal2 s 298834 159200 298890 160000 6 new_PC0[5]
port 825 nsew signal input
rlabel metal2 s 299846 159200 299902 160000 6 new_PC0[6]
port 826 nsew signal input
rlabel metal2 s 300858 159200 300914 160000 6 new_PC0[7]
port 827 nsew signal input
rlabel metal2 s 301870 159200 301926 160000 6 new_PC0[8]
port 828 nsew signal input
rlabel metal2 s 302882 159200 302938 160000 6 new_PC0[9]
port 829 nsew signal input
rlabel metal3 s 439200 70184 440000 70304 6 new_PC1[0]
port 830 nsew signal input
rlabel metal3 s 439200 75624 440000 75744 6 new_PC1[10]
port 831 nsew signal input
rlabel metal3 s 439200 76168 440000 76288 6 new_PC1[11]
port 832 nsew signal input
rlabel metal3 s 439200 76712 440000 76832 6 new_PC1[12]
port 833 nsew signal input
rlabel metal3 s 439200 77256 440000 77376 6 new_PC1[13]
port 834 nsew signal input
rlabel metal3 s 439200 77800 440000 77920 6 new_PC1[14]
port 835 nsew signal input
rlabel metal3 s 439200 78344 440000 78464 6 new_PC1[15]
port 836 nsew signal input
rlabel metal3 s 439200 78888 440000 79008 6 new_PC1[16]
port 837 nsew signal input
rlabel metal3 s 439200 79432 440000 79552 6 new_PC1[17]
port 838 nsew signal input
rlabel metal3 s 439200 79976 440000 80096 6 new_PC1[18]
port 839 nsew signal input
rlabel metal3 s 439200 80520 440000 80640 6 new_PC1[19]
port 840 nsew signal input
rlabel metal3 s 439200 70728 440000 70848 6 new_PC1[1]
port 841 nsew signal input
rlabel metal3 s 439200 81064 440000 81184 6 new_PC1[20]
port 842 nsew signal input
rlabel metal3 s 439200 81608 440000 81728 6 new_PC1[21]
port 843 nsew signal input
rlabel metal3 s 439200 82152 440000 82272 6 new_PC1[22]
port 844 nsew signal input
rlabel metal3 s 439200 82696 440000 82816 6 new_PC1[23]
port 845 nsew signal input
rlabel metal3 s 439200 83240 440000 83360 6 new_PC1[24]
port 846 nsew signal input
rlabel metal3 s 439200 83784 440000 83904 6 new_PC1[25]
port 847 nsew signal input
rlabel metal3 s 439200 84328 440000 84448 6 new_PC1[26]
port 848 nsew signal input
rlabel metal3 s 439200 84872 440000 84992 6 new_PC1[27]
port 849 nsew signal input
rlabel metal3 s 439200 71272 440000 71392 6 new_PC1[2]
port 850 nsew signal input
rlabel metal3 s 439200 71816 440000 71936 6 new_PC1[3]
port 851 nsew signal input
rlabel metal3 s 439200 72360 440000 72480 6 new_PC1[4]
port 852 nsew signal input
rlabel metal3 s 439200 72904 440000 73024 6 new_PC1[5]
port 853 nsew signal input
rlabel metal3 s 439200 73448 440000 73568 6 new_PC1[6]
port 854 nsew signal input
rlabel metal3 s 439200 73992 440000 74112 6 new_PC1[7]
port 855 nsew signal input
rlabel metal3 s 439200 74536 440000 74656 6 new_PC1[8]
port 856 nsew signal input
rlabel metal3 s 439200 75080 440000 75200 6 new_PC1[9]
port 857 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 new_PC2[0]
port 858 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 new_PC2[10]
port 859 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 new_PC2[11]
port 860 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 new_PC2[12]
port 861 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 new_PC2[13]
port 862 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 new_PC2[14]
port 863 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 new_PC2[15]
port 864 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 new_PC2[16]
port 865 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 new_PC2[17]
port 866 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 new_PC2[18]
port 867 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 new_PC2[19]
port 868 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 new_PC2[1]
port 869 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 new_PC2[20]
port 870 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 new_PC2[21]
port 871 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 new_PC2[22]
port 872 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 new_PC2[23]
port 873 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 new_PC2[24]
port 874 nsew signal input
rlabel metal3 s 0 82696 800 82816 6 new_PC2[25]
port 875 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 new_PC2[26]
port 876 nsew signal input
rlabel metal3 s 0 83784 800 83904 6 new_PC2[27]
port 877 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 new_PC2[2]
port 878 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 new_PC2[3]
port 879 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 new_PC2[4]
port 880 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 new_PC2[5]
port 881 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 new_PC2[6]
port 882 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 new_PC2[7]
port 883 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 new_PC2[8]
port 884 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 new_PC2[9]
port 885 nsew signal input
rlabel metal2 s 248234 159200 248290 160000 6 pred_idx0[0]
port 886 nsew signal input
rlabel metal2 s 249246 159200 249302 160000 6 pred_idx0[1]
port 887 nsew signal input
rlabel metal2 s 250258 159200 250314 160000 6 pred_idx0[2]
port 888 nsew signal input
rlabel metal3 s 439200 45704 440000 45824 6 pred_idx1[0]
port 889 nsew signal input
rlabel metal3 s 439200 46248 440000 46368 6 pred_idx1[1]
port 890 nsew signal input
rlabel metal3 s 439200 46792 440000 46912 6 pred_idx1[2]
port 891 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 pred_idx2[0]
port 892 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 pred_idx2[1]
port 893 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 pred_idx2[2]
port 894 nsew signal input
rlabel metal2 s 430394 159200 430450 160000 6 pred_val0
port 895 nsew signal output
rlabel metal3 s 439200 143624 440000 143744 6 pred_val1
port 896 nsew signal output
rlabel metal3 s 0 142536 800 142656 6 pred_val2
port 897 nsew signal output
rlabel metal2 s 195610 159200 195666 160000 6 reg1_idx0[0]
port 898 nsew signal input
rlabel metal2 s 196622 159200 196678 160000 6 reg1_idx0[1]
port 899 nsew signal input
rlabel metal2 s 197634 159200 197690 160000 6 reg1_idx0[2]
port 900 nsew signal input
rlabel metal2 s 198646 159200 198702 160000 6 reg1_idx0[3]
port 901 nsew signal input
rlabel metal2 s 199658 159200 199714 160000 6 reg1_idx0[4]
port 902 nsew signal input
rlabel metal2 s 200670 159200 200726 160000 6 reg1_idx0[5]
port 903 nsew signal input
rlabel metal3 s 439200 17416 440000 17536 6 reg1_idx1[0]
port 904 nsew signal input
rlabel metal3 s 439200 17960 440000 18080 6 reg1_idx1[1]
port 905 nsew signal input
rlabel metal3 s 439200 18504 440000 18624 6 reg1_idx1[2]
port 906 nsew signal input
rlabel metal3 s 439200 19048 440000 19168 6 reg1_idx1[3]
port 907 nsew signal input
rlabel metal3 s 439200 19592 440000 19712 6 reg1_idx1[4]
port 908 nsew signal input
rlabel metal3 s 439200 20136 440000 20256 6 reg1_idx1[5]
port 909 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 reg1_idx2[0]
port 910 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 reg1_idx2[1]
port 911 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 reg1_idx2[2]
port 912 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 reg1_idx2[3]
port 913 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 reg1_idx2[4]
port 914 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 reg1_idx2[5]
port 915 nsew signal input
rlabel metal2 s 365626 159200 365682 160000 6 reg1_val0[0]
port 916 nsew signal output
rlabel metal2 s 375746 159200 375802 160000 6 reg1_val0[10]
port 917 nsew signal output
rlabel metal2 s 376758 159200 376814 160000 6 reg1_val0[11]
port 918 nsew signal output
rlabel metal2 s 377770 159200 377826 160000 6 reg1_val0[12]
port 919 nsew signal output
rlabel metal2 s 378782 159200 378838 160000 6 reg1_val0[13]
port 920 nsew signal output
rlabel metal2 s 379794 159200 379850 160000 6 reg1_val0[14]
port 921 nsew signal output
rlabel metal2 s 380806 159200 380862 160000 6 reg1_val0[15]
port 922 nsew signal output
rlabel metal2 s 381818 159200 381874 160000 6 reg1_val0[16]
port 923 nsew signal output
rlabel metal2 s 382830 159200 382886 160000 6 reg1_val0[17]
port 924 nsew signal output
rlabel metal2 s 383842 159200 383898 160000 6 reg1_val0[18]
port 925 nsew signal output
rlabel metal2 s 384854 159200 384910 160000 6 reg1_val0[19]
port 926 nsew signal output
rlabel metal2 s 366638 159200 366694 160000 6 reg1_val0[1]
port 927 nsew signal output
rlabel metal2 s 385866 159200 385922 160000 6 reg1_val0[20]
port 928 nsew signal output
rlabel metal2 s 386878 159200 386934 160000 6 reg1_val0[21]
port 929 nsew signal output
rlabel metal2 s 387890 159200 387946 160000 6 reg1_val0[22]
port 930 nsew signal output
rlabel metal2 s 388902 159200 388958 160000 6 reg1_val0[23]
port 931 nsew signal output
rlabel metal2 s 389914 159200 389970 160000 6 reg1_val0[24]
port 932 nsew signal output
rlabel metal2 s 390926 159200 390982 160000 6 reg1_val0[25]
port 933 nsew signal output
rlabel metal2 s 391938 159200 391994 160000 6 reg1_val0[26]
port 934 nsew signal output
rlabel metal2 s 392950 159200 393006 160000 6 reg1_val0[27]
port 935 nsew signal output
rlabel metal2 s 393962 159200 394018 160000 6 reg1_val0[28]
port 936 nsew signal output
rlabel metal2 s 394974 159200 395030 160000 6 reg1_val0[29]
port 937 nsew signal output
rlabel metal2 s 367650 159200 367706 160000 6 reg1_val0[2]
port 938 nsew signal output
rlabel metal2 s 395986 159200 396042 160000 6 reg1_val0[30]
port 939 nsew signal output
rlabel metal2 s 396998 159200 397054 160000 6 reg1_val0[31]
port 940 nsew signal output
rlabel metal2 s 368662 159200 368718 160000 6 reg1_val0[3]
port 941 nsew signal output
rlabel metal2 s 369674 159200 369730 160000 6 reg1_val0[4]
port 942 nsew signal output
rlabel metal2 s 370686 159200 370742 160000 6 reg1_val0[5]
port 943 nsew signal output
rlabel metal2 s 371698 159200 371754 160000 6 reg1_val0[6]
port 944 nsew signal output
rlabel metal2 s 372710 159200 372766 160000 6 reg1_val0[7]
port 945 nsew signal output
rlabel metal2 s 373722 159200 373778 160000 6 reg1_val0[8]
port 946 nsew signal output
rlabel metal2 s 374734 159200 374790 160000 6 reg1_val0[9]
port 947 nsew signal output
rlabel metal3 s 439200 108808 440000 108928 6 reg1_val1[0]
port 948 nsew signal output
rlabel metal3 s 439200 114248 440000 114368 6 reg1_val1[10]
port 949 nsew signal output
rlabel metal3 s 439200 114792 440000 114912 6 reg1_val1[11]
port 950 nsew signal output
rlabel metal3 s 439200 115336 440000 115456 6 reg1_val1[12]
port 951 nsew signal output
rlabel metal3 s 439200 115880 440000 116000 6 reg1_val1[13]
port 952 nsew signal output
rlabel metal3 s 439200 116424 440000 116544 6 reg1_val1[14]
port 953 nsew signal output
rlabel metal3 s 439200 116968 440000 117088 6 reg1_val1[15]
port 954 nsew signal output
rlabel metal3 s 439200 117512 440000 117632 6 reg1_val1[16]
port 955 nsew signal output
rlabel metal3 s 439200 118056 440000 118176 6 reg1_val1[17]
port 956 nsew signal output
rlabel metal3 s 439200 118600 440000 118720 6 reg1_val1[18]
port 957 nsew signal output
rlabel metal3 s 439200 119144 440000 119264 6 reg1_val1[19]
port 958 nsew signal output
rlabel metal3 s 439200 109352 440000 109472 6 reg1_val1[1]
port 959 nsew signal output
rlabel metal3 s 439200 119688 440000 119808 6 reg1_val1[20]
port 960 nsew signal output
rlabel metal3 s 439200 120232 440000 120352 6 reg1_val1[21]
port 961 nsew signal output
rlabel metal3 s 439200 120776 440000 120896 6 reg1_val1[22]
port 962 nsew signal output
rlabel metal3 s 439200 121320 440000 121440 6 reg1_val1[23]
port 963 nsew signal output
rlabel metal3 s 439200 121864 440000 121984 6 reg1_val1[24]
port 964 nsew signal output
rlabel metal3 s 439200 122408 440000 122528 6 reg1_val1[25]
port 965 nsew signal output
rlabel metal3 s 439200 122952 440000 123072 6 reg1_val1[26]
port 966 nsew signal output
rlabel metal3 s 439200 123496 440000 123616 6 reg1_val1[27]
port 967 nsew signal output
rlabel metal3 s 439200 124040 440000 124160 6 reg1_val1[28]
port 968 nsew signal output
rlabel metal3 s 439200 124584 440000 124704 6 reg1_val1[29]
port 969 nsew signal output
rlabel metal3 s 439200 109896 440000 110016 6 reg1_val1[2]
port 970 nsew signal output
rlabel metal3 s 439200 125128 440000 125248 6 reg1_val1[30]
port 971 nsew signal output
rlabel metal3 s 439200 125672 440000 125792 6 reg1_val1[31]
port 972 nsew signal output
rlabel metal3 s 439200 110440 440000 110560 6 reg1_val1[3]
port 973 nsew signal output
rlabel metal3 s 439200 110984 440000 111104 6 reg1_val1[4]
port 974 nsew signal output
rlabel metal3 s 439200 111528 440000 111648 6 reg1_val1[5]
port 975 nsew signal output
rlabel metal3 s 439200 112072 440000 112192 6 reg1_val1[6]
port 976 nsew signal output
rlabel metal3 s 439200 112616 440000 112736 6 reg1_val1[7]
port 977 nsew signal output
rlabel metal3 s 439200 113160 440000 113280 6 reg1_val1[8]
port 978 nsew signal output
rlabel metal3 s 439200 113704 440000 113824 6 reg1_val1[9]
port 979 nsew signal output
rlabel metal3 s 0 107720 800 107840 6 reg1_val2[0]
port 980 nsew signal output
rlabel metal3 s 0 113160 800 113280 6 reg1_val2[10]
port 981 nsew signal output
rlabel metal3 s 0 113704 800 113824 6 reg1_val2[11]
port 982 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 reg1_val2[12]
port 983 nsew signal output
rlabel metal3 s 0 114792 800 114912 6 reg1_val2[13]
port 984 nsew signal output
rlabel metal3 s 0 115336 800 115456 6 reg1_val2[14]
port 985 nsew signal output
rlabel metal3 s 0 115880 800 116000 6 reg1_val2[15]
port 986 nsew signal output
rlabel metal3 s 0 116424 800 116544 6 reg1_val2[16]
port 987 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 reg1_val2[17]
port 988 nsew signal output
rlabel metal3 s 0 117512 800 117632 6 reg1_val2[18]
port 989 nsew signal output
rlabel metal3 s 0 118056 800 118176 6 reg1_val2[19]
port 990 nsew signal output
rlabel metal3 s 0 108264 800 108384 6 reg1_val2[1]
port 991 nsew signal output
rlabel metal3 s 0 118600 800 118720 6 reg1_val2[20]
port 992 nsew signal output
rlabel metal3 s 0 119144 800 119264 6 reg1_val2[21]
port 993 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 reg1_val2[22]
port 994 nsew signal output
rlabel metal3 s 0 120232 800 120352 6 reg1_val2[23]
port 995 nsew signal output
rlabel metal3 s 0 120776 800 120896 6 reg1_val2[24]
port 996 nsew signal output
rlabel metal3 s 0 121320 800 121440 6 reg1_val2[25]
port 997 nsew signal output
rlabel metal3 s 0 121864 800 121984 6 reg1_val2[26]
port 998 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 reg1_val2[27]
port 999 nsew signal output
rlabel metal3 s 0 122952 800 123072 6 reg1_val2[28]
port 1000 nsew signal output
rlabel metal3 s 0 123496 800 123616 6 reg1_val2[29]
port 1001 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 reg1_val2[2]
port 1002 nsew signal output
rlabel metal3 s 0 124040 800 124160 6 reg1_val2[30]
port 1003 nsew signal output
rlabel metal3 s 0 124584 800 124704 6 reg1_val2[31]
port 1004 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 reg1_val2[3]
port 1005 nsew signal output
rlabel metal3 s 0 109896 800 110016 6 reg1_val2[4]
port 1006 nsew signal output
rlabel metal3 s 0 110440 800 110560 6 reg1_val2[5]
port 1007 nsew signal output
rlabel metal3 s 0 110984 800 111104 6 reg1_val2[6]
port 1008 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 reg1_val2[7]
port 1009 nsew signal output
rlabel metal3 s 0 112072 800 112192 6 reg1_val2[8]
port 1010 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 reg1_val2[9]
port 1011 nsew signal output
rlabel metal2 s 201682 159200 201738 160000 6 reg2_idx0[0]
port 1012 nsew signal input
rlabel metal2 s 202694 159200 202750 160000 6 reg2_idx0[1]
port 1013 nsew signal input
rlabel metal2 s 203706 159200 203762 160000 6 reg2_idx0[2]
port 1014 nsew signal input
rlabel metal2 s 204718 159200 204774 160000 6 reg2_idx0[3]
port 1015 nsew signal input
rlabel metal2 s 205730 159200 205786 160000 6 reg2_idx0[4]
port 1016 nsew signal input
rlabel metal2 s 206742 159200 206798 160000 6 reg2_idx0[5]
port 1017 nsew signal input
rlabel metal3 s 439200 20680 440000 20800 6 reg2_idx1[0]
port 1018 nsew signal input
rlabel metal3 s 439200 21224 440000 21344 6 reg2_idx1[1]
port 1019 nsew signal input
rlabel metal3 s 439200 21768 440000 21888 6 reg2_idx1[2]
port 1020 nsew signal input
rlabel metal3 s 439200 22312 440000 22432 6 reg2_idx1[3]
port 1021 nsew signal input
rlabel metal3 s 439200 22856 440000 22976 6 reg2_idx1[4]
port 1022 nsew signal input
rlabel metal3 s 439200 23400 440000 23520 6 reg2_idx1[5]
port 1023 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 reg2_idx2[0]
port 1024 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 reg2_idx2[1]
port 1025 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 reg2_idx2[2]
port 1026 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 reg2_idx2[3]
port 1027 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 reg2_idx2[4]
port 1028 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 reg2_idx2[5]
port 1029 nsew signal input
rlabel metal2 s 398010 159200 398066 160000 6 reg2_val0[0]
port 1030 nsew signal output
rlabel metal2 s 408130 159200 408186 160000 6 reg2_val0[10]
port 1031 nsew signal output
rlabel metal2 s 409142 159200 409198 160000 6 reg2_val0[11]
port 1032 nsew signal output
rlabel metal2 s 410154 159200 410210 160000 6 reg2_val0[12]
port 1033 nsew signal output
rlabel metal2 s 411166 159200 411222 160000 6 reg2_val0[13]
port 1034 nsew signal output
rlabel metal2 s 412178 159200 412234 160000 6 reg2_val0[14]
port 1035 nsew signal output
rlabel metal2 s 413190 159200 413246 160000 6 reg2_val0[15]
port 1036 nsew signal output
rlabel metal2 s 414202 159200 414258 160000 6 reg2_val0[16]
port 1037 nsew signal output
rlabel metal2 s 415214 159200 415270 160000 6 reg2_val0[17]
port 1038 nsew signal output
rlabel metal2 s 416226 159200 416282 160000 6 reg2_val0[18]
port 1039 nsew signal output
rlabel metal2 s 417238 159200 417294 160000 6 reg2_val0[19]
port 1040 nsew signal output
rlabel metal2 s 399022 159200 399078 160000 6 reg2_val0[1]
port 1041 nsew signal output
rlabel metal2 s 418250 159200 418306 160000 6 reg2_val0[20]
port 1042 nsew signal output
rlabel metal2 s 419262 159200 419318 160000 6 reg2_val0[21]
port 1043 nsew signal output
rlabel metal2 s 420274 159200 420330 160000 6 reg2_val0[22]
port 1044 nsew signal output
rlabel metal2 s 421286 159200 421342 160000 6 reg2_val0[23]
port 1045 nsew signal output
rlabel metal2 s 422298 159200 422354 160000 6 reg2_val0[24]
port 1046 nsew signal output
rlabel metal2 s 423310 159200 423366 160000 6 reg2_val0[25]
port 1047 nsew signal output
rlabel metal2 s 424322 159200 424378 160000 6 reg2_val0[26]
port 1048 nsew signal output
rlabel metal2 s 425334 159200 425390 160000 6 reg2_val0[27]
port 1049 nsew signal output
rlabel metal2 s 426346 159200 426402 160000 6 reg2_val0[28]
port 1050 nsew signal output
rlabel metal2 s 427358 159200 427414 160000 6 reg2_val0[29]
port 1051 nsew signal output
rlabel metal2 s 400034 159200 400090 160000 6 reg2_val0[2]
port 1052 nsew signal output
rlabel metal2 s 428370 159200 428426 160000 6 reg2_val0[30]
port 1053 nsew signal output
rlabel metal2 s 429382 159200 429438 160000 6 reg2_val0[31]
port 1054 nsew signal output
rlabel metal2 s 401046 159200 401102 160000 6 reg2_val0[3]
port 1055 nsew signal output
rlabel metal2 s 402058 159200 402114 160000 6 reg2_val0[4]
port 1056 nsew signal output
rlabel metal2 s 403070 159200 403126 160000 6 reg2_val0[5]
port 1057 nsew signal output
rlabel metal2 s 404082 159200 404138 160000 6 reg2_val0[6]
port 1058 nsew signal output
rlabel metal2 s 405094 159200 405150 160000 6 reg2_val0[7]
port 1059 nsew signal output
rlabel metal2 s 406106 159200 406162 160000 6 reg2_val0[8]
port 1060 nsew signal output
rlabel metal2 s 407118 159200 407174 160000 6 reg2_val0[9]
port 1061 nsew signal output
rlabel metal3 s 439200 126216 440000 126336 6 reg2_val1[0]
port 1062 nsew signal output
rlabel metal3 s 439200 131656 440000 131776 6 reg2_val1[10]
port 1063 nsew signal output
rlabel metal3 s 439200 132200 440000 132320 6 reg2_val1[11]
port 1064 nsew signal output
rlabel metal3 s 439200 132744 440000 132864 6 reg2_val1[12]
port 1065 nsew signal output
rlabel metal3 s 439200 133288 440000 133408 6 reg2_val1[13]
port 1066 nsew signal output
rlabel metal3 s 439200 133832 440000 133952 6 reg2_val1[14]
port 1067 nsew signal output
rlabel metal3 s 439200 134376 440000 134496 6 reg2_val1[15]
port 1068 nsew signal output
rlabel metal3 s 439200 134920 440000 135040 6 reg2_val1[16]
port 1069 nsew signal output
rlabel metal3 s 439200 135464 440000 135584 6 reg2_val1[17]
port 1070 nsew signal output
rlabel metal3 s 439200 136008 440000 136128 6 reg2_val1[18]
port 1071 nsew signal output
rlabel metal3 s 439200 136552 440000 136672 6 reg2_val1[19]
port 1072 nsew signal output
rlabel metal3 s 439200 126760 440000 126880 6 reg2_val1[1]
port 1073 nsew signal output
rlabel metal3 s 439200 137096 440000 137216 6 reg2_val1[20]
port 1074 nsew signal output
rlabel metal3 s 439200 137640 440000 137760 6 reg2_val1[21]
port 1075 nsew signal output
rlabel metal3 s 439200 138184 440000 138304 6 reg2_val1[22]
port 1076 nsew signal output
rlabel metal3 s 439200 138728 440000 138848 6 reg2_val1[23]
port 1077 nsew signal output
rlabel metal3 s 439200 139272 440000 139392 6 reg2_val1[24]
port 1078 nsew signal output
rlabel metal3 s 439200 139816 440000 139936 6 reg2_val1[25]
port 1079 nsew signal output
rlabel metal3 s 439200 140360 440000 140480 6 reg2_val1[26]
port 1080 nsew signal output
rlabel metal3 s 439200 140904 440000 141024 6 reg2_val1[27]
port 1081 nsew signal output
rlabel metal3 s 439200 141448 440000 141568 6 reg2_val1[28]
port 1082 nsew signal output
rlabel metal3 s 439200 141992 440000 142112 6 reg2_val1[29]
port 1083 nsew signal output
rlabel metal3 s 439200 127304 440000 127424 6 reg2_val1[2]
port 1084 nsew signal output
rlabel metal3 s 439200 142536 440000 142656 6 reg2_val1[30]
port 1085 nsew signal output
rlabel metal3 s 439200 143080 440000 143200 6 reg2_val1[31]
port 1086 nsew signal output
rlabel metal3 s 439200 127848 440000 127968 6 reg2_val1[3]
port 1087 nsew signal output
rlabel metal3 s 439200 128392 440000 128512 6 reg2_val1[4]
port 1088 nsew signal output
rlabel metal3 s 439200 128936 440000 129056 6 reg2_val1[5]
port 1089 nsew signal output
rlabel metal3 s 439200 129480 440000 129600 6 reg2_val1[6]
port 1090 nsew signal output
rlabel metal3 s 439200 130024 440000 130144 6 reg2_val1[7]
port 1091 nsew signal output
rlabel metal3 s 439200 130568 440000 130688 6 reg2_val1[8]
port 1092 nsew signal output
rlabel metal3 s 439200 131112 440000 131232 6 reg2_val1[9]
port 1093 nsew signal output
rlabel metal3 s 0 125128 800 125248 6 reg2_val2[0]
port 1094 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 reg2_val2[10]
port 1095 nsew signal output
rlabel metal3 s 0 131112 800 131232 6 reg2_val2[11]
port 1096 nsew signal output
rlabel metal3 s 0 131656 800 131776 6 reg2_val2[12]
port 1097 nsew signal output
rlabel metal3 s 0 132200 800 132320 6 reg2_val2[13]
port 1098 nsew signal output
rlabel metal3 s 0 132744 800 132864 6 reg2_val2[14]
port 1099 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 reg2_val2[15]
port 1100 nsew signal output
rlabel metal3 s 0 133832 800 133952 6 reg2_val2[16]
port 1101 nsew signal output
rlabel metal3 s 0 134376 800 134496 6 reg2_val2[17]
port 1102 nsew signal output
rlabel metal3 s 0 134920 800 135040 6 reg2_val2[18]
port 1103 nsew signal output
rlabel metal3 s 0 135464 800 135584 6 reg2_val2[19]
port 1104 nsew signal output
rlabel metal3 s 0 125672 800 125792 6 reg2_val2[1]
port 1105 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 reg2_val2[20]
port 1106 nsew signal output
rlabel metal3 s 0 136552 800 136672 6 reg2_val2[21]
port 1107 nsew signal output
rlabel metal3 s 0 137096 800 137216 6 reg2_val2[22]
port 1108 nsew signal output
rlabel metal3 s 0 137640 800 137760 6 reg2_val2[23]
port 1109 nsew signal output
rlabel metal3 s 0 138184 800 138304 6 reg2_val2[24]
port 1110 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 reg2_val2[25]
port 1111 nsew signal output
rlabel metal3 s 0 139272 800 139392 6 reg2_val2[26]
port 1112 nsew signal output
rlabel metal3 s 0 139816 800 139936 6 reg2_val2[27]
port 1113 nsew signal output
rlabel metal3 s 0 140360 800 140480 6 reg2_val2[28]
port 1114 nsew signal output
rlabel metal3 s 0 140904 800 141024 6 reg2_val2[29]
port 1115 nsew signal output
rlabel metal3 s 0 126216 800 126336 6 reg2_val2[2]
port 1116 nsew signal output
rlabel metal3 s 0 141448 800 141568 6 reg2_val2[30]
port 1117 nsew signal output
rlabel metal3 s 0 141992 800 142112 6 reg2_val2[31]
port 1118 nsew signal output
rlabel metal3 s 0 126760 800 126880 6 reg2_val2[3]
port 1119 nsew signal output
rlabel metal3 s 0 127304 800 127424 6 reg2_val2[4]
port 1120 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 reg2_val2[5]
port 1121 nsew signal output
rlabel metal3 s 0 128392 800 128512 6 reg2_val2[6]
port 1122 nsew signal output
rlabel metal3 s 0 128936 800 129056 6 reg2_val2[7]
port 1123 nsew signal output
rlabel metal3 s 0 129480 800 129600 6 reg2_val2[8]
port 1124 nsew signal output
rlabel metal3 s 0 130024 800 130144 6 reg2_val2[9]
port 1125 nsew signal output
rlabel metal2 s 166262 159200 166318 160000 6 rst_eu
port 1126 nsew signal output
rlabel metal2 s 422666 0 422722 800 6 rst_n
port 1127 nsew signal input
rlabel metal2 s 289726 159200 289782 160000 6 sign_extend0
port 1128 nsew signal input
rlabel metal3 s 439200 68008 440000 68128 6 sign_extend1
port 1129 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 sign_extend2
port 1130 nsew signal input
rlabel metal2 s 292762 159200 292818 160000 6 take_branch0
port 1131 nsew signal input
rlabel metal3 s 439200 69640 440000 69760 6 take_branch1
port 1132 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 take_branch2
port 1133 nsew signal input
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 157808 6 vccd1
port 1134 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 157808 6 vssd1
port 1135 nsew ground bidirectional
rlabel metal2 s 420918 0 420974 800 6 wb_clk_i
port 1136 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 440000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 162843634
string GDS_FILE /home/lucah/Desktop/ci2406-rej-pommedeterrible-tholin/openlane/VLIW/runs/24_06_06_12_50/results/signoff/vliw.magic.gds
string GDS_START 1470480
<< end >>

