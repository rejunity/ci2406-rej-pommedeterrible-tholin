* NGSPICE file created from execution_unit.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_2 abstract view
.subckt sky130_fd_sc_hd__a41oi_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

.subckt execution_unit busy curr_PC[0] curr_PC[10] curr_PC[11] curr_PC[12] curr_PC[13]
+ curr_PC[14] curr_PC[15] curr_PC[16] curr_PC[17] curr_PC[18] curr_PC[19] curr_PC[1]
+ curr_PC[20] curr_PC[21] curr_PC[22] curr_PC[23] curr_PC[24] curr_PC[25] curr_PC[26]
+ curr_PC[27] curr_PC[2] curr_PC[3] curr_PC[4] curr_PC[5] curr_PC[6] curr_PC[7] curr_PC[8]
+ curr_PC[9] dest_idx[0] dest_idx[1] dest_idx[2] dest_idx[3] dest_idx[4] dest_idx[5]
+ dest_mask[0] dest_mask[1] dest_pred[0] dest_pred[1] dest_pred[2] dest_pred_val dest_val[0]
+ dest_val[10] dest_val[11] dest_val[12] dest_val[13] dest_val[14] dest_val[15] dest_val[16]
+ dest_val[17] dest_val[18] dest_val[19] dest_val[1] dest_val[20] dest_val[21] dest_val[22]
+ dest_val[23] dest_val[24] dest_val[25] dest_val[26] dest_val[27] dest_val[28] dest_val[29]
+ dest_val[2] dest_val[30] dest_val[31] dest_val[3] dest_val[4] dest_val[5] dest_val[6]
+ dest_val[7] dest_val[8] dest_val[9] instruction[0] instruction[10] instruction[11]
+ instruction[12] instruction[13] instruction[14] instruction[15] instruction[16]
+ instruction[17] instruction[18] instruction[19] instruction[1] instruction[20] instruction[21]
+ instruction[22] instruction[23] instruction[24] instruction[25] instruction[26]
+ instruction[27] instruction[28] instruction[29] instruction[2] instruction[30] instruction[31]
+ instruction[32] instruction[33] instruction[34] instruction[35] instruction[36]
+ instruction[37] instruction[38] instruction[39] instruction[3] instruction[40] instruction[41]
+ instruction[4] instruction[5] instruction[6] instruction[7] instruction[8] instruction[9]
+ int_return is_load is_store loadstore_address[0] loadstore_address[10] loadstore_address[11]
+ loadstore_address[12] loadstore_address[13] loadstore_address[14] loadstore_address[15]
+ loadstore_address[16] loadstore_address[17] loadstore_address[18] loadstore_address[19]
+ loadstore_address[1] loadstore_address[20] loadstore_address[21] loadstore_address[22]
+ loadstore_address[23] loadstore_address[24] loadstore_address[25] loadstore_address[26]
+ loadstore_address[27] loadstore_address[28] loadstore_address[29] loadstore_address[2]
+ loadstore_address[30] loadstore_address[31] loadstore_address[3] loadstore_address[4]
+ loadstore_address[5] loadstore_address[6] loadstore_address[7] loadstore_address[8]
+ loadstore_address[9] loadstore_dest[0] loadstore_dest[1] loadstore_dest[2] loadstore_dest[3]
+ loadstore_dest[4] loadstore_dest[5] loadstore_size[0] loadstore_size[1] new_PC[0]
+ new_PC[10] new_PC[11] new_PC[12] new_PC[13] new_PC[14] new_PC[15] new_PC[16] new_PC[17]
+ new_PC[18] new_PC[19] new_PC[1] new_PC[20] new_PC[21] new_PC[22] new_PC[23] new_PC[24]
+ new_PC[25] new_PC[26] new_PC[27] new_PC[2] new_PC[3] new_PC[4] new_PC[5] new_PC[6]
+ new_PC[7] new_PC[8] new_PC[9] pred_idx[0] pred_idx[1] pred_idx[2] pred_val reg1_idx[0]
+ reg1_idx[1] reg1_idx[2] reg1_idx[3] reg1_idx[4] reg1_idx[5] reg1_val[0] reg1_val[10]
+ reg1_val[11] reg1_val[12] reg1_val[13] reg1_val[14] reg1_val[15] reg1_val[16] reg1_val[17]
+ reg1_val[18] reg1_val[19] reg1_val[1] reg1_val[20] reg1_val[21] reg1_val[22] reg1_val[23]
+ reg1_val[24] reg1_val[25] reg1_val[26] reg1_val[27] reg1_val[28] reg1_val[29] reg1_val[2]
+ reg1_val[30] reg1_val[31] reg1_val[3] reg1_val[4] reg1_val[5] reg1_val[6] reg1_val[7]
+ reg1_val[8] reg1_val[9] reg2_idx[0] reg2_idx[1] reg2_idx[2] reg2_idx[3] reg2_idx[4]
+ reg2_idx[5] reg2_val[0] reg2_val[10] reg2_val[11] reg2_val[12] reg2_val[13] reg2_val[14]
+ reg2_val[15] reg2_val[16] reg2_val[17] reg2_val[18] reg2_val[19] reg2_val[1] reg2_val[20]
+ reg2_val[21] reg2_val[22] reg2_val[23] reg2_val[24] reg2_val[25] reg2_val[26] reg2_val[27]
+ reg2_val[28] reg2_val[29] reg2_val[2] reg2_val[30] reg2_val[31] reg2_val[3] reg2_val[4]
+ reg2_val[5] reg2_val[6] reg2_val[7] reg2_val[8] reg2_val[9] rst sign_extend take_branch
+ vccd1 vssd1 wb_clk_i
XFILLER_0_94_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06883_ reg1_idx[0] reg1_idx[1] reg1_idx[4] vssd1 vssd1 vccd1 vccd1 _06885_/C sky130_fd_sc_hd__and3_1
XFILLER_0_118_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09671_ _09669_/X _09670_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09671_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11866__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08622_ _09058_/A _09060_/A _09058_/B _08405_/Y _08370_/Y vssd1 vssd1 vccd1 vccd1
+ _09061_/B sky130_fd_sc_hd__o32ai_4
XFILLER_0_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08553_ _08538_/B _08552_/X _08551_/X _08542_/Y vssd1 vssd1 vccd1 vccd1 _08553_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08484_ _08484_/A _08484_/B vssd1 vssd1 vccd1 vccd1 _08485_/C sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout162_A _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11135__A _12255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07504_ _09452_/A _07504_/B vssd1 vssd1 vccd1 vccd1 _07506_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07435_ _09968_/A _07434_/X _06622_/X vssd1 vssd1 vccd1 vccd1 _07435_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07366_ fanout52/X fanout83/X fanout81/X fanout51/X vssd1 vssd1 vccd1 vccd1 _07367_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10693__B _12255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09105_ _09660_/B _10230_/A vssd1 vssd1 vccd1 vccd1 _12360_/A sky130_fd_sc_hd__xor2_2
X_07297_ _07087_/B _06939_/C _07165_/A vssd1 vssd1 vccd1 vccd1 _07300_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09036_ _08589_/A _08597_/A _08591_/X _09034_/A vssd1 vssd1 vccd1 vccd1 _09037_/B
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_32_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12897__A2 _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09762__A2 _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10109__B1 _12228_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ _09938_/A _09938_/B vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__or2_1
XANTENNA_fanout75_A _12768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09869_ _09869_/A _09869_/B vssd1 vssd1 vccd1 vccd1 _09870_/B sky130_fd_sc_hd__nor2_1
X_12880_ _13139_/A _13140_/A _13139_/B vssd1 vssd1 vccd1 vccd1 _13144_/B sky130_fd_sc_hd__a21bo_1
X_11900_ _11848_/X _11972_/D _11899_/Y vssd1 vssd1 vccd1 vccd1 _11900_/Y sky130_fd_sc_hd__a21oi_2
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _10518_/Y _11830_/Y _11831_/S vssd1 vssd1 vccd1 vccd1 _11831_/X sky130_fd_sc_hd__mux2_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _07052_/B _12250_/B _11761_/X vssd1 vssd1 vccd1 vccd1 _11762_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_68_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11693_ _12019_/A _11693_/B vssd1 vssd1 vccd1 vccd1 _11695_/B sky130_fd_sc_hd__xnor2_1
X_10713_ _10596_/A _10596_/B _10594_/Y vssd1 vssd1 vccd1 vccd1 _10720_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_125_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10644_ _09205_/B _10631_/X _10643_/X _10622_/X vssd1 vssd1 vccd1 vccd1 _10644_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10575_ fanout56/X fanout20/X fanout18/X fanout98/X vssd1 vssd1 vccd1 vccd1 _10576_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_51_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12314_ _12214_/A _12266_/A _12313_/B _12217_/X vssd1 vssd1 vccd1 vccd1 _12314_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_0_2_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13294_ _13296_/CLK _13294_/D vssd1 vssd1 vccd1 vccd1 hold295/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_121_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12245_ _09183_/Y _12235_/B _12244_/X _06591_/B _12243_/Y vssd1 vssd1 vccd1 vccd1
+ _12245_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12176_ reg1_val[27] curr_PC[27] vssd1 vssd1 vccd1 vccd1 _12176_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09753__A2 _07308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10899__B2 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10899__A1 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__A1 _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__B2 _07869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11127_ _12301_/A _10677_/B fanout8/X fanout52/X vssd1 vssd1 vccd1 vccd1 _11128_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11058_ _11058_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11060_/B sky130_fd_sc_hd__xnor2_1
X_10009_ _12762_/A fanout46/X fanout12/X _12760_/A vssd1 vssd1 vccd1 vccd1 _10010_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13065__A2 _13151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07819__A2 _07168_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12273__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07220_ _07221_/A _07221_/B vssd1 vssd1 vccd1 vccd1 _07220_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09079__B _09079_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07151_ _07128_/B _07128_/C _07128_/D _07135_/B vssd1 vssd1 vccd1 vccd1 _07153_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_77 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07082_ _11688_/A _10156_/B2 fanout69/X _10156_/A1 vssd1 vssd1 vccd1 vccd1 _07083_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout105 _07034_/Y vssd1 vssd1 vccd1 vccd1 _12760_/A sky130_fd_sc_hd__buf_8
Xfanout138 _12736_/A vssd1 vssd1 vccd1 vccd1 _07969_/A sky130_fd_sc_hd__clkbuf_8
Xfanout127 _07894_/A vssd1 vssd1 vccd1 vccd1 _08857_/A sky130_fd_sc_hd__buf_12
Xfanout116 _11780_/A vssd1 vssd1 vccd1 vccd1 _12019_/A sky130_fd_sc_hd__clkbuf_16
X_07984_ _07984_/A _07984_/B vssd1 vssd1 vccd1 vccd1 _07999_/A sky130_fd_sc_hd__nor2_2
Xfanout149 _12131_/A vssd1 vssd1 vccd1 vccd1 _11973_/A sky130_fd_sc_hd__buf_4
X_06935_ reg1_val[10] reg1_val[11] reg1_val[12] _07027_/B vssd1 vssd1 vccd1 vccd1
+ _07165_/B sky130_fd_sc_hd__or4_4
XANTENNA__11839__B1 _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09723_ _10306_/A _09723_/B vssd1 vssd1 vccd1 vccd1 _09725_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07507__A1 _10553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06866_ _06866_/A _10621_/A _10498_/A _06866_/D vssd1 vssd1 vccd1 vccd1 _06871_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__07507__B2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ _09655_/A _09655_/B vssd1 vssd1 vccd1 vccd1 _09654_/X sky130_fd_sc_hd__and2_1
XANTENNA__08180__B2 _08692_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08180__A1 _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07343__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08605_ _08568_/Y _08605_/B vssd1 vssd1 vccd1 vccd1 _09043_/B sky130_fd_sc_hd__and2b_1
X_06797_ _06996_/A reg1_val[6] vssd1 vssd1 vccd1 vccd1 _06797_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09585_ fanout57/X fanout46/X fanout12/X _07553_/A vssd1 vssd1 vccd1 vccd1 _09586_/B
+ sky130_fd_sc_hd__o22a_1
X_08536_ _08531_/A _08531_/C _08531_/B vssd1 vssd1 vccd1 vccd1 _08537_/C sky130_fd_sc_hd__a21oi_1
X_08467_ _08471_/A _08471_/B vssd1 vssd1 vccd1 vccd1 _08467_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_108_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08398_ _08432_/A _08397_/B _08390_/X vssd1 vssd1 vccd1 vccd1 _08407_/A sky130_fd_sc_hd__a21oi_1
X_07418_ _07624_/B _07624_/A vssd1 vssd1 vccd1 vccd1 _07418_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12016__B1 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07349_ _07349_/A _07349_/B vssd1 vssd1 vccd1 vccd1 _07421_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10042__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10360_ _10360_/A _10360_/B vssd1 vssd1 vccd1 vccd1 _10607_/A sky130_fd_sc_hd__xnor2_2
X_09019_ _09007_/X _09016_/X _08340_/A _09060_/A _08621_/B vssd1 vssd1 vccd1 vccd1
+ _09020_/B sky130_fd_sc_hd__a2111o_1
X_10291_ _10292_/A _10292_/B vssd1 vssd1 vccd1 vccd1 _10435_/A sky130_fd_sc_hd__or2_1
Xhold170 hold170/A vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
X_12030_ _12098_/A _12030_/B vssd1 vssd1 vccd1 vccd1 _12032_/C sky130_fd_sc_hd__nand2_1
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 hold226/X vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
X_12932_ _12946_/A hold169/X vssd1 vssd1 vccd1 vccd1 hold170/A sky130_fd_sc_hd__and2_1
X_12863_ _13107_/B _13108_/A _12806_/X vssd1 vssd1 vccd1 vccd1 _13113_/A sky130_fd_sc_hd__a21o_1
X_12794_ hold7/X hold254/X vssd1 vssd1 vccd1 vccd1 _12885_/A sky130_fd_sc_hd__and2b_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11814_ _11814_/A _11969_/A vssd1 vssd1 vccd1 vccd1 _11814_/Y sky130_fd_sc_hd__nor2_1
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11745_/A _11745_/B vssd1 vssd1 vccd1 vccd1 _11746_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11676_ _12200_/A _11676_/B vssd1 vssd1 vccd1 vccd1 _11680_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11222__B _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10627_ _09525_/X _09531_/X _11194_/S vssd1 vssd1 vccd1 vccd1 _10628_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_3_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09423__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09423__A1 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10558_ _07308_/A _07308_/B fanout62/X vssd1 vssd1 vccd1 vccd1 _10559_/C sky130_fd_sc_hd__a21o_1
XANTENNA__09908__A _10819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13277_ _13277_/CLK _13277_/D vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11781__A2 _06987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12228_ _06605_/B _12227_/X _12228_/B1 vssd1 vssd1 vccd1 vccd1 _12228_/Y sky130_fd_sc_hd__o21ai_1
X_10489_ _10232_/Y _10732_/A _10488_/Y vssd1 vssd1 vccd1 vccd1 _10961_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12191__C1 _12382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11533__A2 _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__B _07148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12159_ _12159_/A vssd1 vssd1 vccd1 vccd1 _12161_/A sky130_fd_sc_hd__inv_2
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06720_ reg1_val[11] _07018_/A vssd1 vssd1 vccd1 vccd1 _06722_/B sky130_fd_sc_hd__and2_1
X_06651_ _06649_/Y _06680_/B1 _06778_/B reg2_val[20] vssd1 vssd1 vccd1 vccd1 _06653_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_06582_ reg2_val[29] _06752_/A _06688_/B1 _06581_/Y vssd1 vssd1 vccd1 vccd1 _07243_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_93_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09370_ _09355_/X _09369_/X _11195_/A vssd1 vssd1 vccd1 vccd1 _09370_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_115_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08321_ _08345_/A _08345_/B _08317_/Y vssd1 vssd1 vccd1 vccd1 _08334_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_86_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08465__A2 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13104__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08252_ _08250_/A _08250_/B _08251_/X vssd1 vssd1 vccd1 vccd1 _08294_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07673__B1 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10272__A2 _10269_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11413__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07203_ fanout77/X _07058_/A fanout62/X _08532_/B vssd1 vssd1 vccd1 vccd1 _07204_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_222 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_767 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08183_ _08183_/A _08183_/B vssd1 vssd1 vccd1 vccd1 _08245_/B sky130_fd_sc_hd__xor2_1
XANTENNA_fanout125_A _07319_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09414__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09414__A1 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07134_ _07134_/A reg1_val[1] vssd1 vssd1 vccd1 vccd1 _07869_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_15_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10024__A2 _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06779__A2 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07065_ _07066_/A _07066_/B vssd1 vssd1 vccd1 vccd1 _07065_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12182__C1 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07967_ _07968_/B vssd1 vssd1 vccd1 vccd1 _07967_/Y sky130_fd_sc_hd__inv_2
X_09706_ _06768_/Y _09191_/X _09383_/B _06868_/D _09705_/X vssd1 vssd1 vccd1 vccd1
+ _09706_/X sky130_fd_sc_hd__o221a_1
X_06918_ _09198_/C instruction[5] _09188_/C vssd1 vssd1 vccd1 vccd1 _06918_/X sky130_fd_sc_hd__or3_2
XANTENNA__06896__B _06897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07898_ _07892_/A _07892_/B _07897_/B _08053_/A _08053_/B vssd1 vssd1 vccd1 vccd1
+ _07928_/A sky130_fd_sc_hd__o32a_1
X_06849_ _12357_/A _06847_/X _06848_/Y _06833_/Y vssd1 vssd1 vccd1 vccd1 _06849_/X
+ sky130_fd_sc_hd__o211a_1
X_09637_ _09637_/A _09637_/B vssd1 vssd1 vccd1 vccd1 _09638_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09568_ _09569_/A _09569_/B vssd1 vssd1 vccd1 vccd1 _09570_/A sky130_fd_sc_hd__or2_1
XFILLER_0_93_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08519_ _08540_/A _08540_/B _08516_/C vssd1 vssd1 vccd1 vccd1 _08520_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_93_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12419__A _12588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11323__A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09499_ _09500_/B _09500_/A vssd1 vssd1 vccd1 vccd1 _09499_/Y sky130_fd_sc_hd__nand2b_1
X_11530_ _11439_/A _11439_/B _11438_/A vssd1 vssd1 vccd1 vccd1 _11540_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11461_ _11276_/Y _11636_/A _11459_/Y vssd1 vssd1 vccd1 vccd1 _11461_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13200_ _13296_/CLK hold67/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
X_11392_ _11197_/S _11390_/X _11391_/X _06917_/Y vssd1 vssd1 vccd1 vccd1 _11404_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10412_ _12776_/A fanout52/X _10677_/B _11935_/A vssd1 vssd1 vccd1 vccd1 _10413_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09728__A _10301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12960__B2 _12980_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13131_ _13131_/A _13131_/B vssd1 vssd1 vccd1 vccd1 _13131_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10343_ _10209_/A _10209_/B _10193_/A vssd1 vssd1 vccd1 vccd1 _10353_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13062_ _13062_/A _13062_/B vssd1 vssd1 vccd1 vccd1 _13063_/B sky130_fd_sc_hd__nand2_1
X_10274_ _10523_/A _10523_/B _12278_/A vssd1 vssd1 vccd1 vccd1 _10274_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07307__A_N _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ _12776_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _12014_/B sky130_fd_sc_hd__or2_1
XANTENNA__06942__A2 _07087_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12915_ hold205/X _12947_/A2 _12947_/B1 hold219/X vssd1 vssd1 vccd1 vccd1 hold220/A
+ sky130_fd_sc_hd__a22o_1
X_12846_ _13062_/A _13063_/A _13062_/B vssd1 vssd1 vccd1 vccd1 _13068_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__12228__B1 _12228_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12779__A1 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12777_ hold17/X _12778_/B _12776_/Y _13147_/A vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__o211a_1
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06972__D _07001_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11233__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11728_ _11376_/B _11552_/B _11725_/Y _11727_/X vssd1 vssd1 vccd1 vccd1 _11729_/B
+ sky130_fd_sc_hd__a31o_1
X_11659_ hold234/A _11559_/A _11657_/X _11920_/C1 vssd1 vssd1 vccd1 vccd1 _11659_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13329_ instruction[10] vssd1 vssd1 vccd1 vccd1 pred_idx[2] sky130_fd_sc_hd__buf_12
XFILLER_0_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11506__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08870_ _08870_/A _08870_/B vssd1 vssd1 vccd1 vccd1 _08872_/B sky130_fd_sc_hd__nor2_2
X_07821_ _09180_/A _07821_/B _07821_/C vssd1 vssd1 vccd1 vccd1 _07824_/B sky130_fd_sc_hd__and3_1
X_07752_ _07751_/A _07785_/A vssd1 vssd1 vccd1 vccd1 _07753_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_79_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06703_ reg1_val[14] _07192_/A vssd1 vssd1 vccd1 vccd1 _06704_/B sky130_fd_sc_hd__and2_1
X_07683_ _08812_/A _08812_/B vssd1 vssd1 vccd1 vccd1 _08813_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09883__A1 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06634_ _06641_/A _12598_/B vssd1 vssd1 vccd1 vccd1 _06634_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09883__B2 _07098_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ _09232_/A _09232_/B _09237_/A vssd1 vssd1 vccd1 vccd1 _09437_/A sky130_fd_sc_hd__o21ai_2
X_09353_ _09351_/X _09352_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09353_/X sky130_fd_sc_hd__mux2_1
X_06565_ instruction[0] instruction[1] instruction[2] pred_val vssd1 vssd1 vccd1 vccd1
+ _06567_/B sky130_fd_sc_hd__or4bb_4
X_08304_ _08775_/A _08304_/B vssd1 vssd1 vccd1 vccd1 _08309_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11978__C1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07646__B1 _07182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09284_ _07525_/A _07525_/B _07523_/Y vssd1 vssd1 vccd1 vccd1 _09288_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_35_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08235_ _08235_/A _08235_/B vssd1 vssd1 vccd1 vccd1 _08285_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08166_ _08166_/A _08166_/B vssd1 vssd1 vccd1 vccd1 _08207_/A sky130_fd_sc_hd__nand2_2
X_07117_ _09898_/A _09764_/A _07115_/X vssd1 vssd1 vccd1 vccd1 _07117_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_43_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08097_ _07969_/A _08348_/B fanout56/X _12734_/A vssd1 vssd1 vccd1 vccd1 _08098_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07068__A _07068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07048_ _08532_/B vssd1 vssd1 vccd1 vccd1 _09252_/A sky130_fd_sc_hd__inv_2
XFILLER_0_100_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07177__A2 _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__A _09283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06924__A2 _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _09507_/B _09660_/B _08998_/X _09509_/C _09509_/B vssd1 vssd1 vccd1 vccd1
+ _09000_/B sky130_fd_sc_hd__o32a_1
XANTENNA__08126__B2 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10961_ _10960_/Y _10961_/B vssd1 vssd1 vccd1 vccd1 _10961_/Y sky130_fd_sc_hd__nand2b_1
X_12700_ _12700_/A _12700_/B _12700_/C vssd1 vssd1 vccd1 vccd1 _12701_/B sky130_fd_sc_hd__and3_2
XANTENNA__07531__A _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12631_ reg1_val[14] _12632_/B vssd1 vssd1 vccd1 vccd1 _12639_/A sky130_fd_sc_hd__nand2_1
X_10892_ _11429_/A _10892_/B vssd1 vssd1 vccd1 vccd1 _10894_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12562_ reg1_val[1] _12563_/B vssd1 vssd1 vccd1 vccd1 _12564_/A sky130_fd_sc_hd__or2_1
XFILLER_0_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12493_ _12551_/A _12493_/B vssd1 vssd1 vccd1 vccd1 _12500_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_81_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10892__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11513_ _11513_/A _11513_/B vssd1 vssd1 vccd1 vccd1 _11514_/B sky130_fd_sc_hd__and2_1
X_11444_ _11444_/A _11444_/B _11442_/Y vssd1 vssd1 vccd1 vccd1 _11445_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11375_ _10965_/B _11374_/Y _11373_/Y vssd1 vssd1 vccd1 vccd1 _11376_/B sky130_fd_sc_hd__o21ai_2
X_13114_ hold289/A _13113_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13114_/X sky130_fd_sc_hd__mux2_1
X_10326_ _10326_/A _10326_/B vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__nand2_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ hold284/X _12721_/B _13044_/X _12722_/A vssd1 vssd1 vccd1 vccd1 hold285/A
+ sky130_fd_sc_hd__a22o_1
X_10257_ _09385_/C _10514_/C hold292/A vssd1 vssd1 vccd1 vccd1 _10257_/Y sky130_fd_sc_hd__a21oi_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06680__A2_N _06569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10188_ _10346_/A _10188_/B vssd1 vssd1 vccd1 vccd1 _10190_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11228__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13110__B2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08668__A2 _10811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07340__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12829_ hold240/X hold45/X vssd1 vssd1 vccd1 vccd1 _12830_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_84_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11424__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11424__A1 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13177__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08020_ _08020_/A _08020_/B vssd1 vssd1 vccd1 vccd1 _08023_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08272__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout7 fanout7/A vssd1 vssd1 vccd1 vccd1 fanout7/X sky130_fd_sc_hd__buf_6
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09971_ _10750_/S _09528_/X _11195_/C vssd1 vssd1 vccd1 vccd1 _09971_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08922_ _08922_/A _08922_/B vssd1 vssd1 vccd1 vccd1 _08923_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_110_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08356__B2 _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08356__A1 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09553__B1 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ _08853_/A _08853_/B vssd1 vssd1 vccd1 vccd1 _08861_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07804_ _07804_/A _07804_/B vssd1 vssd1 vccd1 vccd1 _08020_/A sky130_fd_sc_hd__nor2_2
X_08784_ _08784_/A _08784_/B vssd1 vssd1 vccd1 vccd1 _08785_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07735_ _08841_/A1 _08217_/B fanout55/X _08841_/B2 vssd1 vssd1 vccd1 vccd1 _07736_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08659__A2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07666_ _07687_/B _08904_/A _07687_/A vssd1 vssd1 vccd1 vccd1 _07688_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__07331__A2 _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09405_ _09323_/A _09323_/B _09324_/Y vssd1 vssd1 vccd1 vccd1 _09503_/A sky130_fd_sc_hd__o21ai_4
X_06617_ _06619_/A vssd1 vssd1 vccd1 vccd1 _06617_/Y sky130_fd_sc_hd__inv_2
X_07597_ _07604_/B vssd1 vssd1 vccd1 vccd1 _07597_/Y sky130_fd_sc_hd__inv_2
X_06548_ instruction[0] pred_val vssd1 vssd1 vccd1 vccd1 _06881_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_118_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09336_ _09224_/X _09559_/C _09335_/Y vssd1 vssd1 vccd1 vccd1 _09336_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09267_ _09267_/A _09267_/B vssd1 vssd1 vccd1 vccd1 _09271_/A sky130_fd_sc_hd__xor2_1
X_08218_ _08857_/A _08218_/B vssd1 vssd1 vccd1 vccd1 _08283_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09278__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09198_ instruction[4] _09198_/B _09198_/C _09200_/B vssd1 vssd1 vccd1 vccd1 _09198_/X
+ sky130_fd_sc_hd__and4_2
X_08149_ _08149_/A _08149_/B vssd1 vssd1 vccd1 vccd1 _08153_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11160_ _11160_/A _11160_/B vssd1 vssd1 vccd1 vccd1 _11162_/B sky130_fd_sc_hd__xnor2_1
X_10111_ _10251_/S _10110_/X _09214_/A vssd1 vssd1 vccd1 vccd1 _10111_/Y sky130_fd_sc_hd__o21ai_2
X_11091_ _10251_/S _09395_/Y _11090_/X vssd1 vssd1 vccd1 vccd1 _11092_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__12432__A _12598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10042_ _10677_/A fanout98/X fanout56/X fanout58/X vssd1 vssd1 vccd1 vccd1 _10043_/B
+ sky130_fd_sc_hd__o22a_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ _12124_/B _12059_/B hold173/A vssd1 vssd1 vccd1 vccd1 _11995_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08357__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07261__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10944_ _10942_/X _10944_/B vssd1 vssd1 vccd1 vccd1 _10945_/B sky130_fd_sc_hd__and2b_1
X_10875_ _11559_/A _10983_/B hold195/A vssd1 vssd1 vccd1 vccd1 _10875_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12614_ reg1_val[11] _12614_/B vssd1 vssd1 vccd1 vccd1 _12615_/B sky130_fd_sc_hd__or2_1
X_12545_ _12551_/A _12545_/B vssd1 vssd1 vccd1 vccd1 _12546_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11511__A _11511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12476_ _12485_/A _12476_/B vssd1 vssd1 vccd1 vccd1 _12478_/C sky130_fd_sc_hd__nand2_1
XANTENNA_5 _11092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11427_ _11427_/A _11427_/B vssd1 vssd1 vccd1 vccd1 _11428_/B sky130_fd_sc_hd__or2_1
XFILLER_0_111_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08586__B2 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08586__A1 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ _11358_/A _11358_/B vssd1 vssd1 vccd1 vccd1 _11360_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09783__B1 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08820__A _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ _10461_/B _10309_/B vssd1 vssd1 vccd1 vccd1 _10311_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11590__B1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11289_ _11289_/A _11289_/B vssd1 vssd1 vccd1 vccd1 _11289_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_67_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ _13028_/A _13028_/B vssd1 vssd1 vccd1 vccd1 _13282_/D sky130_fd_sc_hd__and2_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09073__D _09073_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07520_ _09618_/B2 _12782_/A fanout22/X _09618_/A1 vssd1 vssd1 vccd1 vccd1 _07521_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10797__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07171__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08510__A1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08510__B2 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07451_ _07451_/A _07451_/B vssd1 vssd1 vccd1 vccd1 _07464_/B sky130_fd_sc_hd__xnor2_4
X_07382_ _07385_/A _07385_/B vssd1 vssd1 vccd1 vccd1 _07382_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_45_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09121_ _09119_/X _09120_/X _09359_/S vssd1 vssd1 vccd1 vccd1 _09121_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09052_ _09052_/A _09052_/B vssd1 vssd1 vccd1 vccd1 _10617_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08003_ _07738_/B _07738_/C _07738_/A vssd1 vssd1 vccd1 vccd1 _08007_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_13_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout205_A _08311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09774__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08730__A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09954_ _09954_/A _09954_/B vssd1 vssd1 vccd1 vccd1 _09955_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_110_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08905_ _07686_/A _07685_/C _08813_/A vssd1 vssd1 vccd1 vccd1 _08908_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_57_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07346__A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11333__B1 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09885_ _12736_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _09887_/B sky130_fd_sc_hd__or2_1
X_08836_ _08836_/A _08836_/B vssd1 vssd1 vccd1 vccd1 _08840_/A sky130_fd_sc_hd__xnor2_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08767_ _08870_/B _08767_/B vssd1 vssd1 vccd1 vccd1 _08768_/C sky130_fd_sc_hd__or2_1
XANTENNA__09829__A1 _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08698_ _08699_/B _08699_/A vssd1 vssd1 vccd1 vccd1 _08698_/X sky130_fd_sc_hd__and2b_1
X_07718_ _08855_/A _07718_/B vssd1 vssd1 vccd1 vccd1 _07722_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10439__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07649_ _08888_/A _08888_/B vssd1 vssd1 vccd1 vccd1 _08889_/A sky130_fd_sc_hd__or2_1
XFILLER_0_94_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10660_ _10660_/A _10660_/B vssd1 vssd1 vccd1 vccd1 _10662_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout20_A _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09319_ _09320_/A _09320_/B vssd1 vssd1 vccd1 vccd1 _09319_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08265__B1 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10591_ _10418_/A _10418_/B _10421_/A vssd1 vssd1 vccd1 vccd1 _10596_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_118_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12330_ _13246_/Q _12330_/B vssd1 vssd1 vccd1 vccd1 _12332_/C sky130_fd_sc_hd__or2_1
XFILLER_0_63_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12261_ _12204_/A _12204_/B _12201_/Y vssd1 vssd1 vccd1 vccd1 _12263_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11212_ curr_PC[15] _11213_/B vssd1 vssd1 vccd1 vccd1 _11212_/Y sky130_fd_sc_hd__nor2_1
X_12192_ _06612_/B _12243_/B1 _12190_/Y _06610_/Y _12191_/X vssd1 vssd1 vccd1 vccd1
+ _12192_/Y sky130_fd_sc_hd__o221ai_4
XANTENNA__10989__A1_N _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ _11262_/B _11143_/B _11143_/C vssd1 vssd1 vccd1 vccd1 _11143_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__07256__A _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11074_ _12278_/A _11000_/X _11215_/C vssd1 vssd1 vccd1 vccd1 _11076_/A sky130_fd_sc_hd__a21oi_1
X_10025_ _10559_/A _10025_/B vssd1 vssd1 vccd1 vccd1 _10027_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07543__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ _09075_/Y _09076_/Y _12131_/A vssd1 vssd1 vccd1 vccd1 _11977_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_53_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10410__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10927_ _10927_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _10928_/B sky130_fd_sc_hd__or2_1
XFILLER_0_128_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10858_ _10740_/B _10740_/C _12131_/A vssd1 vssd1 vccd1 vccd1 _10859_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10789_ _10789_/A _10789_/B vssd1 vssd1 vccd1 vccd1 _10793_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_124_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12528_ _12513_/B _12521_/B _12551_/A vssd1 vssd1 vccd1 vccd1 _12541_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_124_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12459_ reg1_val[12] curr_PC[12] _12487_/S vssd1 vssd1 vccd1 vccd1 _12461_/B sky130_fd_sc_hd__mux2_1
XANTENNA__06989__B _11782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10118__A1 _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _10752_/S _07135_/B _06951_/C vssd1 vssd1 vccd1 vccd1 _08544_/B sky130_fd_sc_hd__or3_2
XANTENNA__11315__B1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _09345_/X _09348_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09670_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11866__A1 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06990__B1 _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ _08621_/A _08621_/B vssd1 vssd1 vccd1 vccd1 _09058_/B sky130_fd_sc_hd__or2_2
X_06882_ _06915_/B dest_pred_val _12345_/A vssd1 vssd1 vccd1 vccd1 take_branch sky130_fd_sc_hd__a21o_4
XANTENNA__11866__B2 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08552_ _08538_/A _08537_/C _08537_/B vssd1 vssd1 vccd1 vccd1 _08552_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_89_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08483_ _08502_/B _08502_/A vssd1 vssd1 vccd1 vccd1 _08485_/B sky130_fd_sc_hd__and2b_1
X_07503_ _10156_/B2 _10557_/A fanout62/X _10156_/A1 vssd1 vssd1 vccd1 vccd1 _07504_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07434_ _07434_/A _07434_/B _07434_/C _07434_/D vssd1 vssd1 vccd1 vccd1 _07434_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_43_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07365_ _07626_/A _07626_/B _07361_/Y vssd1 vssd1 vccd1 vccd1 _07376_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09104_ _09095_/X _09102_/Y _09103_/X _09085_/X _09101_/X vssd1 vssd1 vccd1 vccd1
+ _10230_/A sky130_fd_sc_hd__o221a_2
X_07296_ _07601_/B _07294_/B _07420_/B _07295_/B _07295_/A vssd1 vssd1 vccd1 vccd1
+ _07353_/A sky130_fd_sc_hd__o32a_2
XFILLER_0_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09035_ _09514_/A _09035_/B vssd1 vssd1 vccd1 vccd1 _09668_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07773__A2 _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ _09938_/A _09938_/B vssd1 vssd1 vccd1 vccd1 _09939_/A sky130_fd_sc_hd__nand2_1
XANTENNA_fanout68_A _07090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09868_ _09869_/A _09869_/B vssd1 vssd1 vccd1 vccd1 _09870_/A sky130_fd_sc_hd__and2_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08819_ _09772_/A _08681_/A _09295_/A _08819_/B2 vssd1 vssd1 vccd1 vccd1 _08820_/B
+ sky130_fd_sc_hd__o22a_1
X_09799_ _09577_/A _09577_/B _09576_/A vssd1 vssd1 vccd1 vccd1 _09804_/A sky130_fd_sc_hd__a21o_2
X_11830_ _11830_/A _11830_/B vssd1 vssd1 vccd1 vccd1 _11830_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__10230__A _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11761_ _11733_/Y _11735_/X _11760_/X _06930_/Y vssd1 vssd1 vccd1 vccd1 _11761_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10712_ _10589_/A _10589_/B _10572_/Y vssd1 vssd1 vccd1 vccd1 _10722_/A sky130_fd_sc_hd__a21bo_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11692_ fanout29/X _12203_/A fanout19/X fanout32/X vssd1 vssd1 vccd1 vccd1 _11693_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10643_ _09184_/X _10629_/X _10642_/Y _09115_/X _10641_/X vssd1 vssd1 vccd1 vccd1
+ _10643_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_91_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09986__B1 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10574_ _10435_/A _10435_/C _10435_/B vssd1 vssd1 vccd1 vccd1 _10588_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_121_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12313_ _12313_/A _12313_/B vssd1 vssd1 vccd1 vccd1 _12313_/Y sky130_fd_sc_hd__nor2_1
X_13293_ _13296_/CLK _13293_/D vssd1 vssd1 vccd1 vccd1 hold274/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12244_ _06591_/A _09194_/Y _10638_/B vssd1 vssd1 vccd1 vccd1 _12244_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_121_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08410__B1 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12175_ _12112_/X _12113_/Y _12115_/Y vssd1 vssd1 vccd1 vccd1 _12179_/A sky130_fd_sc_hd__o21a_1
XANTENNA__09185__B _09199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10899__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ _11126_/A _11126_/B vssd1 vssd1 vccd1 vccd1 _11129_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_64_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11057_ _11058_/A _11058_/B vssd1 vssd1 vccd1 vccd1 _11167_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__10520__A1 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10008_ _10306_/A _10008_/B vssd1 vssd1 vccd1 vccd1 _10012_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11959_ _12036_/A _11959_/B vssd1 vssd1 vccd1 vccd1 _11961_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_117_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07150_ _07150_/A _07150_/B vssd1 vssd1 vccd1 vccd1 _07150_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_82_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07081_ _10458_/A _07073_/A _07080_/X vssd1 vssd1 vccd1 vccd1 _07081_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08280__A _10819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10315__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout106 _10452_/B2 vssd1 vssd1 vccd1 vccd1 _08420_/B sky130_fd_sc_hd__clkbuf_8
Xfanout117 _07364_/A vssd1 vssd1 vccd1 vccd1 _11780_/A sky130_fd_sc_hd__buf_4
X_07983_ _07982_/B _07982_/C _07982_/A vssd1 vssd1 vccd1 vccd1 _07984_/B sky130_fd_sc_hd__a21oi_1
Xfanout139 _07004_/X vssd1 vssd1 vccd1 vccd1 _12736_/A sky130_fd_sc_hd__buf_8
X_09722_ _08680_/B fanout83/X fanout81/X fanout30/X vssd1 vssd1 vccd1 vccd1 _09723_/B
+ sky130_fd_sc_hd__o22a_1
X_06934_ reg1_val[7] reg1_val[8] reg1_val[9] _07038_/B vssd1 vssd1 vccd1 vccd1 _07027_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07507__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06865_ _06865_/A _06865_/B _06865_/C _11289_/A vssd1 vssd1 vccd1 vccd1 _06872_/C
+ sky130_fd_sc_hd__nor4_1
XANTENNA__09901__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09653_ _09653_/A _09653_/B vssd1 vssd1 vccd1 vccd1 _09655_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08180__A2 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08604_ _08605_/B _09043_/A _08568_/Y vssd1 vssd1 vccd1 vccd1 _09045_/A sky130_fd_sc_hd__a21o_1
X_09584_ _09584_/A _09584_/B vssd1 vssd1 vccd1 vccd1 _09588_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06730__A3 _12607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06796_ _09970_/A _06794_/Y _06795_/Y vssd1 vssd1 vccd1 vccd1 _06796_/X sky130_fd_sc_hd__o21a_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _10155_/A _08541_/B _08541_/A vssd1 vssd1 vccd1 vccd1 _08537_/B sky130_fd_sc_hd__mux2_1
XANTENNA__08468__B1 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08466_ _08595_/A _08466_/B vssd1 vssd1 vccd1 vccd1 _08471_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07140__B1 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08397_ _08390_/X _08397_/B vssd1 vssd1 vccd1 vccd1 _08432_/B sky130_fd_sc_hd__nand2b_1
X_07417_ _07417_/A _07417_/B vssd1 vssd1 vccd1 vccd1 _07624_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10290__A3 _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12016__A1 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12016__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07348_ _07344_/A _07344_/B _07388_/A vssd1 vssd1 vccd1 vccd1 _07421_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07279_ _07279_/A _07279_/B vssd1 vssd1 vccd1 vccd1 _08681_/B sky130_fd_sc_hd__xnor2_4
X_09018_ _08339_/A _08339_/B _09006_/X vssd1 vssd1 vccd1 vccd1 _09020_/A sky130_fd_sc_hd__a21o_1
X_10290_ _10458_/A _07073_/A _12349_/A _10289_/Y vssd1 vssd1 vccd1 vccd1 _10292_/B
+ sky130_fd_sc_hd__a31o_2
XANTENNA__09286__A _12349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold171 hold298/X vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__clkbuf_2
Xhold160 hold160/A vssd1 vssd1 vccd1 vccd1 hold160/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__A1 _12228_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 hold193/A vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12440__A _12603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12931_ hold168/X _13146_/B2 _12947_/B1 _13236_/Q vssd1 vssd1 vccd1 vccd1 hold169/A
+ sky130_fd_sc_hd__a22o_1
X_12862_ _13102_/A _13103_/A _13102_/B vssd1 vssd1 vccd1 vccd1 _13108_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_87_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11813_ _11634_/Y _11969_/A _11811_/X vssd1 vssd1 vccd1 vccd1 _11813_/Y sky130_fd_sc_hd__o21ai_1
X_12793_ hold270/X hold21/X vssd1 vssd1 vccd1 vccd1 _13157_/A sky130_fd_sc_hd__nand2b_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _11652_/B _11654_/B _11652_/A vssd1 vssd1 vccd1 vccd1 _11745_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_56_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11675_ _12772_/A fanout15/X fanout6/X _11794_/A vssd1 vssd1 vccd1 vccd1 _11676_/B
+ sky130_fd_sc_hd__o22a_1
X_10626_ _10504_/A _10501_/Y _10503_/B vssd1 vssd1 vccd1 vccd1 _10630_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09423__A2 _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10557_ _10557_/A _10557_/B vssd1 vssd1 vccd1 vccd1 _10559_/B sky130_fd_sc_hd__or2_1
X_13276_ _13277_/CLK hold94/X vssd1 vssd1 vccd1 vccd1 hold142/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11781__A3 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10488_ _10225_/X _10358_/X _10359_/X vssd1 vssd1 vccd1 vccd1 _10488_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12227_ _12322_/S _12226_/Y _12225_/Y vssd1 vssd1 vccd1 vccd1 _12227_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08934__A1 _08932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07198__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12191__B1 _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11533__A3 _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__A _10180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ _12160_/A _12160_/B _12160_/C vssd1 vssd1 vccd1 vccd1 _12159_/A sky130_fd_sc_hd__a21o_1
Xclkbuf_4_12_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13310_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11109_ _12005_/A _11213_/B _11108_/Y _11106_/X vssd1 vssd1 vccd1 vccd1 dest_val[14]
+ sky130_fd_sc_hd__o31ai_4
X_12089_ _12090_/A _12090_/B vssd1 vssd1 vccd1 vccd1 _12160_/A sky130_fd_sc_hd__nand2_1
X_06650_ reg2_val[20] _06729_/B _06680_/B1 _06649_/Y vssd1 vssd1 vccd1 vccd1 _07068_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06712__A3 _12626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06581_ _06687_/A _12632_/B vssd1 vssd1 vccd1 vccd1 _06581_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09111__A1 _09559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08320_ _08320_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _08345_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08251_ _08261_/B _08261_/A vssd1 vssd1 vccd1 vccd1 _08251_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07673__A1 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07673__B2 _07119_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07202_ _10658_/A _07202_/B vssd1 vssd1 vccd1 vccd1 _07205_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10009__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08182_ _08245_/A vssd1 vssd1 vccd1 vccd1 _08182_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_55_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09414__A2 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07133_ _07134_/A _12563_/A vssd1 vssd1 vccd1 vccd1 _08544_/C sky130_fd_sc_hd__and2_4
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07064_ _09610_/A _07064_/B vssd1 vssd1 vccd1 vccd1 _07066_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06779__A3 _12568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout118_A _07364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10980__A1 _11194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10045__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ _08777_/A _07966_/B vssd1 vssd1 vccd1 vccd1 _07968_/B sky130_fd_sc_hd__xnor2_1
X_09705_ _06964_/A _12250_/B _12243_/B1 _06771_/B _09704_/X vssd1 vssd1 vccd1 vccd1
+ _09705_/X sky130_fd_sc_hd__o221a_1
X_06917_ _09198_/C instruction[5] _09188_/C vssd1 vssd1 vccd1 vccd1 _06917_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07897_ _07897_/A _07897_/B vssd1 vssd1 vccd1 vccd1 _08053_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09636_ _09637_/A _09637_/B vssd1 vssd1 vccd1 vccd1 _09636_/Y sky130_fd_sc_hd__nand2_1
X_06848_ reg1_val[31] _06622_/X _09200_/A vssd1 vssd1 vccd1 vccd1 _06848_/Y sky130_fd_sc_hd__a21oi_1
X_06779_ _06783_/A _06649_/A _12568_/B _06778_/X vssd1 vssd1 vccd1 vccd1 _09679_/S
+ sky130_fd_sc_hd__a31oi_4
X_09567_ _10306_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _09569_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_81_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08518_ _10155_/A _08518_/B vssd1 vssd1 vccd1 vccd1 _08520_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11604__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09498_ _09498_/A _09498_/B vssd1 vssd1 vccd1 vccd1 _09500_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08449_ _08773_/A _08449_/B vssd1 vssd1 vccd1 vccd1 _08487_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11996__B1 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11460_ _11460_/A _11550_/A vssd1 vssd1 vccd1 vccd1 _11636_/A sky130_fd_sc_hd__or2_1
XFILLER_0_123_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11391_ _11831_/S _11391_/B vssd1 vssd1 vccd1 vccd1 _11391_/X sky130_fd_sc_hd__or2_1
XFILLER_0_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10411_ _10411_/A _10411_/B vssd1 vssd1 vccd1 vccd1 _10415_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13130_ _13130_/A _13130_/B vssd1 vssd1 vccd1 vccd1 _13131_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10342_ _10342_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _10356_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_21_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13061_ _13066_/A hold269/X vssd1 vssd1 vccd1 vccd1 _13289_/D sky130_fd_sc_hd__and2_1
XFILLER_0_104_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07719__A2 _11222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12173__B1 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10273_ _10235_/Y _10273_/B _10273_/C _10273_/D vssd1 vssd1 vccd1 vccd1 _10523_/B
+ sky130_fd_sc_hd__nand4b_2
X_12012_ _12012_/A _12012_/B vssd1 vssd1 vccd1 vccd1 _12014_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09744__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06942__A3 _07086_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07264__A _10180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12914_ _12946_/A hold206/X vssd1 vssd1 vccd1 vccd1 _13227_/D sky130_fd_sc_hd__and2_1
X_12845_ hold63/X hold268/X vssd1 vssd1 vccd1 vccd1 _13062_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__12779__A2 _12781_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12776_ _12776_/A _12778_/B vssd1 vssd1 vccd1 vccd1 _12776_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10239__B1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11727_ _11549_/X _11725_/Y _11894_/A vssd1 vssd1 vccd1 vccd1 _11727_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08852__B1 _07197_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11658_ _12187_/A1 _11657_/X hold234/A vssd1 vssd1 vccd1 vccd1 _11658_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12345__A _12345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11589_ _11540_/A _11540_/B _11538_/Y vssd1 vssd1 vccd1 vccd1 _11629_/A sky130_fd_sc_hd__a21o_1
X_10609_ _09816_/X _10609_/B _10609_/C _10850_/A vssd1 vssd1 vccd1 vccd1 _10609_/Y
+ sky130_fd_sc_hd__nand4b_2
X_13328_ instruction[9] vssd1 vssd1 vccd1 vccd1 pred_idx[1] sky130_fd_sc_hd__buf_12
XFILLER_0_107_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12951__A2 _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13259_ _13264_/CLK _13259_/D vssd1 vssd1 vccd1 vccd1 hold144/A sky130_fd_sc_hd__dfxtp_1
X_07820_ _08775_/A _07820_/B vssd1 vssd1 vccd1 vccd1 _07825_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07751_ _07751_/A _07751_/B _07749_/X vssd1 vssd1 vccd1 vccd1 _07785_/A sky130_fd_sc_hd__or3b_1
X_06702_ reg1_val[14] _07192_/A vssd1 vssd1 vccd1 vccd1 _06702_/X sky130_fd_sc_hd__or2_1
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07682_ _09452_/A _07682_/B vssd1 vssd1 vccd1 vccd1 _08812_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09883__A2 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06633_ instruction[33] _06633_/B vssd1 vssd1 vccd1 vccd1 _12598_/B sky130_fd_sc_hd__and2_4
XFILLER_0_126_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07902__A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09421_ _09421_/A _09421_/B vssd1 vssd1 vccd1 vccd1 _09489_/A sky130_fd_sc_hd__xnor2_4
X_06564_ instruction[15] _06552_/X _06563_/X _06633_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[4]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_87_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09352_ _09142_/X _09162_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09352_/X sky130_fd_sc_hd__mux2_1
X_08303_ _10281_/A _08572_/B _07117_/Y _10149_/A vssd1 vssd1 vccd1 vccd1 _08304_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07646__A1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout235_A _09384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07646__B2 _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09283_ _09283_/A _09775_/A vssd1 vssd1 vccd1 vccd1 _09289_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08234_ _08773_/A _08234_/B vssd1 vssd1 vccd1 vccd1 _08235_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08733__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10650__B1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08165_ _08165_/A _08165_/B vssd1 vssd1 vccd1 vccd1 _08166_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09399__A1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12255__A _12255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07116_ _09898_/A _09764_/A _07115_/X vssd1 vssd1 vccd1 vccd1 _07116_/X sky130_fd_sc_hd__o21a_1
X_08096_ _08857_/A _08096_/B vssd1 vssd1 vccd1 vccd1 _08099_/B sky130_fd_sc_hd__xnor2_2
X_07047_ _07047_/A _07056_/B vssd1 vssd1 vccd1 vccd1 _07047_/X sky130_fd_sc_hd__or2_2
XFILLER_0_100_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07177__A3 _07303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11902__B1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__A1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__B2 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09283__B _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ _08962_/X _08977_/Y _08976_/X vssd1 vssd1 vccd1 vccd1 _08998_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08126__A2 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ _07949_/A _07949_/B vssd1 vssd1 vccd1 vccd1 _07982_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11666__C1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout50_A fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ _10960_/A _11174_/A vssd1 vssd1 vccd1 vccd1 _10960_/Y sky130_fd_sc_hd__nand2_1
X_09619_ _09898_/A _09619_/B vssd1 vssd1 vccd1 vccd1 _09621_/B sky130_fd_sc_hd__xnor2_2
X_10891_ _12784_/A fanout52/X _10677_/B _12782_/A vssd1 vssd1 vccd1 vccd1 _10892_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07531__B _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11334__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12630_ _12635_/B _12630_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[13] sky130_fd_sc_hd__and2_4
XFILLER_0_93_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12561_ _12565_/A _12561_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[0] sky130_fd_sc_hd__and2_4
XFILLER_0_25_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12492_ reg1_val[17] curr_PC[17] _12524_/S vssd1 vssd1 vccd1 vccd1 _12493_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_65_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11512_ _11513_/A _11513_/B vssd1 vssd1 vccd1 vccd1 _11618_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_19_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11443_ _11444_/A _11444_/B _11442_/Y vssd1 vssd1 vccd1 vccd1 _11443_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_123_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12933__A2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07259__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13113_ _13113_/A _13113_/B vssd1 vssd1 vccd1 vccd1 _13113_/Y sky130_fd_sc_hd__xnor2_1
X_11374_ _11374_/A _11552_/A vssd1 vssd1 vccd1 vccd1 _11374_/Y sky130_fd_sc_hd__nand2_1
X_10325_ _10325_/A _10325_/B vssd1 vssd1 vccd1 vccd1 _10326_/B sky130_fd_sc_hd__or2_1
XANTENNA__12146__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13044_ hold288/A _13043_/Y hold243/X vssd1 vssd1 vccd1 vccd1 _13044_/X sky130_fd_sc_hd__mux2_1
X_10256_ hold266/A _10256_/B vssd1 vssd1 vccd1 vccd1 _10514_/C sky130_fd_sc_hd__or2_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11509__A _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10413__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ _10187_/A _10187_/B _10187_/C vssd1 vssd1 vccd1 vccd1 _10188_/B sky130_fd_sc_hd__and3_1
XANTENNA__13110__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12828_ hold45/X hold240/X vssd1 vssd1 vccd1 vccd1 _12830_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_84_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12759_ _07168_/Y _12781_/A2 hold59/X _13166_/A vssd1 vssd1 vccd1 vccd1 hold60/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08825__B1 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11424__A2 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13177__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09250__B1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout8 fanout9/A vssd1 vssd1 vccd1 vccd1 fanout8/X sky130_fd_sc_hd__buf_6
XFILLER_0_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09970_ _09970_/A _09970_/B vssd1 vssd1 vccd1 vccd1 _09970_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12137__B1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08921_ _08919_/A _08919_/B _08922_/B vssd1 vssd1 vccd1 vccd1 _08921_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08356__A2 _08692_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08852_ _08348_/B fanout94/X _07197_/Y _07181_/Y vssd1 vssd1 vccd1 vccd1 _08853_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09553__A1 _10249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07803_ _07802_/A _07802_/B _07802_/C vssd1 vssd1 vccd1 vccd1 _07804_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07564__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08783_ _08784_/A _08784_/B vssd1 vssd1 vccd1 vccd1 _08783_/X sky130_fd_sc_hd__and2b_1
XANTENNA_fanout185_A _08415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07734_ _07734_/A _07734_/B vssd1 vssd1 vccd1 vccd1 _07737_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07665_ _08903_/A _08903_/B vssd1 vssd1 vccd1 vccd1 _08904_/A sky130_fd_sc_hd__and2_1
X_06616_ reg1_val[26] _07153_/A vssd1 vssd1 vccd1 vccd1 _06619_/A sky130_fd_sc_hd__nand2_2
X_09404_ _09328_/A _09328_/B _09326_/X vssd1 vssd1 vccd1 vccd1 _09506_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_48_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07596_ _07596_/A _07596_/B vssd1 vssd1 vccd1 vccd1 _07604_/B sky130_fd_sc_hd__or2_2
X_06547_ rst vssd1 vssd1 vccd1 vccd1 _06547_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_118_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09335_ _09224_/X _09559_/C _12223_/B1 vssd1 vssd1 vccd1 vccd1 _09335_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09559__A _09559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09266_ _09267_/A _09267_/B vssd1 vssd1 vccd1 vccd1 _09438_/A sky130_fd_sc_hd__nand2b_1
X_08217_ _08821_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08218_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_62_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09197_ _09197_/A _09197_/B _09197_/C vssd1 vssd1 vccd1 vccd1 _09197_/X sky130_fd_sc_hd__or3_1
XFILLER_0_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08148_ _08158_/B _08158_/A vssd1 vssd1 vccd1 vccd1 _08160_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_70_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ _08133_/A _08133_/B vssd1 vssd1 vccd1 vccd1 _08149_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12713__A _12713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10110_ _10750_/S _09361_/X _11195_/C vssd1 vssd1 vccd1 vccd1 _10110_/X sky130_fd_sc_hd__o21a_1
X_11090_ _10750_/S _10114_/X _11089_/X _10752_/S vssd1 vssd1 vccd1 vccd1 _11090_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout98_A _08348_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09294__A _09294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12679__B2 _07087_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10041_ _09932_/A _09932_/B _09929_/A vssd1 vssd1 vccd1 vccd1 _10052_/A sky130_fd_sc_hd__a21o_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__buf_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07526__B _07526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ hold226/A _11992_/B vssd1 vssd1 vccd1 vccd1 _12059_/B sky130_fd_sc_hd__or2_1
X_10943_ _10943_/A _10943_/B _10941_/Y vssd1 vssd1 vccd1 vccd1 _10944_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_97_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10874_ hold219/A _10874_/B vssd1 vssd1 vccd1 vccd1 _10983_/B sky130_fd_sc_hd__or2_1
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12613_ reg1_val[11] _12614_/B vssd1 vssd1 vccd1 vccd1 _12623_/A sky130_fd_sc_hd__nand2_1
X_12544_ _12551_/A _12545_/B vssd1 vssd1 vccd1 vccd1 _12546_/A sky130_fd_sc_hd__and2_1
XFILLER_0_81_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09469__A _09620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12607__B _12607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11511__B _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12475_ _12632_/B _12475_/B vssd1 vssd1 vccd1 vccd1 _12476_/B sky130_fd_sc_hd__or2_1
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_6 instruction[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11426_ _11427_/A _11427_/B vssd1 vssd1 vccd1 vccd1 _11532_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08586__A2 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09783__B2 _09295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09783__A1 _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ _11355_/X _11357_/B vssd1 vssd1 vccd1 vccd1 _11358_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07794__B1 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10308_ _10308_/A _10308_/B vssd1 vssd1 vccd1 vccd1 _10309_/B sky130_fd_sc_hd__nor2_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11590__B2 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__A1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13027_ hold279/X _13151_/A2 _13026_/X _06537_/A vssd1 vssd1 vccd1 vccd1 _13028_/B
+ sky130_fd_sc_hd__a22o_1
X_11288_ _06816_/Y _11287_/Y _11738_/S vssd1 vssd1 vccd1 vccd1 _11289_/B sky130_fd_sc_hd__mux2_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ _12278_/A _09046_/A _09046_/B _11184_/A _10238_/Y vssd1 vssd1 vccd1 vccd1
+ _10269_/B sky130_fd_sc_hd__a311oi_1
XANTENNA__13095__B2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08548__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08510__A2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07450_ _11125_/A _07450_/B vssd1 vssd1 vccd1 vccd1 _07451_/B sky130_fd_sc_hd__xnor2_4
X_07381_ _07381_/A _07381_/B vssd1 vssd1 vccd1 vccd1 _07385_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09120_ reg1_val[3] reg1_val[28] _09158_/S vssd1 vssd1 vccd1 vccd1 _09120_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09051_ _09050_/A _09050_/B _10370_/C _10370_/B vssd1 vssd1 vccd1 vccd1 _10617_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08002_ _07783_/A _07783_/B _07781_/B _07780_/B _07780_/A vssd1 vssd1 vccd1 vccd1
+ _08008_/A sky130_fd_sc_hd__o32ai_4
XANTENNA__12358__B1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10752__S _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap242 _09192_/Y vssd1 vssd1 vccd1 vccd1 _12228_/B1 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09774__B2 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09774__A1 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout100_A _09925_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11581__A1 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10384__A2 _11838_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09953_ _09954_/A _09954_/B vssd1 vssd1 vccd1 vccd1 _09953_/Y sky130_fd_sc_hd__nand2_1
X_08904_ _08904_/A _08904_/B vssd1 vssd1 vccd1 vccd1 _08910_/A sky130_fd_sc_hd__nor2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11333__A1 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09884_ _10280_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _09887_/A sky130_fd_sc_hd__xnor2_1
X_08835_ _08134_/B _08672_/B _08835_/B1 fanout51/X vssd1 vssd1 vccd1 vccd1 _08836_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_57_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11333__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ _08766_/A _08766_/B _08766_/C vssd1 vssd1 vccd1 vccd1 _08767_/B sky130_fd_sc_hd__nor3_1
XANTENNA__11097__B1 _09200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07717_ _08420_/B fanout84/X fanout81/X _08854_/B2 vssd1 vssd1 vccd1 vccd1 _07718_/B
+ sky130_fd_sc_hd__o22a_1
X_08697_ _07968_/A _07967_/Y _07963_/Y vssd1 vssd1 vccd1 vccd1 _08699_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07648_ _07648_/A _07648_/B vssd1 vssd1 vccd1 vccd1 _08888_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12046__C1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ _07579_/A _07579_/B vssd1 vssd1 vccd1 vccd1 _07580_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08265__A1 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09318_ _07577_/A _07577_/B _07575_/X vssd1 vssd1 vccd1 vccd1 _09320_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_118_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08265__B2 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout13_A fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10590_ _10466_/A _10466_/C _10466_/B vssd1 vssd1 vccd1 vccd1 _10600_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_106_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09249_ _09249_/A _09249_/B vssd1 vssd1 vccd1 vccd1 _09292_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__13010__A1 _06965_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12260_ _12308_/A _12260_/B vssd1 vssd1 vccd1 vccd1 _12263_/A sky130_fd_sc_hd__or2_1
XFILLER_0_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11211_ _11181_/X _11184_/X _11188_/X _11210_/X _06898_/C vssd1 vssd1 vccd1 vccd1
+ _11211_/X sky130_fd_sc_hd__a41o_2
XANTENNA__09765__B2 _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12191_ _06837_/B _12250_/B _10377_/B reg1_val[27] _12382_/S vssd1 vssd1 vccd1 vccd1
+ _12191_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11021__B1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__B1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142_ _11142_/A _11142_/B vssd1 vssd1 vccd1 vccd1 _11143_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10127__A2 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ _11462_/A _11073_/B vssd1 vssd1 vccd1 vccd1 _11215_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__09752__A _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _10553_/B _09752_/B fanout14/X fanout69/X vssd1 vssd1 vccd1 vccd1 _10025_/B
+ sky130_fd_sc_hd__o22a_1
X_11975_ _12072_/A _11975_/B vssd1 vssd1 vccd1 vccd1 _11975_/X sky130_fd_sc_hd__or2_1
XFILLER_0_58_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10926_ _10926_/A _10926_/B vssd1 vssd1 vccd1 vccd1 _10928_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_85_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10857_ _10776_/Y _11215_/A _10856_/Y vssd1 vssd1 vccd1 vccd1 _10857_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ _10789_/A _10789_/B vssd1 vssd1 vccd1 vccd1 _10934_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12527_ _12525_/X _12527_/B vssd1 vssd1 vccd1 vccd1 _12539_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_41_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12458_ _12464_/B _12458_/B vssd1 vssd1 vccd1 vccd1 new_PC[11] sky130_fd_sc_hd__and2_4
XFILLER_0_41_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11409_ _12206_/A _11409_/B vssd1 vssd1 vccd1 vccd1 _11416_/A sky130_fd_sc_hd__xnor2_2
X_12389_ reg1_val[2] curr_PC[2] _12556_/S vssd1 vssd1 vccd1 vccd1 _12391_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06950_ _07303_/B _07175_/A _07001_/C vssd1 vssd1 vccd1 vccd1 _08544_/A sky130_fd_sc_hd__a21o_1
X_06881_ instruction[2] _06881_/B _06881_/C vssd1 vssd1 vccd1 vccd1 _06881_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__06990__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06990__A1 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08620_ _08620_/A _08620_/B _08620_/C vssd1 vssd1 vccd1 vccd1 _08621_/B sky130_fd_sc_hd__nor3_1
XANTENNA_clkbuf_4_10_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07534__A3 _07277_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11866__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08551_ _08559_/A _08555_/B vssd1 vssd1 vccd1 vccd1 _08551_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08482_ _08482_/A _08482_/B vssd1 vssd1 vccd1 vccd1 _08502_/B sky130_fd_sc_hd__xnor2_2
X_07502_ _07502_/A _07502_/B vssd1 vssd1 vccd1 vccd1 _07506_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_77_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07433_ _09467_/A _07433_/B vssd1 vssd1 vccd1 vccd1 _07440_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_43_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13123__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11432__A _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09103_ _09103_/A _09103_/B _09102_/A _09102_/B vssd1 vssd1 vccd1 vccd1 _09103_/X
+ sky130_fd_sc_hd__or4bb_1
X_07364_ _07364_/A _07364_/B vssd1 vssd1 vccd1 vccd1 _07626_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09995__B2 _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07295_ _07295_/A _07295_/B vssd1 vssd1 vccd1 vccd1 _07420_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09034_ _09034_/A _09034_/B vssd1 vssd1 vccd1 vccd1 _09035_/B sky130_fd_sc_hd__and2_1
XFILLER_0_5_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09936_ _09936_/A _09936_/B vssd1 vssd1 vccd1 vccd1 _09938_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09572__A _10301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09867_ _10555_/A _09867_/B vssd1 vssd1 vccd1 vccd1 _09869_/B sky130_fd_sc_hd__xnor2_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08818_ _08818_/A _08818_/B vssd1 vssd1 vccd1 vccd1 _08850_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07092__A _09679_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09798_ _09642_/A _09642_/B _09641_/A vssd1 vssd1 vccd1 vccd1 _09808_/A sky130_fd_sc_hd__a21bo_2
X_08749_ _10306_/A _08749_/B vssd1 vssd1 vccd1 vccd1 _08750_/C sky130_fd_sc_hd__xnor2_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11739_/Y _11740_/X _11747_/X _11759_/X vssd1 vssd1 vccd1 vccd1 _11760_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07820__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10880__A2_N _06928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ _10711_/A _10711_/B vssd1 vssd1 vccd1 vccd1 _10724_/A sky130_fd_sc_hd__and2_1
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _11691_/A _11691_/B vssd1 vssd1 vccd1 vccd1 _11701_/A sky130_fd_sc_hd__nand2_1
X_10642_ _10251_/S _09977_/X _09214_/A vssd1 vssd1 vccd1 vccd1 _10642_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10573_ _10573_/A _10573_/B vssd1 vssd1 vccd1 vccd1 _10589_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_24_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13292_ _13296_/CLK _13292_/D vssd1 vssd1 vccd1 vccd1 hold291/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12312_ _12312_/A _12312_/B vssd1 vssd1 vccd1 vccd1 _12313_/B sky130_fd_sc_hd__or2_1
X_12243_ reg1_val[28] _09202_/B _12243_/B1 _06591_/A vssd1 vssd1 vccd1 vccd1 _12243_/Y
+ sky130_fd_sc_hd__o22ai_1
XFILLER_0_51_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08410__A1 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08410__B2 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12174_ _12174_/A _12174_/B vssd1 vssd1 vccd1 vccd1 _12174_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_102_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11125_ _11125_/A _11125_/B vssd1 vssd1 vccd1 vccd1 _11126_/B sky130_fd_sc_hd__nor2_1
X_11056_ _10945_/A _10945_/B _10942_/X vssd1 vssd1 vccd1 vccd1 _11058_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12620__B _12620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10007_ _08680_/B _07553_/A _10927_/A fanout30/X vssd1 vssd1 vccd1 vccd1 _10008_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08098__A _08853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07921__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07730__A _08853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08826__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11958_ _11958_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _11959_/B sky130_fd_sc_hd__or2_1
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10909_ _10910_/A _10910_/B vssd1 vssd1 vccd1 vccd1 _10909_/Y sky130_fd_sc_hd__nor2_1
X_11889_ _11889_/A vssd1 vssd1 vccd1 vccd1 _11890_/B sky130_fd_sc_hd__inv_2
XFILLER_0_117_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07080_ _10458_/A _10155_/A _07080_/C vssd1 vssd1 vccd1 vccd1 _07080_/X sky130_fd_sc_hd__and3b_1
XFILLER_0_14_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08561__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout107 _07031_/Y vssd1 vssd1 vccd1 vccd1 _10452_/B2 sky130_fd_sc_hd__buf_8
X_07982_ _07982_/A _07982_/B _07982_/C vssd1 vssd1 vccd1 vccd1 _07984_/A sky130_fd_sc_hd__and3_1
Xfanout129 _09742_/A vssd1 vssd1 vccd1 vccd1 _10894_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout118 _07364_/A vssd1 vssd1 vccd1 vccd1 _10306_/A sky130_fd_sc_hd__buf_12
X_06933_ reg1_val[4] reg1_val[5] reg1_val[6] _07105_/B vssd1 vssd1 vccd1 vccd1 _07038_/B
+ sky130_fd_sc_hd__or4_2
X_09721_ _10280_/A _09721_/B vssd1 vssd1 vccd1 vccd1 _09725_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13118__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06864_ _06864_/A _12726_/A vssd1 vssd1 vccd1 vccd1 _06864_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09901__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09901__B2 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10331__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09652_ _09653_/B _09653_/A vssd1 vssd1 vccd1 vccd1 _09652_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06795_ reg1_val[5] _06795_/B vssd1 vssd1 vccd1 vccd1 _06795_/Y sky130_fd_sc_hd__nand2_1
X_08603_ _08576_/X _09041_/A _08577_/X vssd1 vssd1 vccd1 vccd1 _09043_/A sky130_fd_sc_hd__a21oi_2
X_09583_ _09584_/A _09584_/B vssd1 vssd1 vccd1 vccd1 _09736_/A sky130_fd_sc_hd__and2_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08468__A1 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08534_ _09898_/A _08534_/B vssd1 vssd1 vccd1 vccd1 _08541_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08468__B2 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11472__B1 _12228_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08465_ _06864_/A _08841_/A1 _08841_/B2 _08758_/A2 vssd1 vssd1 vccd1 vccd1 _08466_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07140__B2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07140__A1 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08396_ _08390_/A _08390_/B _08390_/C vssd1 vssd1 vccd1 vccd1 _08397_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_80_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07416_ _07414_/A _07414_/B _07415_/Y vssd1 vssd1 vccd1 vccd1 _07624_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12016__A2 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07347_ _07387_/A _07387_/B vssd1 vssd1 vccd1 vccd1 _07388_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09567__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09017_ _09007_/X _09016_/X _08621_/B vssd1 vssd1 vccd1 vccd1 _09060_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07278_ _08588_/A _07278_/B vssd1 vssd1 vccd1 vccd1 _07591_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_33_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06703__B _07192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06651__B1 _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold161 hold161/A vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 hold150/A vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__A2 _11838_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold172 hold172/A vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 hold194/A vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 hold183/A vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07815__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09919_ _09919_/A _09919_/B _09919_/C vssd1 vssd1 vccd1 vccd1 _09921_/A sky130_fd_sc_hd__and3_1
X_12930_ _13147_/A hold179/X vssd1 vssd1 vccd1 vccd1 _13235_/D sky130_fd_sc_hd__and2_1
X_12861_ hold11/X hold294/A vssd1 vssd1 vccd1 vccd1 _13102_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11812_ _11812_/A _11892_/A vssd1 vssd1 vccd1 vccd1 _11969_/A sky130_fd_sc_hd__nand2_1
X_12792_ _12891_/B _12792_/B vssd1 vssd1 vccd1 vccd1 _13162_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08646__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11743_ _11743_/A _11743_/B vssd1 vssd1 vccd1 vccd1 _11745_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11674_ _12345_/A _11670_/X _11673_/X vssd1 vssd1 vccd1 vccd1 dest_val[20] sky130_fd_sc_hd__o21ai_4
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06890__B1 _09199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10625_ _10625_/A _10625_/B vssd1 vssd1 vccd1 vccd1 _10630_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11766__A1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10556_ _10555_/B _10555_/C _10555_/A vssd1 vssd1 vccd1 vccd1 _10562_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_122_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13275_ _13277_/CLK _13275_/D vssd1 vssd1 vccd1 vccd1 hold124/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__06642__B1 _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10487_ _10487_/A _10732_/A vssd1 vssd1 vccd1 vccd1 _10487_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06613__B _06633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12226_ _06612_/B _12169_/X _06610_/Y vssd1 vssd1 vccd1 vccd1 _12226_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07198__A1 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07198__B2 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _12157_/A _12157_/B vssd1 vssd1 vccd1 vccd1 _12160_/C sky130_fd_sc_hd__xnor2_1
X_11108_ curr_PC[13] _11107_/C curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11108_/Y sky130_fd_sc_hd__a21oi_1
X_12088_ _12088_/A _12088_/B vssd1 vssd1 vccd1 vccd1 _12090_/B sky130_fd_sc_hd__xnor2_1
X_11039_ _07195_/B fanout9/X _11038_/X vssd1 vssd1 vccd1 vccd1 _11041_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__09895__B1 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06580_ instruction[39] _06633_/B vssd1 vssd1 vccd1 vccd1 _12632_/B sky130_fd_sc_hd__and2_4
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08250_ _08250_/A _08250_/B vssd1 vssd1 vccd1 vccd1 _08261_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07673__A2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08181_ _08443_/A _08181_/B vssd1 vssd1 vccd1 vccd1 _08245_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07201_ _11431_/A _10527_/A fanout69/X _10452_/B2 vssd1 vssd1 vccd1 vccd1 _07202_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10009__B2 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10009__A1 _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07132_ _12250_/A _07132_/B vssd1 vssd1 vccd1 vccd1 _07132_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07063_ _08532_/B _07055_/Y _07058_/A _12768_/A vssd1 vssd1 vccd1 vccd1 _07064_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07965_ _07074_/Y _07179_/A fanout94/X _08776_/B1 vssd1 vssd1 vccd1 vccd1 _07966_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_4_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06916_ instruction[23] _06552_/X _06915_/X _06678_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[5]
+ sky130_fd_sc_hd__o211a_4
X_09704_ _11400_/A _09702_/Y _09703_/X _11099_/B reg1_val[3] vssd1 vssd1 vccd1 vccd1
+ _09704_/X sky130_fd_sc_hd__o32a_1
X_07896_ _08733_/A _07896_/B vssd1 vssd1 vccd1 vccd1 _08053_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_97_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09635_ _09635_/A _09635_/B vssd1 vssd1 vccd1 vccd1 _09637_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_69_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06847_ _06856_/A _06846_/X _06834_/Y vssd1 vssd1 vccd1 vccd1 _06847_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08466__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06778_ reg2_val[1] _06778_/B vssd1 vssd1 vccd1 vccd1 _06778_/X sky130_fd_sc_hd__and2_1
X_09566_ _08680_/B fanout81/X _09295_/B fanout30/X vssd1 vssd1 vccd1 vccd1 _09567_/B
+ sky130_fd_sc_hd__o22a_1
X_08517_ _08588_/A _07058_/A _08825_/A2 _08532_/B vssd1 vssd1 vccd1 vccd1 _08518_/B
+ sky130_fd_sc_hd__o22a_1
X_09497_ _09321_/A _09321_/B _09319_/Y vssd1 vssd1 vccd1 vccd1 _09498_/B sky130_fd_sc_hd__a21boi_4
XFILLER_0_93_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08310__B1 _07325_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08448_ _09478_/B2 _08532_/B _07058_/A _09476_/A vssd1 vssd1 vccd1 vccd1 _08449_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08379_ _08777_/A _08379_/B vssd1 vssd1 vccd1 vccd1 _08383_/B sky130_fd_sc_hd__xnor2_1
X_10410_ _11125_/A _10410_/B vssd1 vssd1 vccd1 vccd1 _10411_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11390_ _11390_/A _11390_/B vssd1 vssd1 vccd1 vccd1 _11390_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_73_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10341_ _10341_/A _10341_/B vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__xnor2_2
X_13060_ hold268/X _12721_/B _13059_/X _12722_/A vssd1 vssd1 vccd1 vccd1 hold269/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10272_ _12005_/A _10269_/X _10270_/X _10271_/Y vssd1 vssd1 vccd1 vccd1 dest_val[7]
+ sky130_fd_sc_hd__a22o_4
X_12011_ _12011_/A _12011_/B vssd1 vssd1 vccd1 vccd1 _12012_/B sky130_fd_sc_hd__or2_1
X_12913_ hold198/X _12947_/A2 _12947_/B1 hold205/X vssd1 vssd1 vccd1 vccd1 hold206/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09760__A _10578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12844_ _13057_/A _13058_/A _13057_/B vssd1 vssd1 vccd1 vccd1 _13063_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_69_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12775_ hold19/X _12778_/B _12774_/Y _13147_/A vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__o211a_1
XFILLER_0_96_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10239__A1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _11548_/A _11631_/Y _11633_/B vssd1 vssd1 vccd1 vccd1 _11894_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08852__A1 _08348_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08852__B2 _07181_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11657_ _13236_/Q _11751_/C vssd1 vssd1 vccd1 vccd1 _11657_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06624__A _12713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11588_ _11973_/A _11972_/A vssd1 vssd1 vccd1 vccd1 _11588_/Y sky130_fd_sc_hd__nor2_1
X_10608_ _10609_/C _10850_/A vssd1 vssd1 vccd1 vccd1 _10608_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13327_ instruction[8] vssd1 vssd1 vccd1 vccd1 pred_idx[0] sky130_fd_sc_hd__buf_12
XANTENNA__06615__B1 _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10539_ _10539_/A _10539_/B vssd1 vssd1 vccd1 vccd1 _10540_/B sky130_fd_sc_hd__and2_1
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13258_ _13264_/CLK _13258_/D vssd1 vssd1 vccd1 vccd1 hold140/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13189_ _13310_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12209_ _12209_/A _12264_/A _12209_/C vssd1 vssd1 vccd1 vccd1 _12264_/B sky130_fd_sc_hd__nor3_1
X_07750_ _07747_/A _07747_/B _07747_/C vssd1 vssd1 vccd1 vccd1 _07751_/B sky130_fd_sc_hd__a21oi_1
X_06701_ reg1_val[14] _07192_/A vssd1 vssd1 vccd1 vccd1 _06704_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07681_ _07023_/Y _10156_/B2 _10156_/A1 _07034_/Y vssd1 vssd1 vccd1 vccd1 _07682_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11675__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06632_ _06632_/A _06632_/B _12357_/A _06856_/A vssd1 vssd1 vccd1 vccd1 _06632_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_35_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09420_ _09421_/B _09421_/A vssd1 vssd1 vccd1 vccd1 _09645_/B sky130_fd_sc_hd__nand2b_1
X_06563_ instruction[22] _06915_/B vssd1 vssd1 vccd1 vccd1 _06563_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07190__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09351_ _09139_/X _09141_/X _09359_/S vssd1 vssd1 vccd1 vccd1 _09351_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08302_ _08302_/A _08302_/B vssd1 vssd1 vccd1 vccd1 _08334_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11978__A1 _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09282_ _09282_/A _09282_/B vssd1 vssd1 vccd1 vccd1 _09291_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08233_ _08841_/A1 _08772_/B2 _08772_/A2 _08841_/B2 vssd1 vssd1 vccd1 vccd1 _08234_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07646__A2 _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout130_A _09742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08164_ _08633_/A _08633_/B _08163_/Y vssd1 vssd1 vccd1 vccd1 _08643_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_117_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12927__B1 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08095_ _08819_/B2 _08217_/B fanout55/X _12730_/A vssd1 vssd1 vccd1 vccd1 _08096_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07115_ _08589_/A _07115_/B _09898_/A vssd1 vssd1 vccd1 vccd1 _07115_/X sky130_fd_sc_hd__or3b_2
XANTENNA__12255__B _12255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07046_ _09898_/A _07046_/B vssd1 vssd1 vccd1 vccd1 _07056_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_100_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11902__A1 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09571__A2 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _08995_/A _08995_/B _08990_/A vssd1 vssd1 vccd1 vccd1 _09509_/C sky130_fd_sc_hd__a21boi_1
X_07948_ _07948_/A _07948_/B vssd1 vssd1 vccd1 vccd1 _07949_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09580__A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07879_ _07974_/A _07877_/B _07936_/A vssd1 vssd1 vccd1 vccd1 _07888_/A sky130_fd_sc_hd__o21ai_4
X_09618_ _09618_/A1 fanout18/X fanout9/X _09618_/B2 vssd1 vssd1 vccd1 vccd1 _09619_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout43_A _11147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ _11000_/A _11316_/A _11215_/A _12278_/A vssd1 vssd1 vccd1 vccd1 _10890_/X
+ sky130_fd_sc_hd__o31a_1
X_09549_ hold250/A _09549_/B vssd1 vssd1 vccd1 vccd1 _09549_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12560_ reg1_val[0] _12560_/B vssd1 vssd1 vccd1 vccd1 _12561_/B sky130_fd_sc_hd__or2_1
X_12491_ _12500_/A _12491_/B vssd1 vssd1 vccd1 vccd1 new_PC[16] sky130_fd_sc_hd__and2_4
XANTENNA__12446__A _12607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11511_ _11511_/A _12200_/A vssd1 vssd1 vccd1 vccd1 _11513_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11442_ _11340_/A _11340_/B _11337_/A vssd1 vssd1 vccd1 vccd1 _11442_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_18_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07259__B _07259_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08598__A0 _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11373_ _11175_/Y _11552_/A _11371_/X vssd1 vssd1 vccd1 vccd1 _11373_/Y sky130_fd_sc_hd__a21oi_1
X_13112_ _13112_/A _13112_/B vssd1 vssd1 vccd1 vccd1 _13113_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_104_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10324_ _10325_/A _10325_/B vssd1 vssd1 vccd1 vccd1 _10326_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12146__A1 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13043_ _13043_/A _13043_/B vssd1 vssd1 vccd1 vccd1 _13043_/Y sky130_fd_sc_hd__xnor2_1
X_10255_ _06986_/A _06928_/X _10377_/B reg1_val[7] vssd1 vssd1 vccd1 vccd1 _10255_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12181__A _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09474__B _09474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12146__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ _10187_/A _10187_/B _10187_/C vssd1 vssd1 vccd1 vccd1 _10346_/A sky130_fd_sc_hd__a21oi_1
Xfanout290 _13116_/A vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_4_15_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12827_ hold279/A hold29/X vssd1 vssd1 vccd1 vccd1 _13029_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12758_ hold58/X _12786_/B vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__or2_1
XANTENNA__08825__B2 _07000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08825__A1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12689_ _12708_/B _07086_/C _12698_/B vssd1 vssd1 vccd1 vccd1 _12690_/B sky130_fd_sc_hd__a21bo_2
XFILLER_0_16_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11709_ _11709_/A _11709_/B vssd1 vssd1 vccd1 vccd1 _11710_/B sky130_fd_sc_hd__and2_1
XFILLER_0_126_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout9 fanout9/A vssd1 vssd1 vccd1 vccd1 fanout9/X sky130_fd_sc_hd__buf_6
XANTENNA__09250__A1 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09250__B2 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09384__B _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08920_ _08830_/Y _08848_/B _08846_/X vssd1 vssd1 vccd1 vccd1 _08922_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08851_ _08731_/A _08731_/B _08727_/Y vssd1 vssd1 vccd1 vccd1 _08862_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__09553__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _07802_/A _07802_/B _07802_/C vssd1 vssd1 vccd1 vccd1 _07804_/A sky130_fd_sc_hd__and3_1
XANTENNA__07564__A1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07564__B2 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08782_ _08782_/A _08782_/B vssd1 vssd1 vccd1 vccd1 _08784_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07733_ _07734_/A _07734_/B vssd1 vssd1 vccd1 vccd1 _07733_/X sky130_fd_sc_hd__or2_1
XANTENNA__11648__B1 _12228_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07664_ _10306_/A _07664_/B vssd1 vssd1 vccd1 vccd1 _08903_/B sky130_fd_sc_hd__xnor2_1
X_06615_ _06614_/Y _06688_/B1 _06752_/A reg2_val[26] vssd1 vssd1 vccd1 vccd1 _07153_/A
+ sky130_fd_sc_hd__a2bb2o_4
X_09403_ _09559_/A wire3/X _09559_/C _10617_/A vssd1 vssd1 vccd1 vccd1 _09403_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_48_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07595_ _07595_/A _07595_/B _07595_/C vssd1 vssd1 vccd1 vccd1 _07596_/B sky130_fd_sc_hd__nor3_1
XANTENNA__08744__A _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09334_ _09660_/C _09334_/B vssd1 vssd1 vccd1 vccd1 _09559_/C sky130_fd_sc_hd__xnor2_2
X_06546_ _11823_/S vssd1 vssd1 vccd1 vccd1 _11647_/S sky130_fd_sc_hd__inv_2
XFILLER_0_117_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09265_ _10180_/A _09265_/B vssd1 vssd1 vccd1 vccd1 _09267_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08216_ _08853_/A _08216_/B vssd1 vssd1 vccd1 vccd1 _08283_/A sky130_fd_sc_hd__xnor2_1
X_09196_ _12228_/B1 _11838_/A2 _08594_/B vssd1 vssd1 vccd1 vccd1 _09197_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08147_ _08169_/A _08169_/B _08136_/X vssd1 vssd1 vccd1 vccd1 _08158_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08078_ _08443_/A _08078_/B vssd1 vssd1 vccd1 vccd1 _08133_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12128__A1 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07029_ _08777_/A _07030_/B vssd1 vssd1 vccd1 vccd1 _07031_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12128__B2 _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10139__B1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09294__B _10694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10040_ _10040_/A _10040_/B vssd1 vssd1 vccd1 vccd1 _10073_/A sky130_fd_sc_hd__xor2_2
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10541__A2_N fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ hold262/A _12119_/B1 _12056_/B _11990_/Y _11400_/A vssd1 vssd1 vccd1 vccd1
+ _11991_/X sky130_fd_sc_hd__a311o_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13036__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12300__B2 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10942_ _10943_/A _10943_/B _10941_/Y vssd1 vssd1 vccd1 vccd1 _10942_/X sky130_fd_sc_hd__o21ba_1
X_10873_ _11831_/S _10867_/Y _10872_/X vssd1 vssd1 vccd1 vccd1 _10873_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_109_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12612_ _12617_/B _12612_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[10] sky130_fd_sc_hd__and2_4
XFILLER_0_108_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12543_ reg1_val[25] curr_PC[25] _12556_/S vssd1 vssd1 vccd1 vccd1 _12545_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10614__A1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12474_ _12632_/B _12475_/B vssd1 vssd1 vccd1 vccd1 _12485_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_7 instruction[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10378__B1 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11425_ _11853_/A _11425_/B vssd1 vssd1 vccd1 vccd1 _11427_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09783__A2 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11356_ _11356_/A _11356_/B _11356_/C vssd1 vssd1 vccd1 vccd1 _11357_/B sky130_fd_sc_hd__or3_1
XFILLER_0_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07794__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07794__A1 _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10307_ _10308_/A _10308_/B vssd1 vssd1 vccd1 vccd1 _10461_/B sky130_fd_sc_hd__and2_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11590__A2 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06621__B _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13026_ hold240/X _13025_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _13026_/X sky130_fd_sc_hd__mux2_1
X_11287_ _11187_/A _11185_/Y _06698_/B vssd1 vssd1 vccd1 vccd1 _11287_/Y sky130_fd_sc_hd__o21ai_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08743__B1 _08681_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10238_ _12278_/A _09046_/A _09046_/B vssd1 vssd1 vccd1 vccd1 _10238_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10169_ _10169_/A _10169_/B vssd1 vssd1 vccd1 vccd1 _10170_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13095__A2 _13151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11645__A3 _09073_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07380_ _07380_/A _07380_/B vssd1 vssd1 vccd1 vccd1 _07381_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_32_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09471__A1 _08311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09050_ _09050_/A _09050_/B vssd1 vssd1 vccd1 vccd1 _09050_/X sky130_fd_sc_hd__or2_1
XFILLER_0_4_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08001_ _07841_/A _07839_/Y _07838_/X vssd1 vssd1 vccd1 vccd1 _08009_/A sky130_fd_sc_hd__a21boi_4
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10369__B1 _10370_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09774__A2 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09952_ _09952_/A _09952_/B vssd1 vssd1 vccd1 vccd1 _09954_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_12_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08903_ _08903_/A _08903_/B vssd1 vssd1 vccd1 vccd1 _08904_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout295_A _13028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08734__B1 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11869__B1 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09883_ _10144_/B2 fanout26/X _10433_/A _07098_/Y vssd1 vssd1 vccd1 vccd1 _09884_/B
+ sky130_fd_sc_hd__o22a_1
X_08834_ _08834_/A _08834_/B vssd1 vssd1 vccd1 vccd1 _08847_/A sky130_fd_sc_hd__xor2_2
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10541__B1 _11222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08765_ _08766_/A _08766_/B _08766_/C vssd1 vssd1 vccd1 vccd1 _08870_/B sky130_fd_sc_hd__o21a_1
XANTENNA__07643__A _08232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07716_ _07716_/A _07716_/B _07716_/C vssd1 vssd1 vccd1 vccd1 _07727_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06760__A2 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08696_ _08696_/A _08696_/B vssd1 vssd1 vccd1 vccd1 _08699_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_67_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07647_ _08853_/A _07647_/B vssd1 vssd1 vccd1 vccd1 _08888_/A sky130_fd_sc_hd__xor2_1
X_07578_ _07579_/A _07579_/B vssd1 vssd1 vccd1 vccd1 _07578_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09317_ _07542_/A _07542_/B _07540_/X vssd1 vssd1 vccd1 vccd1 _09320_/A sky130_fd_sc_hd__a21o_2
XANTENNA__08265__A2 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09248_ _09249_/A _09249_/B vssd1 vssd1 vccd1 vccd1 _09418_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07473__B1 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13010__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09179_ _09180_/A curr_PC[0] vssd1 vssd1 vccd1 vccd1 _09374_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11210_ _09205_/B _11197_/X _11207_/X _11209_/X vssd1 vssd1 vccd1 vccd1 _11210_/X
+ sky130_fd_sc_hd__o211a_1
X_12190_ _06612_/B _09194_/Y _10638_/B vssd1 vssd1 vccd1 vccd1 _12190_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09765__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11021__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11021__A1 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07776__B2 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__A1 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11141_ _11142_/A _11142_/B vssd1 vssd1 vccd1 vccd1 _11262_/D sky130_fd_sc_hd__and2b_1
XANTENNA__10780__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11072_ _10613_/B _10850_/B _11279_/A _11071_/X vssd1 vssd1 vccd1 vccd1 _11073_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08725__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__B _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ _10180_/A _10023_/B vssd1 vssd1 vccd1 vccd1 _10027_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07553__A _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ _12072_/A _11975_/B vssd1 vssd1 vccd1 vccd1 _11974_/Y sky130_fd_sc_hd__nand2_1
X_10925_ _10925_/A _10925_/B _10925_/C vssd1 vssd1 vccd1 vccd1 _10926_/B sky130_fd_sc_hd__or3_1
X_10856_ _10776_/Y _11215_/A _09110_/X vssd1 vssd1 vccd1 vccd1 _10856_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09199__B _09199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06616__B _07153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10787_ _11604_/A _10787_/B vssd1 vssd1 vccd1 vccd1 _10789_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12526_ _12551_/A _12526_/B vssd1 vssd1 vccd1 vccd1 _12527_/B sky130_fd_sc_hd__or2_1
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12457_ _12457_/A _12457_/B _12457_/C vssd1 vssd1 vccd1 vccd1 _12458_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11408_ _11794_/A fanout27/X _12205_/A _11704_/A vssd1 vssd1 vccd1 vccd1 _11409_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_111_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12388_ _12394_/B _12388_/B vssd1 vssd1 vccd1 vccd1 new_PC[1] sky130_fd_sc_hd__and2_4
XFILLER_0_1_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11339_ _12019_/A _11339_/B vssd1 vssd1 vccd1 vccd1 _11340_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_120_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06880_ instruction[2] _06881_/B _06881_/C vssd1 vssd1 vccd1 vccd1 _06898_/C sky130_fd_sc_hd__and3_4
XFILLER_0_94_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13009_ hold118/X _13013_/A2 _13020_/A2 hold124/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold125/A sky130_fd_sc_hd__o221a_1
XANTENNA__06990__A2 _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07534__A4 _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08550_ _08550_/A _08550_/B vssd1 vssd1 vccd1 vccd1 _08555_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_77_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08481_ _08489_/A _08489_/B _08474_/Y vssd1 vssd1 vccd1 vccd1 _08502_/A sky130_fd_sc_hd__a21bo_1
X_07501_ _07502_/A _07502_/B vssd1 vssd1 vccd1 vccd1 _07501_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_119_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07432_ _09618_/B2 fanout22/X _10677_/A _09618_/A1 vssd1 vssd1 vccd1 vccd1 _07433_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_92_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09102_ _09102_/A _09102_/B vssd1 vssd1 vccd1 vccd1 _09102_/Y sky130_fd_sc_hd__nand2_1
X_07363_ _09772_/A _08680_/B fanout30/X _09478_/B2 vssd1 vssd1 vccd1 vccd1 _07364_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10329__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07294_ _07601_/B _07294_/B vssd1 vssd1 vccd1 vccd1 _07420_/A sky130_fd_sc_hd__or2_1
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07455__B1 _10553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09033_ _08595_/A _09514_/A _08595_/B vssd1 vssd1 vccd1 vccd1 _09034_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12751__A1 _10811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09935_ _09935_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09936_/B sky130_fd_sc_hd__xor2_2
X_09866_ _08681_/A fanout57/X fanout94/X _09295_/A vssd1 vssd1 vccd1 vccd1 _09867_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _08818_/A _08818_/B vssd1 vssd1 vccd1 vccd1 _08919_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08469__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09797_ _09797_/A _09797_/B vssd1 vssd1 vccd1 vccd1 _09810_/A sky130_fd_sc_hd__xor2_4
X_08748_ _08821_/A fanout30/X _08748_/B1 _08680_/B vssd1 vssd1 vccd1 vccd1 _08749_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08679_ _08678_/B _08678_/C _08678_/A vssd1 vssd1 vccd1 vccd1 _08679_/X sky130_fd_sc_hd__a21o_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10710_ _10710_/A _10710_/B vssd1 vssd1 vccd1 vccd1 _10711_/B sky130_fd_sc_hd__nand2_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11690_ _11690_/A _11690_/B vssd1 vssd1 vccd1 vccd1 _11691_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_119_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ _10641_/A _10641_/B _10641_/C vssd1 vssd1 vccd1 vccd1 _10641_/X sky130_fd_sc_hd__and3_1
XFILLER_0_63_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08932__A _08932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10572_ _10573_/A _10573_/B vssd1 vssd1 vccd1 vccd1 _10572_/Y sky130_fd_sc_hd__nand2b_1
X_13291_ _13296_/CLK _13291_/D vssd1 vssd1 vccd1 vccd1 hold301/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12990__A1 _07259_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12311_ _12311_/A _12311_/B vssd1 vssd1 vccd1 vccd1 _12316_/A sky130_fd_sc_hd__nand2_1
X_12242_ hold270/A _11398_/B _12285_/B _11400_/A vssd1 vssd1 vccd1 vccd1 _12242_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12454__A _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08410__A2 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ _12131_/B _12133_/A _12131_/A vssd1 vssd1 vccd1 vccd1 _12174_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09763__A _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11124_ _11125_/A _11125_/B vssd1 vssd1 vccd1 vccd1 _11126_/A sky130_fd_sc_hd__and2_1
X_11055_ _11055_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11058_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08379__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10006_ _10006_/A _10006_/B vssd1 vssd1 vccd1 vccd1 _10020_/A sky130_fd_sc_hd__nor2_2
XANTENNA__07921__A1 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07921__B2 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11957_ _11958_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _12036_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10808__A1 _10453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10908_ _10908_/A _10908_/B vssd1 vssd1 vccd1 vccd1 _10910_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_67_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09003__A _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11888_ _11888_/A _11888_/B _11888_/C vssd1 vssd1 vccd1 vccd1 _11889_/A sky130_fd_sc_hd__and3_1
XANTENNA__10149__A _10149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10839_ _10839_/A _10839_/B vssd1 vssd1 vccd1 vccd1 _10842_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08842__A _08842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07437__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12509_ _12516_/A _12509_/B vssd1 vssd1 vccd1 vccd1 _12510_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_89_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12733__A1 _09600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10744__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07981_ _07980_/B _07980_/C _07980_/A vssd1 vssd1 vccd1 vccd1 _07982_/C sky130_fd_sc_hd__o21ai_1
Xfanout108 _12762_/A vssd1 vssd1 vccd1 vccd1 _11431_/A sky130_fd_sc_hd__buf_6
XFILLER_0_1_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06932_ _09180_/A _12563_/A reg1_val[2] reg1_val[3] vssd1 vssd1 vccd1 vccd1 _07105_/B
+ sky130_fd_sc_hd__or4_2
X_09720_ _10144_/B2 _07389_/B fanout26/X _10064_/B2 vssd1 vssd1 vccd1 vccd1 _09721_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07193__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06863_ _09180_/A _09362_/S vssd1 vssd1 vccd1 vccd1 _08594_/B sky130_fd_sc_hd__nand2_2
XANTENNA__09901__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09651_ _09651_/A _09651_/B vssd1 vssd1 vccd1 vccd1 _09653_/B sky130_fd_sc_hd__xnor2_2
X_06794_ _06868_/C _06792_/Y _06793_/X vssd1 vssd1 vccd1 vccd1 _06794_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08602_ _08602_/A _08602_/B vssd1 vssd1 vccd1 vccd1 _09041_/B sky130_fd_sc_hd__xnor2_1
X_09582_ _10555_/A _09582_/B vssd1 vssd1 vccd1 vccd1 _09584_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08533_ _08825_/A2 _09618_/A1 _09476_/A _09618_/B2 vssd1 vssd1 vccd1 vccd1 _08534_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout160_A _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _12345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08468__A2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06537__A _06537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08464_ _09467_/A _08464_/B vssd1 vssd1 vccd1 vccd1 _08471_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07140__A2 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08395_ _08421_/A _08421_/B vssd1 vssd1 vccd1 vccd1 _08432_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_64_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07415_ _07696_/B _07696_/A vssd1 vssd1 vccd1 vccd1 _07415_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_58_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07346_ _09580_/A _07346_/B vssd1 vssd1 vccd1 vccd1 _07387_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12972__A1 _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09016_ _09009_/X _09014_/Y _08457_/X _09057_/A vssd1 vssd1 vccd1 vccd1 _09016_/X
+ sky130_fd_sc_hd__a211o_1
X_07277_ _12255_/A _07277_/B vssd1 vssd1 vccd1 vccd1 _07277_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__12185__C1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold140 hold140/A vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 hold162/A vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 hold184/A vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12721__B _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09918_ _10006_/B _09917_/C _09917_/A vssd1 vssd1 vccd1 vccd1 _09919_/C sky130_fd_sc_hd__o21ai_2
XANTENNA_fanout73_A _07069_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10499__C1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09849_ _09847_/Y _09849_/B vssd1 vssd1 vccd1 vccd1 _09850_/B sky130_fd_sc_hd__nand2b_1
X_12860_ _13097_/A _13098_/A _13097_/B vssd1 vssd1 vccd1 vccd1 _13103_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__11209__A1_N _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11633_/A _11721_/A _11723_/B vssd1 vssd1 vccd1 vccd1 _11811_/X sky130_fd_sc_hd__a21o_1
X_12791_ _13163_/A hold3/X vssd1 vssd1 vccd1 vccd1 _12792_/B sky130_fd_sc_hd__nand2_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11742_ reg1_val[21] curr_PC[21] vssd1 vssd1 vccd1 vccd1 _11743_/B sky130_fd_sc_hd__or2_1
XFILLER_0_56_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11673_ _12556_/S _11764_/B _11673_/C vssd1 vssd1 vccd1 vccd1 _11673_/X sky130_fd_sc_hd__or3_2
XFILLER_0_49_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06890__A1 _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10624_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10625_/B sky130_fd_sc_hd__or2_1
XFILLER_0_64_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08662__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10555_ _10555_/A _10555_/B _10555_/C vssd1 vssd1 vccd1 vccd1 _10562_/A sky130_fd_sc_hd__and3_1
X_13274_ _13277_/CLK hold120/X vssd1 vssd1 vccd1 vccd1 hold118/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07278__A _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10486_ _10486_/A _10607_/A vssd1 vssd1 vccd1 vccd1 _10732_/A sky130_fd_sc_hd__nor2_1
X_12225_ _12322_/S _12225_/B vssd1 vssd1 vccd1 vccd1 _12225_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12191__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07198__A2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12156_ _12157_/A _12157_/B vssd1 vssd1 vccd1 vccd1 _12213_/B sky130_fd_sc_hd__and2_1
X_11107_ curr_PC[13] curr_PC[14] _11107_/C vssd1 vssd1 vccd1 vccd1 _11213_/B sky130_fd_sc_hd__and3_1
XANTENNA__12631__B _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12087_ _12087_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _12088_/B sky130_fd_sc_hd__nor2_1
X_11038_ _08733_/A _07194_/C _07435_/Y _08857_/A vssd1 vssd1 vccd1 vccd1 _11038_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09895__A1 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09895__B2 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12989_ hold42/X _13013_/A2 _13020_/A2 _13265_/Q _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold43/A sky130_fd_sc_hd__o221a_1
XFILLER_0_87_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07658__B1 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12078__B _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08180_ _08692_/A2 _12752_/A fanout84/X _08692_/B1 vssd1 vssd1 vccd1 vccd1 _08181_/B
+ sky130_fd_sc_hd__o22a_1
X_07200_ _07631_/A _07631_/B vssd1 vssd1 vccd1 vccd1 _07632_/A sky130_fd_sc_hd__or2_2
XFILLER_0_55_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10009__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07131_ _06837_/B _07128_/X _07135_/B vssd1 vssd1 vccd1 vccd1 _07132_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08572__A _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07062_ _07062_/A _07062_/B vssd1 vssd1 vccd1 vccd1 _07062_/X sky130_fd_sc_hd__and2_1
XFILLER_0_30_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11914__C1 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07964_ _07964_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _07968_/A sky130_fd_sc_hd__xor2_2
X_06915_ instruction[30] _06915_/B vssd1 vssd1 vccd1 vccd1 _06915_/X sky130_fd_sc_hd__or2_1
X_09703_ hold246/A _09842_/B _09841_/B vssd1 vssd1 vccd1 vccd1 _09703_/X sky130_fd_sc_hd__and3_1
X_07895_ _10149_/A _07173_/Y _07182_/X _10035_/A vssd1 vssd1 vccd1 vccd1 _07896_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09335__B1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06846_ _12276_/A _06845_/Y _06835_/Y vssd1 vssd1 vccd1 vccd1 _06846_/X sky130_fd_sc_hd__o21a_1
X_09634_ _09634_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09635_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07005__A_N _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06777_ _09694_/A _06777_/B vssd1 vssd1 vccd1 vccd1 _06870_/A sky130_fd_sc_hd__nand2b_2
X_09565_ _10280_/A _09565_/B vssd1 vssd1 vccd1 vccd1 _09569_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08516_ _08540_/A _08540_/B _08516_/C vssd1 vssd1 vccd1 vccd1 _08521_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_38_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09496_ _09496_/A _09496_/B vssd1 vssd1 vccd1 vccd1 _09498_/A sky130_fd_sc_hd__xnor2_4
X_08447_ _08453_/A _08453_/B vssd1 vssd1 vccd1 vccd1 _08447_/X sky130_fd_sc_hd__and2_1
XFILLER_0_46_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08378_ _08819_/B2 _08477_/B _08776_/B1 _12730_/A vssd1 vssd1 vccd1 vccd1 _08379_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_92_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06714__B _07303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07329_ _07329_/A _07329_/B vssd1 vssd1 vccd1 vccd1 _07330_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_6_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10340_ _10340_/A _10340_/B vssd1 vssd1 vccd1 vccd1 _10341_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10271_ curr_PC[7] _10397_/C _12005_/A vssd1 vssd1 vccd1 vccd1 _10271_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12173__A2 _12133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ _12011_/A _12011_/B vssd1 vssd1 vccd1 vccd1 _12012_/A sky130_fd_sc_hd__nand2_1
X_12912_ _12946_/A hold199/X vssd1 vssd1 vccd1 vccd1 _13226_/D sky130_fd_sc_hd__and2_1
X_12843_ hold73/X hold292/A vssd1 vssd1 vccd1 vccd1 _13057_/B sky130_fd_sc_hd__nand2b_1
X_12774_ _12774_/A _12778_/B vssd1 vssd1 vccd1 vccd1 _12774_/Y sky130_fd_sc_hd__nand2_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11725_ _11893_/A vssd1 vssd1 vccd1 vccd1 _11725_/Y sky130_fd_sc_hd__inv_2
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08852__A2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11656_ _11746_/A _10765_/Y _11655_/Y _06918_/X vssd1 vssd1 vccd1 vccd1 _11668_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__08392__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout90 _07255_/Y vssd1 vssd1 vccd1 vccd1 _08836_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__12626__B _12626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06624__B _12370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11587_ _11730_/A _11730_/B _11730_/C vssd1 vssd1 vccd1 vccd1 _11972_/A sky130_fd_sc_hd__nor3_1
XANTENNA__10427__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10607_ _10607_/A _10730_/A vssd1 vssd1 vccd1 vccd1 _10850_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13326_ instruction[6] vssd1 vssd1 vccd1 vccd1 loadstore_size[1] sky130_fd_sc_hd__buf_12
X_10538_ _10539_/A _10539_/B vssd1 vssd1 vccd1 vccd1 _10662_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_3_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13257_ _13264_/CLK hold136/X vssd1 vssd1 vccd1 vccd1 hold134/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07736__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12208_ _12208_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12209_/C sky130_fd_sc_hd__and2_1
X_10469_ _10342_/A _10342_/B _10326_/A vssd1 vssd1 vccd1 vccd1 _10479_/A sky130_fd_sc_hd__o21ai_4
X_13188_ _13280_/CLK _13188_/D vssd1 vssd1 vccd1 vccd1 hold105/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12361__B _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12139_ curr_PC[27] _12139_/B vssd1 vssd1 vccd1 vccd1 _12139_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06700_ _06898_/A _06641_/A _12637_/B _06699_/X vssd1 vssd1 vccd1 vccd1 _07192_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__11675__A1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07680_ _08415_/A _07680_/B vssd1 vssd1 vccd1 vccd1 _08812_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11675__B2 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06631_ _06631_/A _06631_/B vssd1 vssd1 vccd1 vccd1 _06856_/A sky130_fd_sc_hd__nor2_2
X_06562_ instruction[12] _06552_/X _06561_/X _06678_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[1]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_75_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09350_ _09348_/X _09349_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09350_/X sky130_fd_sc_hd__mux2_1
X_08301_ _08301_/A _08301_/B vssd1 vssd1 vccd1 vccd1 _08341_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_75_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09281_ _09281_/A _09281_/B vssd1 vssd1 vccd1 vccd1 _09282_/B sky130_fd_sc_hd__xnor2_2
X_08232_ _08232_/A _08232_/B vssd1 vssd1 vccd1 vccd1 _08235_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_90_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08163_ _08635_/B _08635_/A vssd1 vssd1 vccd1 vccd1 _08163_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout123_A _07324_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08094_ _08855_/A _08094_/B vssd1 vssd1 vccd1 vccd1 _08099_/A sky130_fd_sc_hd__xnor2_2
X_07114_ _07126_/B _07114_/B vssd1 vssd1 vccd1 vccd1 _12774_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07045_ _09898_/A _07046_/B vssd1 vssd1 vccd1 vccd1 _07045_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08996_ _09090_/A _09090_/B _08979_/Y _09507_/B _09660_/B vssd1 vssd1 vccd1 vccd1
+ _09000_/A sky130_fd_sc_hd__a2111o_1
X_07947_ _07948_/A _07948_/B vssd1 vssd1 vccd1 vccd1 _07947_/X sky130_fd_sc_hd__and2b_1
X_07878_ _07935_/A _07935_/B _07935_/C vssd1 vssd1 vccd1 vccd1 _07936_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_97_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08477__A _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06829_ _11824_/A _06829_/B vssd1 vssd1 vccd1 vccd1 _06829_/X sky130_fd_sc_hd__or2_1
X_09617_ _09736_/D _09617_/B vssd1 vssd1 vccd1 vccd1 _09635_/A sky130_fd_sc_hd__nor2_1
X_09548_ hold279/A hold240/A _09385_/C vssd1 vssd1 vccd1 vccd1 _09549_/B sky130_fd_sc_hd__o21a_1
XANTENNA__06709__B _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11510_ _11618_/C _11510_/B vssd1 vssd1 vccd1 vccd1 _11513_/A sky130_fd_sc_hd__or2_1
XFILLER_0_19_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09479_ _09775_/A _09479_/B vssd1 vssd1 vccd1 vccd1 _09481_/B sky130_fd_sc_hd__xnor2_2
X_12490_ _12490_/A _12490_/B _12490_/C vssd1 vssd1 vccd1 vccd1 _12491_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_93_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08047__B1 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11441_ _11350_/A _11350_/B _11349_/A vssd1 vssd1 vccd1 vccd1 _11446_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_116_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11372_ _11462_/B _11460_/A vssd1 vssd1 vccd1 vccd1 _11552_/A sky130_fd_sc_hd__nor2_1
X_13111_ _13116_/A hold290/X vssd1 vssd1 vccd1 vccd1 _13299_/D sky130_fd_sc_hd__and2_1
XFILLER_0_61_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10323_ _10323_/A _10323_/B vssd1 vssd1 vccd1 vccd1 _10325_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12146__A2 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13042_ _13086_/A _13042_/B vssd1 vssd1 vccd1 vccd1 _13285_/D sky130_fd_sc_hd__and2_1
X_10254_ _13224_/Q _12124_/B _10509_/C _12290_/C1 vssd1 vssd1 vccd1 vccd1 _10254_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10185_ _10185_/A _10185_/B vssd1 vssd1 vccd1 vccd1 _10187_/C sky130_fd_sc_hd__xnor2_1
Xfanout291 _06547_/Y vssd1 vssd1 vccd1 vccd1 _13116_/A sky130_fd_sc_hd__buf_2
XANTENNA__11106__B1 _06898_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout280 _06569_/X vssd1 vssd1 vccd1 vccd1 _06778_/B sky130_fd_sc_hd__clkbuf_4
X_12826_ hold250/X hold105/X vssd1 vssd1 vccd1 vccd1 _13034_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12757_ _11147_/A _12781_/A2 hold66/X _13166_/A vssd1 vssd1 vccd1 vccd1 hold67/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08825__A2 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12688_ _12688_/A _12688_/B vssd1 vssd1 vccd1 vccd1 _12698_/B sky130_fd_sc_hd__or2_1
XFILLER_0_37_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11708_ _11709_/A _11709_/B vssd1 vssd1 vccd1 vccd1 _11797_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_126_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08038__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10157__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11639_ _11459_/Y _11814_/A _11638_/Y _11634_/Y vssd1 vssd1 vccd1 vccd1 _11639_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13309_ _13309_/CLK _13309_/D vssd1 vssd1 vccd1 vccd1 hold270/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09250__A2 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10396__A1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11345__B1 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08850_ _08850_/A _08850_/B vssd1 vssd1 vccd1 vccd1 _08866_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_20_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07801_ _07801_/A _07801_/B vssd1 vssd1 vccd1 vccd1 _07802_/C sky130_fd_sc_hd__xor2_1
XANTENNA__07564__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08781_ _08667_/A _08667_/B _08663_/X vssd1 vssd1 vccd1 vccd1 _08782_/B sky130_fd_sc_hd__a21o_1
X_07732_ _10578_/A _07732_/B vssd1 vssd1 vccd1 vccd1 _07734_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07663_ _09478_/B2 _08680_/B fanout30/X _09476_/A vssd1 vssd1 vccd1 vccd1 _07664_/B
+ sky130_fd_sc_hd__o22a_1
X_06614_ _06687_/A _12614_/B vssd1 vssd1 vccd1 vccd1 _06614_/Y sky130_fd_sc_hd__nor2_1
X_09402_ _09712_/B _09402_/B vssd1 vssd1 vccd1 vccd1 _09402_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09333_ _09660_/A _09660_/B _10230_/A _09332_/X vssd1 vssd1 vccd1 vccd1 _09334_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07594_ _07595_/A _07595_/B _07595_/C vssd1 vssd1 vccd1 vccd1 _07596_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06545_ reg1_val[31] vssd1 vssd1 vccd1 vccd1 _12713_/A sky130_fd_sc_hd__inv_6
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09264_ _11347_/A fanout52/X _10677_/B _11134_/B2 vssd1 vssd1 vccd1 vccd1 _09265_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08215_ _08748_/B1 _07181_/Y _12730_/A fanout98/X vssd1 vssd1 vccd1 vccd1 _08216_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09195_ _09200_/A _09200_/B _09201_/B vssd1 vssd1 vccd1 vccd1 _09383_/B sky130_fd_sc_hd__or3_4
XFILLER_0_7_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10067__A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08146_ _08146_/A _08146_/B vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_16_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10387__A1 _09198_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11584__B1 _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08077_ _08692_/A2 fanout94/X _12752_/A _08692_/B1 vssd1 vssd1 vccd1 vccd1 _08078_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07028_ reg1_val[10] _07028_/B vssd1 vssd1 vccd1 vccd1 _07030_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
X_08979_ _09103_/B _09102_/A vssd1 vssd1 vccd1 vccd1 _08979_/Y sky130_fd_sc_hd__nand2b_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _12119_/B1 _12056_/B hold262/A vssd1 vssd1 vccd1 vccd1 _11990_/Y sky130_fd_sc_hd__a21oi_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ _10813_/A _10813_/B _10811_/X vssd1 vssd1 vccd1 vccd1 _10941_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10872_ _11197_/S _10872_/B _10871_/X vssd1 vssd1 vccd1 vccd1 _10872_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09530__S _09679_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ _12611_/A _12611_/B _12611_/C vssd1 vssd1 vccd1 vccd1 _12612_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12542_ _12542_/A _12542_/B vssd1 vssd1 vccd1 vccd1 new_PC[24] sky130_fd_sc_hd__xor2_4
XFILLER_0_38_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12473_ reg1_val[14] curr_PC[14] _12524_/S vssd1 vssd1 vccd1 vccd1 _12475_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11424_ _10553_/A _12203_/A _12150_/A fanout33/X vssd1 vssd1 vccd1 vccd1 _11425_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_8 instruction[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11355_ _11356_/A _11356_/B _11356_/C vssd1 vssd1 vccd1 vccd1 _11355_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_21_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11286_ _11285_/A _11285_/B _11184_/A vssd1 vssd1 vccd1 vccd1 _11286_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07794__A2 _07322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10306_ _10306_/A _10306_/B vssd1 vssd1 vccd1 vccd1 _10308_/B sky130_fd_sc_hd__xnor2_1
X_13025_ _13025_/A _13025_/B vssd1 vssd1 vccd1 vccd1 _13025_/X sky130_fd_sc_hd__xor2_1
X_10237_ _10141_/Y _10235_/Y _10236_/Y vssd1 vssd1 vccd1 vccd1 _10269_/A sky130_fd_sc_hd__o21a_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08743__A1 _06989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06754__B1 _12284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10168_ _08821_/B _10927_/A fanout83/X fanout36/X vssd1 vssd1 vccd1 vccd1 _10169_/B
+ sky130_fd_sc_hd__o22a_1
X_10099_ _09511_/B _10229_/B _09816_/X _10229_/C _10098_/X vssd1 vssd1 vccd1 vccd1
+ _10100_/B sky130_fd_sc_hd__o41a_2
XANTENNA__10440__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12809_ hold258/X hold58/X vssd1 vssd1 vccd1 vccd1 _13097_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_84_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12055__A1 _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10066__B1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08000_ _07756_/B _07782_/B _07756_/A vssd1 vssd1 vccd1 vccd1 _08011_/A sky130_fd_sc_hd__o21ba_2
XANTENNA__12358__A2 _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09759__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09951_ _09952_/B _09952_/A vssd1 vssd1 vccd1 vccd1 _09951_/Y sky130_fd_sc_hd__nand2b_1
X_08902_ _08902_/A _08902_/B vssd1 vssd1 vccd1 vccd1 _08912_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11318__B1 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08734__A1 _07031_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ _10018_/B _09882_/B vssd1 vssd1 vccd1 vccd1 _09919_/A sky130_fd_sc_hd__and2b_1
XANTENNA__11869__A1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11869__B2 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08734__B2 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08833_ _10169_/A _08833_/B vssd1 vssd1 vccd1 vccd1 _08834_/B sky130_fd_sc_hd__xnor2_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout288_A _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08764_ _08764_/A _08764_/B vssd1 vssd1 vccd1 vccd1 _08766_/C sky130_fd_sc_hd__xnor2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07715_ _07727_/A vssd1 vssd1 vccd1 vccd1 _07998_/A sky130_fd_sc_hd__inv_2
XANTENNA__06760__A3 _12583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08695_ _08695_/A _08695_/B vssd1 vssd1 vccd1 vccd1 _08696_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07646_ _07173_/Y _07179_/A _07182_/X _11012_/A vssd1 vssd1 vccd1 vccd1 _07647_/B
+ sky130_fd_sc_hd__a22o_1
X_07577_ _07577_/A _07577_/B vssd1 vssd1 vccd1 vccd1 _07579_/B sky130_fd_sc_hd__xnor2_1
X_09316_ _09316_/A _09316_/B vssd1 vssd1 vccd1 vccd1 _09321_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09247_ _09247_/A _09247_/B vssd1 vssd1 vccd1 vccd1 _09249_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07473__A1 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08670__B1 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07473__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09178_ _09146_/X _09177_/X _10251_/S vssd1 vssd1 vccd1 vccd1 _09178_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09586__A _11695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08129_ _08129_/A _08129_/B vssd1 vssd1 vccd1 vccd1 _08198_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11021__A2 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07776__A2 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11140_ _11262_/C _11140_/B vssd1 vssd1 vccd1 vccd1 _11142_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_31_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11309__B1 _12382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10780__A1 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10780__B2 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08725__A1 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11071_ _10852_/Y _11279_/A _11069_/Y vssd1 vssd1 vccd1 vccd1 _11071_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08725__B2 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10022_ fanout77/X fanout52/X _10677_/B fanout75/X vssd1 vssd1 vccd1 vccd1 _10023_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07553__B _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11973_ _11973_/A _11973_/B vssd1 vssd1 vccd1 vccd1 _11975_/B sky130_fd_sc_hd__or2_1
XFILLER_0_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10924_ _10925_/A _10925_/B _10925_/C vssd1 vssd1 vccd1 vccd1 _10926_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10855_ _11070_/A _10855_/B vssd1 vssd1 vccd1 vccd1 _11215_/A sky130_fd_sc_hd__xor2_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12525_ _12557_/A _12526_/B vssd1 vssd1 vccd1 vccd1 _12525_/X sky130_fd_sc_hd__and2_1
XFILLER_0_94_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10786_ _11935_/A fanout47/X _11603_/A _12772_/A vssd1 vssd1 vccd1 vccd1 _10787_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08661__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11260__A2 _11148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12456_ _12457_/A _12457_/B _12457_/C vssd1 vssd1 vccd1 vccd1 _12464_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12387_ _12387_/A _12387_/B vssd1 vssd1 vccd1 vccd1 _12388_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07216__A1 _12250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11407_ _11360_/A _11360_/B _11361_/X vssd1 vssd1 vccd1 vccd1 _11455_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11338_ fanout29/X _11935_/A _12776_/A fanout32/X vssd1 vssd1 vccd1 vccd1 _11339_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_9_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13311_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__10154__B _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11269_ _11270_/A _11270_/B vssd1 vssd1 vccd1 vccd1 _11369_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_118_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13008_ _11780_/A _13020_/B2 hold119/X vssd1 vssd1 vccd1 vccd1 hold120/A sky130_fd_sc_hd__o21a_1
XANTENNA__07744__A _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07500_ _10155_/A _07500_/B vssd1 vssd1 vccd1 vccd1 _07502_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08480_ _08480_/A _08480_/B vssd1 vssd1 vccd1 vccd1 _08489_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10287__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07431_ _07431_/A vssd1 vssd1 vccd1 vccd1 _07441_/A sky130_fd_sc_hd__inv_2
XFILLER_0_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07362_ _07362_/A _07362_/B vssd1 vssd1 vccd1 vccd1 _07626_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_18_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09101_ _08977_/Y _08990_/A _08990_/B vssd1 vssd1 vccd1 vccd1 _09101_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07293_ _07293_/A _07293_/B vssd1 vssd1 vccd1 vccd1 _07294_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_45_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07455__A1 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07455__B2 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09032_ _09032_/A _09032_/B vssd1 vssd1 vccd1 vccd1 _09079_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_13_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12544__B _12545_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12751__A2 _12980_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout203_A _08311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09934_ _09935_/A _09935_/B vssd1 vssd1 vccd1 vccd1 _09934_/Y sky130_fd_sc_hd__nand2_1
X_09865_ _10169_/A _09865_/B vssd1 vssd1 vccd1 vccd1 _09869_/A sky130_fd_sc_hd__xnor2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _08919_/A _08816_/B vssd1 vssd1 vccd1 vccd1 _08818_/B sky130_fd_sc_hd__nor2_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _09794_/Y _09796_/B vssd1 vssd1 vccd1 vccd1 _09797_/B sky130_fd_sc_hd__and2b_1
X_08747_ _08696_/A _08696_/B _08744_/Y _08745_/X vssd1 vssd1 vccd1 vccd1 _08750_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_68_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _08678_/A _08678_/B _08678_/C vssd1 vssd1 vccd1 vccd1 _08678_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_68_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _07629_/A _07629_/B vssd1 vssd1 vccd1 vccd1 _08941_/B sky130_fd_sc_hd__xor2_2
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10640_ _06728_/B _12243_/B1 _09383_/B _10621_/A _10639_/X vssd1 vssd1 vccd1 vccd1
+ _10641_/C sky130_fd_sc_hd__o221a_1
XFILLER_0_48_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09840__C1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10571_ _10571_/A _10571_/B vssd1 vssd1 vccd1 vccd1 _10573_/B sky130_fd_sc_hd__xor2_4
X_13290_ _13318_/CLK _13290_/D vssd1 vssd1 vccd1 vccd1 hold272/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12310_ _12308_/A _12308_/B _12308_/C vssd1 vssd1 vccd1 vccd1 _12311_/B sky130_fd_sc_hd__o21ai_1
X_12241_ _11398_/B _12285_/B hold270/A vssd1 vssd1 vccd1 vccd1 _12241_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10202__B1 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12172_ _06843_/A _12170_/X _12171_/Y vssd1 vssd1 vccd1 vccd1 _12172_/X sky130_fd_sc_hd__o21a_1
X_11123_ _11499_/A _11123_/B vssd1 vssd1 vccd1 vccd1 _11125_/B sky130_fd_sc_hd__xnor2_1
X_11054_ _11054_/A _11054_/B _11054_/C vssd1 vssd1 vccd1 vccd1 _11055_/B sky130_fd_sc_hd__or3_1
X_10005_ _09950_/A _09950_/B _09951_/Y vssd1 vssd1 vccd1 vccd1 _10091_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__07921__A2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06724__A3 _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11956_ _12032_/B _11956_/B vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__and2_1
XFILLER_0_59_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10907_ _10908_/A _10908_/B vssd1 vssd1 vccd1 vccd1 _11003_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11887_ _11888_/A _11888_/B _11888_/C vssd1 vssd1 vccd1 vccd1 _11890_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_82_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10149__B _11147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11769__B1 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10838_ _10839_/B _10839_/A vssd1 vssd1 vccd1 vccd1 _10953_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_125_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10769_ _11381_/A _10739_/Y _10740_/X _10768_/Y _10738_/Y vssd1 vssd1 vccd1 vccd1
+ _10769_/X sky130_fd_sc_hd__a311o_2
XANTENNA__07437__B2 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07437__A1 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12508_ _12516_/C _12508_/B vssd1 vssd1 vccd1 vccd1 _12515_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_82_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12439_ _12603_/B _12440_/B vssd1 vssd1 vccd1 vccd1 _12450_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10165__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12733__A2 _12980_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout109 _07023_/Y vssd1 vssd1 vccd1 vccd1 _12762_/A sky130_fd_sc_hd__clkbuf_16
X_07980_ _07980_/A _07980_/B _07980_/C vssd1 vssd1 vccd1 vccd1 _07982_/B sky130_fd_sc_hd__or3_1
XANTENNA__12380__A _12560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06931_ reg1_val[31] _09968_/A vssd1 vssd1 vccd1 vccd1 _06931_/X sky130_fd_sc_hd__and2_1
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07474__A _10301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07193__B _10819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09650_ _09650_/A _09650_/B vssd1 vssd1 vccd1 vccd1 _09651_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07373__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06862_ _09202_/A vssd1 vssd1 vccd1 vccd1 _06928_/D sky130_fd_sc_hd__inv_2
X_08601_ _09039_/A _09039_/B _08584_/X vssd1 vssd1 vccd1 vccd1 _09041_/A sky130_fd_sc_hd__a21o_1
X_06793_ reg1_val[4] _10752_/S vssd1 vssd1 vccd1 vccd1 _06793_/X sky130_fd_sc_hd__and2_1
X_09581_ _08681_/A _10927_/A fanout83/X _09295_/A vssd1 vssd1 vccd1 vccd1 _09582_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08532_ _08588_/A _08532_/B vssd1 vssd1 vccd1 vccd1 _08541_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08463_ _09772_/A _09618_/B2 _09618_/A1 _09478_/B2 vssd1 vssd1 vccd1 vccd1 _08464_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_49_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout153_A _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07414_ _07414_/A _07414_/B vssd1 vssd1 vccd1 vccd1 _07696_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_9_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08394_ _08394_/A _08394_/B vssd1 vssd1 vccd1 vccd1 _08421_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10680__B1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07345_ _10557_/B fanout81/X _09295_/B fanout13/X vssd1 vssd1 vccd1 vccd1 _07346_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12972__A2 _12742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13150__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07276_ reg1_val[30] _07276_/B vssd1 vssd1 vccd1 vccd1 _07277_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ _09009_/X _09014_/Y _08457_/X vssd1 vssd1 vccd1 vccd1 _09057_/B sky130_fd_sc_hd__a21o_1
Xhold152 hold152/A vssd1 vssd1 vccd1 vccd1 hold152/X sky130_fd_sc_hd__buf_1
Xhold141 hold141/A vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold130 hold130/A vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07087__C _07087_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold163 hold163/A vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07061__C1 _07052_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold185 hold185/A vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 hold174/A vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06954__A3 _07087_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09917_ _09917_/A _10006_/B _09917_/C vssd1 vssd1 vccd1 vccd1 _09919_/B sky130_fd_sc_hd__or3_1
X_09848_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _09849_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout66_A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _09780_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09779_/Y sky130_fd_sc_hd__nand2_1
X_12790_ _13163_/A hold3/X vssd1 vssd1 vccd1 vccd1 _12891_/B sky130_fd_sc_hd__or2_1
X_11810_ _11810_/A _11810_/B vssd1 vssd1 vccd1 vccd1 _11967_/A sky130_fd_sc_hd__nor2_2
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ reg1_val[21] curr_PC[21] vssd1 vssd1 vccd1 vccd1 _11743_/A sky130_fd_sc_hd__nand2_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11672_ curr_PC[19] _11671_/C curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11673_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__10671__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10623_ reg1_val[10] curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10625_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10554_ _06989_/A _11782_/A fanout69/X vssd1 vssd1 vccd1 vccd1 _10555_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_24_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07559__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13273_ _13277_/CLK _13273_/D vssd1 vssd1 vccd1 vccd1 hold130/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07278__B _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10485_ _10485_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10730_/A sky130_fd_sc_hd__xnor2_4
X_12224_ _12317_/A _12222_/X _12223_/Y vssd1 vssd1 vccd1 vccd1 _12224_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_102_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11923__B1 _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12155_ _12083_/A _12083_/B _12084_/X vssd1 vssd1 vccd1 vccd1 _12157_/B sky130_fd_sc_hd__a21o_1
X_11106_ _11076_/X _11079_/Y _11083_/X _11105_/X _06898_/C vssd1 vssd1 vccd1 vccd1
+ _11106_/X sky130_fd_sc_hd__a41o_2
XFILLER_0_75_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12086_ _12203_/A fanout15/X fanout6/X _12150_/A vssd1 vssd1 vccd1 vccd1 _12088_/A
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09895__A2 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11037_ _11429_/A _11037_/B vssd1 vssd1 vccd1 vccd1 _11041_/A sky130_fd_sc_hd__xnor2_1
X_12988_ _10819_/A _13020_/B2 hold91/X vssd1 vssd1 vccd1 vccd1 _13264_/D sky130_fd_sc_hd__o21a_1
XANTENNA__07658__A1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07658__B2 _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11939_ _11939_/A _11939_/B vssd1 vssd1 vccd1 vccd1 _11958_/A sky130_fd_sc_hd__and2_1
XFILLER_0_86_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08853__A _08853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11206__A2 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07130_ _07434_/A _07153_/A vssd1 vssd1 vccd1 vccd1 _07130_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08572__B _08572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07469__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07061_ _07303_/B _07129_/B _07059_/Y _07052_/B vssd1 vssd1 vccd1 vccd1 _07062_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_70_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12167__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07963_ _07964_/A _07964_/B vssd1 vssd1 vccd1 vccd1 _07963_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06914_ instruction[22] _06552_/X _06913_/X _06678_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[4]
+ sky130_fd_sc_hd__o211a_4
X_07894_ _07894_/A _07894_/B vssd1 vssd1 vccd1 vccd1 _07897_/B sky130_fd_sc_hd__xnor2_1
X_09702_ _09842_/B _09841_/B hold246/A vssd1 vssd1 vccd1 vccd1 _09702_/Y sky130_fd_sc_hd__a21oi_1
X_06845_ _06845_/A _06845_/B vssd1 vssd1 vccd1 vccd1 _06845_/Y sky130_fd_sc_hd__nor2_1
X_09633_ _09634_/A _09634_/B vssd1 vssd1 vccd1 vccd1 _09633_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__13145__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09564_ _10064_/B2 _07389_/B fanout26/X _09888_/B2 vssd1 vssd1 vccd1 vccd1 _09565_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06776_ reg1_val[2] _07279_/A vssd1 vssd1 vccd1 vccd1 _06777_/B sky130_fd_sc_hd__nand2_1
X_08515_ _09467_/A _08515_/B vssd1 vssd1 vccd1 vccd1 _08516_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09495_ _09495_/A _09495_/B vssd1 vssd1 vccd1 vccd1 _09496_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_93_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08310__A2 _10551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08446_ _08473_/A _08444_/Y _08441_/Y vssd1 vssd1 vccd1 vccd1 _08453_/B sky130_fd_sc_hd__a21o_1
X_08377_ _08775_/A _08377_/B vssd1 vssd1 vccd1 vccd1 _08383_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07328_ _07329_/A _07329_/B vssd1 vssd1 vccd1 vccd1 _07479_/A sky130_fd_sc_hd__and2_1
XFILLER_0_18_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07259_ _11125_/A _07259_/B vssd1 vssd1 vccd1 vccd1 _07260_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10270_ curr_PC[7] _10397_/C vssd1 vssd1 vccd1 vccd1 _10270_/X sky130_fd_sc_hd__or2_1
XFILLER_0_103_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11669__C1 _11643_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ hold187/X _12947_/A2 _12947_/B1 hold198/X vssd1 vssd1 vccd1 vccd1 hold199/A
+ sky130_fd_sc_hd__a22o_1
X_12842_ _13052_/A _13053_/A _13052_/B vssd1 vssd1 vccd1 vccd1 _13058_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_96_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12773_ hold15/X _12778_/B _12772_/Y _13147_/A vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__o211a_1
XFILLER_0_96_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08837__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11724_ _11635_/B _11812_/A vssd1 vssd1 vccd1 vccd1 _11893_/A sky130_fd_sc_hd__nand2b_1
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11655_ _11746_/A _11655_/B vssd1 vssd1 vccd1 vccd1 _11655_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06905__B _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout80 _06982_/Y vssd1 vssd1 vccd1 vccd1 _08681_/A sky130_fd_sc_hd__buf_4
XFILLER_0_36_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout91 _07197_/Y vssd1 vssd1 vccd1 vccd1 _10927_/A sky130_fd_sc_hd__buf_8
XANTENNA__08065__A1 _08018_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11586_ _11586_/A _11586_/B vssd1 vssd1 vccd1 vccd1 _11730_/C sky130_fd_sc_hd__or2_1
XANTENNA__09262__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10606_ _10606_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _10730_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_101_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13325_ instruction[5] vssd1 vssd1 vccd1 vccd1 loadstore_size[0] sky130_fd_sc_hd__buf_12
X_10537_ _12019_/A _10537_/B vssd1 vssd1 vccd1 vccd1 _10539_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_12_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13256_ _13264_/CLK hold123/X vssd1 vssd1 vccd1 vccd1 _13256_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12149__B1 _09252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10468_ _10468_/A _10468_/B vssd1 vssd1 vccd1 vccd1 _10481_/A sky130_fd_sc_hd__nor2_2
X_12207_ _12208_/A _12258_/B vssd1 vssd1 vccd1 vccd1 _12264_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_32_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13187_ _13280_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
X_10399_ _10646_/C _10399_/B vssd1 vssd1 vccd1 vccd1 _10399_/Y sky130_fd_sc_hd__nor2_1
X_12138_ _12556_/S _12135_/X _12139_/B _12137_/X vssd1 vssd1 vccd1 vccd1 dest_val[26]
+ sky130_fd_sc_hd__a22o_4
X_12069_ curr_PC[25] _12069_/B vssd1 vssd1 vccd1 vccd1 _12069_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07879__A1 _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ reg1_val[30] _07434_/B vssd1 vssd1 vccd1 vccd1 _06631_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11675__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06561_ instruction[19] _06915_/B vssd1 vssd1 vccd1 vccd1 _06561_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08300_ _08301_/A _08301_/B vssd1 vssd1 vccd1 vccd1 _08300_/Y sky130_fd_sc_hd__nor2_1
X_09280_ _09280_/A _09280_/B vssd1 vssd1 vccd1 vccd1 _09281_/B sky130_fd_sc_hd__xnor2_4
X_08231_ _12734_/A _08420_/B _07035_/X _08819_/B2 vssd1 vssd1 vccd1 vccd1 _08232_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08162_ _08209_/A _08209_/B _08122_/X vssd1 vssd1 vccd1 vccd1 _08635_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__12927__A2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07199__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08093_ _08841_/B2 _08420_/B _08854_/B2 _08837_/B2 vssd1 vssd1 vccd1 vccd1 _08094_/B
+ sky130_fd_sc_hd__o22a_1
X_07113_ _07128_/B _07128_/C _07135_/B vssd1 vssd1 vccd1 vccd1 _07114_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_43_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07044_ _09898_/A _07046_/B vssd1 vssd1 vccd1 vccd1 _07047_/A sky130_fd_sc_hd__and2_1
XFILLER_0_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout116_A _11780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11902__A3 _09076_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ _08995_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _09660_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_11_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07946_ _10015_/A _07946_/B vssd1 vssd1 vccd1 vccd1 _07948_/B sky130_fd_sc_hd__xnor2_2
X_07877_ _07974_/A _07877_/B vssd1 vssd1 vccd1 vccd1 _07935_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__11184__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08477__B _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06828_ _11739_/A _06827_/Y _06826_/Y vssd1 vssd1 vccd1 vccd1 _06829_/B sky130_fd_sc_hd__o21a_1
X_09616_ _09615_/B _09616_/B vssd1 vssd1 vccd1 vccd1 _09617_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_78_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08819__B1 _09295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09547_ _06870_/A _09545_/X _09546_/Y vssd1 vssd1 vccd1 vccd1 _09547_/Y sky130_fd_sc_hd__o21ai_1
X_06759_ reg2_val[4] _06778_/B vssd1 vssd1 vccd1 vccd1 _06759_/X sky130_fd_sc_hd__and2_1
XFILLER_0_93_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09478_ _09772_/A _07278_/B fanout7/X _09478_/B2 vssd1 vssd1 vccd1 vccd1 _09479_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout29_A _07006_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_11_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13264_/CLK sky130_fd_sc_hd__clkbuf_8
X_08429_ _08427_/A _08427_/B _08428_/X vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10528__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08047__B2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08047__A1 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ _11351_/A _11351_/B _11341_/Y vssd1 vssd1 vccd1 vccd1 _11451_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11371_ _11170_/Y _11275_/A _11275_/B vssd1 vssd1 vccd1 vccd1 _11371_/X sky130_fd_sc_hd__o21ba_1
X_13110_ hold289/X _13165_/A2 _13109_/X _13146_/B2 vssd1 vssd1 vccd1 vccd1 hold290/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09528__S _10249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ _10323_/A _10323_/B vssd1 vssd1 vccd1 vccd1 _10473_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_21_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13041_ hold288/X _12721_/B _13040_/X _12722_/A vssd1 vssd1 vccd1 vccd1 _13042_/B
+ sky130_fd_sc_hd__a22o_1
X_10253_ _12124_/B _10509_/C _13224_/Q vssd1 vssd1 vccd1 vccd1 _10253_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07558__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10184_ _10184_/A _10184_/B vssd1 vssd1 vccd1 vccd1 _10185_/B sky130_fd_sc_hd__xnor2_1
Xfanout270 hold152/X vssd1 vssd1 vccd1 vccd1 _13168_/A2 sky130_fd_sc_hd__buf_2
Xfanout292 _13028_/A vssd1 vssd1 vccd1 vccd1 _13013_/C1 sky130_fd_sc_hd__buf_4
XANTENNA__11106__A1 _11076_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout281 _06569_/X vssd1 vssd1 vccd1 vccd1 _06729_/B sky130_fd_sc_hd__buf_2
XANTENNA__07572__A _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12825_ _12823_/X _12825_/B vssd1 vssd1 vccd1 vccd1 _13039_/A sky130_fd_sc_hd__nand2b_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12756_ hold65/X _12786_/B vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__or2_1
XFILLER_0_84_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12637__B _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12687_ _12685_/X _12687_/B vssd1 vssd1 vccd1 vccd1 _12698_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__10438__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11707_ _11797_/A _11707_/B vssd1 vssd1 vccd1 vccd1 _11709_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_114_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08038__B2 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08038__A1 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11638_ _11638_/A _11638_/B vssd1 vssd1 vccd1 vccd1 _11638_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_126_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13308_ _13309_/CLK _13308_/D vssd1 vssd1 vccd1 vccd1 hold254/A sky130_fd_sc_hd__dfxtp_1
X_11569_ _10883_/Y _11568_/Y _11831_/S vssd1 vssd1 vccd1 vccd1 _11569_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13239_ _13241_/CLK hold202/X vssd1 vssd1 vccd1 vccd1 hold200/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11345__A1 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11345__B2 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07800_ _09580_/A _07800_/B vssd1 vssd1 vccd1 vccd1 _07801_/B sky130_fd_sc_hd__xnor2_1
X_08780_ _08780_/A _08780_/B vssd1 vssd1 vccd1 vccd1 _08782_/A sky130_fd_sc_hd__xor2_2
X_07731_ _08837_/B2 _08134_/B fanout51/X _12736_/A vssd1 vssd1 vccd1 vccd1 _07732_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07662_ _07687_/B _07662_/B vssd1 vssd1 vccd1 vccd1 _08903_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09710__A1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10856__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06613_ instruction[36] _06633_/B vssd1 vssd1 vccd1 vccd1 _12614_/B sky130_fd_sc_hd__and2_4
XANTENNA__12058__C1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09401_ curr_PC[0] curr_PC[1] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09402_/B sky130_fd_sc_hd__a21oi_1
X_07593_ _07593_/A _07593_/B vssd1 vssd1 vccd1 vccd1 _07595_/C sky130_fd_sc_hd__xor2_1
X_09332_ _07705_/X _08994_/Y _07706_/X vssd1 vssd1 vccd1 vccd1 _09332_/X sky130_fd_sc_hd__a21o_1
X_06544_ reg1_val[26] vssd1 vssd1 vccd1 vccd1 _06956_/A sky130_fd_sc_hd__inv_2
XFILLER_0_118_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout233_A _09384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09263_ _10894_/A _09263_/B vssd1 vssd1 vccd1 vccd1 _09267_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08214_ _08253_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _08214_/Y sky130_fd_sc_hd__nor2_1
X_09194_ _09200_/A _09200_/B _09201_/B vssd1 vssd1 vccd1 vccd1 _09194_/Y sky130_fd_sc_hd__nor3_4
XFILLER_0_16_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08145_ _08203_/A _08203_/B _08141_/X vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_105_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07657__A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12563__A _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08076_ _08394_/A _08076_/B vssd1 vssd1 vccd1 vccd1 _08133_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07027_ _07105_/A _07027_/B vssd1 vssd1 vccd1 vccd1 _07028_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09872__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _08978_/A _08978_/B vssd1 vssd1 vccd1 vccd1 _09102_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__10811__A _10811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07929_ _08024_/A _08024_/B _07910_/Y vssd1 vssd1 vccd1 vccd1 _07939_/B sky130_fd_sc_hd__o21ai_2
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
X_10940_ _10826_/A _10825_/B _10825_/A vssd1 vssd1 vccd1 vccd1 _10945_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07712__B1 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10871_ _10868_/Y _10869_/X _10747_/A _10749_/X vssd1 vssd1 vccd1 vccd1 _10871_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_78_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12610_ _12611_/A _12611_/C _12611_/B vssd1 vssd1 vccd1 vccd1 _12617_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_93_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12064__A2 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12541_ _12541_/A _12541_/B _12541_/C _12541_/D vssd1 vssd1 vccd1 vccd1 _12542_/B
+ sky130_fd_sc_hd__and4_2
X_12472_ _12478_/B _12472_/B vssd1 vssd1 vccd1 vccd1 new_PC[13] sky130_fd_sc_hd__and2_4
XFILLER_0_81_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11423_ _11532_/A _11423_/B vssd1 vssd1 vccd1 vccd1 _11427_/A sky130_fd_sc_hd__and2_1
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10378__A2 _06928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_9 reg1_val[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11354_ _11354_/A _11354_/B vssd1 vssd1 vccd1 vccd1 _11356_/C sky130_fd_sc_hd__or2_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11285_ _11285_/A _11285_/B vssd1 vssd1 vccd1 vccd1 _11285_/X sky130_fd_sc_hd__or2_1
XANTENNA__07794__A3 _07322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ _08680_/B _11134_/B2 fanout57/X fanout30/X vssd1 vssd1 vccd1 vccd1 _10306_/B
+ sky130_fd_sc_hd__o22a_1
X_13024_ _13028_/A hold241/X vssd1 vssd1 vccd1 vccd1 _13281_/D sky130_fd_sc_hd__and2_1
X_10236_ _10141_/Y _10235_/Y _09110_/X vssd1 vssd1 vccd1 vccd1 _10236_/Y sky130_fd_sc_hd__a21oi_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08743__A2 _11782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ _10167_/A _10167_/B vssd1 vssd1 vccd1 vccd1 _10171_/B sky130_fd_sc_hd__xor2_1
X_10098_ _09815_/X _10096_/X _10097_/Y vssd1 vssd1 vccd1 vccd1 _10098_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_107_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_202 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12808_ hold294/A hold11/X vssd1 vssd1 vccd1 vccd1 _13102_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09456__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12739_ _10035_/A _12980_/A2 hold78/X _13028_/A vssd1 vssd1 vccd1 vccd1 _13191_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10066__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10066__A1 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09471__A3 _07435_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13004__A1 _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09759__A1 _10553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12383__A _12563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09759__B2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09950_ _09950_/A _09950_/B vssd1 vssd1 vccd1 vccd1 _09952_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08901_ _08902_/B _08902_/A vssd1 vssd1 vccd1 vccd1 _08950_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11318__B2 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11318__A1 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08734__A2 _07179_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _09881_/A _09881_/B _09879_/Y vssd1 vssd1 vccd1 vccd1 _09882_/B sky130_fd_sc_hd__or3b_1
XANTENNA__11869__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08832_ _10169_/A _08833_/B vssd1 vssd1 vccd1 vccd1 _08832_/Y sky130_fd_sc_hd__nand2_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ _08764_/A _08764_/B vssd1 vssd1 vccd1 vccd1 _08870_/A sky130_fd_sc_hd__and2b_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07714_ _07716_/A _07716_/B _07716_/C vssd1 vssd1 vccd1 vccd1 _07727_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout183_A _08415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08694_ _07134_/A _10557_/A _07119_/Y _07869_/B vssd1 vssd1 vccd1 vccd1 _08695_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07645_ _08857_/A _07645_/B vssd1 vssd1 vccd1 vccd1 _07648_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09447__B1 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07576_ _07576_/A _07576_/B vssd1 vssd1 vccd1 vccd1 _07577_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10057__A1 _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09315_ _07581_/A _07580_/B _07578_/Y vssd1 vssd1 vccd1 vccd1 _09325_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_8_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09867__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09246_ _09247_/A _09247_/B vssd1 vssd1 vccd1 vccd1 _09418_/A sky130_fd_sc_hd__or2_1
XFILLER_0_118_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08670__B2 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08670__A1 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07473__A2 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06681__B1 _06569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ _09161_/X _09176_/X _11089_/A vssd1 vssd1 vccd1 vccd1 _09177_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08128_ _08129_/A _08129_/B vssd1 vssd1 vccd1 vccd1 _08128_/X sky130_fd_sc_hd__or2_1
XFILLER_0_16_496 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08059_ _08059_/A _08120_/A vssd1 vssd1 vccd1 vccd1 _08069_/A sky130_fd_sc_hd__nand2_2
XANTENNA_fanout96_A _08672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10780__A2 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ _11070_/A _11173_/A vssd1 vssd1 vccd1 vccd1 _11279_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12740__B _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08186__B1 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10021_ _09870_/B _09873_/B _09870_/A vssd1 vssd1 vccd1 vccd1 _10033_/A sky130_fd_sc_hd__o21bai_1
XANTENNA__08725__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09107__A _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11972_ _11972_/A _11972_/B _11972_/C _11972_/D vssd1 vssd1 vccd1 vccd1 _11973_/B
+ sky130_fd_sc_hd__and4_2
XANTENNA__12468__A _12626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10923_ _12255_/B _10923_/B vssd1 vssd1 vccd1 vccd1 _10925_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10854_ _09818_/B _10362_/Y _10850_/Y _10851_/Y _10853_/Y vssd1 vssd1 vccd1 vccd1
+ _10855_/B sky130_fd_sc_hd__o311a_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11245__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ reg1_val[22] curr_PC[22] _12524_/S vssd1 vssd1 vccd1 vccd1 _12526_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10785_ _11429_/A _10785_/B vssd1 vssd1 vccd1 vccd1 _10789_/A sky130_fd_sc_hd__xnor2_1
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08681__A _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__B2 _06952_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__A1 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06913__B _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12455_ _12464_/A _12455_/B vssd1 vssd1 vccd1 vccd1 _12457_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06672__B1 _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12386_ _12387_/A _12387_/B vssd1 vssd1 vccd1 vccd1 _12394_/B sky130_fd_sc_hd__or2_1
XFILLER_0_50_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11406_ _11730_/A _11730_/B _12230_/A vssd1 vssd1 vccd1 vccd1 _11406_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_120_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11337_ _11337_/A _11337_/B vssd1 vssd1 vccd1 vccd1 _11340_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08177__B1 _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11268_ _11268_/A _11268_/B vssd1 vssd1 vccd1 vccd1 _11270_/B sky130_fd_sc_hd__xnor2_1
X_11199_ hold258/A _11398_/B _11296_/B vssd1 vssd1 vccd1 vccd1 _11199_/X sky130_fd_sc_hd__and3_1
X_13007_ hold130/A _13013_/A2 _13020_/A2 hold118/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold119/A sky130_fd_sc_hd__o221a_1
X_10219_ _10220_/B _10220_/A vssd1 vssd1 vccd1 vccd1 _10219_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07760__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10287__A1 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10287__B2 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07430_ _09622_/A _07430_/B vssd1 vssd1 vccd1 vccd1 _07431_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09429__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07361_ _07362_/A _07362_/B vssd1 vssd1 vccd1 vccd1 _07361_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09100_ _09507_/B _09100_/B vssd1 vssd1 vccd1 vccd1 _12326_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_128_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09031_ _09031_/A _09031_/B vssd1 vssd1 vccd1 vccd1 _09032_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_60_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07292_ _07293_/A _07293_/B vssd1 vssd1 vccd1 vccd1 _07601_/B sky130_fd_sc_hd__and2_1
XFILLER_0_5_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07455__A2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold301 hold301/A vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06966__A1 _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09933_ _08544_/A _08544_/B _10551_/B _09778_/B _09776_/X vssd1 vssd1 vccd1 vccd1
+ _09935_/B sky130_fd_sc_hd__a41o_1
XFILLER_0_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12560__B _12560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09864_ _08821_/B fanout81/X _09295_/B fanout36/X vssd1 vssd1 vccd1 vccd1 _09865_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08815_ _08815_/A _08815_/B _08815_/C vssd1 vssd1 vccd1 vccd1 _08816_/B sky130_fd_sc_hd__and3_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _09795_/A _09795_/B vssd1 vssd1 vccd1 vccd1 _09796_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_84_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08746_ _08744_/Y _08745_/X _08696_/A _08696_/B vssd1 vssd1 vccd1 vccd1 _08864_/A
+ sky130_fd_sc_hd__a211o_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _08677_/A _08677_/B _08677_/C vssd1 vssd1 vccd1 vccd1 _08678_/C sky130_fd_sc_hd__nand3_1
XANTENNA__07143__A1 _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07628_ _07628_/A _07628_/B vssd1 vssd1 vccd1 vccd1 _08941_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11227__B1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07559_ _10555_/A _07559_/B _07559_/C vssd1 vssd1 vccd1 vccd1 _07562_/C sky130_fd_sc_hd__and3_1
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout11_A _07322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10570_ _10570_/A _10570_/B vssd1 vssd1 vccd1 vccd1 _10571_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_91_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09229_ _10280_/A _09229_/B vssd1 vssd1 vccd1 vccd1 _09232_/A sky130_fd_sc_hd__xnor2_2
X_12240_ hold254/A _12240_/B vssd1 vssd1 vccd1 vccd1 _12285_/B sky130_fd_sc_hd__or2_1
XFILLER_0_32_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12171_ _06843_/A _12170_/X _12277_/B1 vssd1 vssd1 vccd1 vccd1 _12171_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10202__B2 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10202__A1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11122_ fanout19/X _10557_/B fanout13/X _12203_/A vssd1 vssd1 vccd1 vccd1 _11123_/B
+ sky130_fd_sc_hd__o22a_1
X_11053_ _11054_/A _11054_/B _11054_/C vssd1 vssd1 vccd1 vccd1 _11055_/A sky130_fd_sc_hd__o21ai_1
X_10004_ _09955_/A _09955_/B _09953_/Y vssd1 vssd1 vccd1 vccd1 _10094_/A sky130_fd_sc_hd__a21boi_4
XFILLER_0_99_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11955_ _11955_/A _11955_/B _11955_/C vssd1 vssd1 vccd1 vccd1 _11956_/B sky130_fd_sc_hd__or3_1
XFILLER_0_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10906_ _12022_/A _10906_/B vssd1 vssd1 vccd1 vccd1 _10908_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11886_ _11886_/A _11886_/B vssd1 vssd1 vccd1 vccd1 _11888_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11769__A1 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11769__B2 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10837_ _10837_/A _10837_/B vssd1 vssd1 vccd1 vccd1 _10839_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10768_ _10743_/Y _10744_/X _10767_/X vssd1 vssd1 vccd1 vccd1 _10768_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07437__A2 _12786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12507_ _12551_/A _12507_/B vssd1 vssd1 vccd1 vccd1 _12508_/B sky130_fd_sc_hd__or2_1
XFILLER_0_82_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09300__A _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12438_ reg1_val[9] curr_PC[9] _12524_/S vssd1 vssd1 vccd1 vccd1 _12440_/B sky130_fd_sc_hd__mux2_1
X_10699_ _10699_/A _10832_/A _10699_/C vssd1 vssd1 vccd1 vccd1 _10700_/A sky130_fd_sc_hd__and3_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12369_ reg1_val[31] _10377_/B _12250_/B vssd1 vssd1 vccd1 vccd1 _12369_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06930_ _06928_/D _09202_/B _12250_/B vssd1 vssd1 vccd1 vccd1 _06930_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07373__B2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07373__A1 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06861_ instruction[4] instruction[3] vssd1 vssd1 vccd1 vccd1 _09202_/A sky130_fd_sc_hd__or2_4
X_08600_ _09034_/A _09037_/A _08599_/Y _08597_/B vssd1 vssd1 vccd1 vccd1 _09039_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_89_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06792_ _06770_/X _06790_/Y _06791_/Y vssd1 vssd1 vccd1 vccd1 _06792_/Y sky130_fd_sc_hd__o21ai_1
X_09580_ _09580_/A _09580_/B vssd1 vssd1 vccd1 vccd1 _09584_/A sky130_fd_sc_hd__xnor2_1
X_08531_ _08531_/A _08531_/B _08531_/C vssd1 vssd1 vccd1 vccd1 _08538_/A sky130_fd_sc_hd__and3_1
XANTENNA__07490__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08462_ _08482_/A _08482_/B vssd1 vssd1 vccd1 vccd1 _08485_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_54_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07413_ _07625_/A _07625_/B _07410_/Y vssd1 vssd1 vccd1 vccd1 _07696_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_58_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10680__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout146_A _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08393_ _09180_/A _10551_/A _07325_/Y _08544_/C vssd1 vssd1 vccd1 vccd1 _08394_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10680__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12957__B1 _12980_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07344_ _07344_/A _07344_/B vssd1 vssd1 vccd1 vccd1 _07387_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09822__B1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09210__A _10249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07275_ reg1_val[29] _07528_/C _07165_/A vssd1 vssd1 vccd1 vccd1 _07276_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_33_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06553__B _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09014_ _09010_/Y _09050_/A _08503_/Y _09054_/A vssd1 vssd1 vccd1 vccd1 _09014_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold153 hold153/A vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 hold142/A vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07087__D _12697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 hold197/A vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
X_09916_ _10006_/A _09915_/B _09900_/Y vssd1 vssd1 vccd1 vccd1 _09917_/C sky130_fd_sc_hd__o21ba_1
XFILLER_0_0_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09847_ reg1_val[4] curr_PC[4] vssd1 vssd1 vccd1 vccd1 _09847_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11696__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ _09778_/A _09778_/B vssd1 vssd1 vccd1 vccd1 _09780_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout59_A _07157_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08729_ _10064_/B2 _09752_/B fanout14/X _08837_/B2 vssd1 vssd1 vccd1 vccd1 _08730_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07116__A1 _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _11739_/A _11739_/B _12277_/B1 vssd1 vssd1 vccd1 vccd1 _11740_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_68_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11999__A1 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ curr_PC[19] curr_PC[20] _11671_/C vssd1 vssd1 vccd1 vccd1 _11764_/B sky130_fd_sc_hd__and3_1
XANTENNA__10671__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10671__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10622_ _10621_/A _10621_/B _10621_/Y _12277_/B1 vssd1 vssd1 vccd1 vccd1 _10622_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06627__B1 _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10553_ _10553_/A _10553_/B vssd1 vssd1 vccd1 vccd1 _10555_/B sky130_fd_sc_hd__or2_1
XFILLER_0_24_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13272_ _13277_/CLK hold102/X vssd1 vssd1 vccd1 vccd1 hold100/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _10485_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10484_/X sky130_fd_sc_hd__and2_1
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12481__A _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12223_ _12317_/A _12222_/X _12223_/B1 vssd1 vssd1 vccd1 vccd1 _12223_/Y sky130_fd_sc_hd__o21ai_1
X_12154_ _12154_/A _12154_/B vssd1 vssd1 vccd1 vccd1 _12157_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11105_ _09184_/X _11092_/A _11093_/X _09205_/B _11104_/Y vssd1 vssd1 vccd1 vccd1
+ _11105_/X sky130_fd_sc_hd__o221a_1
X_12085_ _12085_/A _12085_/B vssd1 vssd1 vccd1 vccd1 _12090_/A sky130_fd_sc_hd__xnor2_1
X_11036_ _12301_/A fanout52/X _10677_/B _12784_/A vssd1 vssd1 vccd1 vccd1 _11037_/B
+ sky130_fd_sc_hd__o22a_1
X_12987_ hold90/X _13013_/A2 _13020_/A2 hold42/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold91/A sky130_fd_sc_hd__o221a_1
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07658__A2 _09295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11938_ _11938_/A _11938_/B _11938_/C vssd1 vssd1 vccd1 vccd1 _11939_/B sky130_fd_sc_hd__or3_1
X_11869_ fanout27/X _12150_/A _12150_/B _12205_/A vssd1 vssd1 vccd1 vccd1 _11870_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07060_ _06653_/B _07129_/B _07303_/B _07052_/B vssd1 vssd1 vccd1 vccd1 _07062_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07115__C_N _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12391__A _12568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11914__A1 _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07962_ _08773_/A _07962_/B vssd1 vssd1 vccd1 vccd1 _07964_/B sky130_fd_sc_hd__xnor2_2
X_09701_ hold250/A hold279/A hold240/A vssd1 vssd1 vccd1 vccd1 _09841_/B sky130_fd_sc_hd__or3_1
XANTENNA__10115__S _10249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06913_ instruction[29] _06915_/B vssd1 vssd1 vccd1 vccd1 _06913_/X sky130_fd_sc_hd__or2_1
X_07893_ _07004_/X _08217_/B fanout55/X _12734_/A vssd1 vssd1 vccd1 vccd1 _07894_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_4_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08543__B1 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06844_ _06837_/Y _06843_/Y _06605_/B vssd1 vssd1 vccd1 vccd1 _06845_/B sky130_fd_sc_hd__a21oi_1
X_09632_ _09632_/A _09632_/B vssd1 vssd1 vccd1 vccd1 _09634_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09205__A _12713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09563_ _09475_/A _09475_/B _09473_/Y vssd1 vssd1 vccd1 vccd1 _09577_/A sky130_fd_sc_hd__a21bo_2
XANTENNA_fanout263_A _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06775_ reg1_val[2] _07279_/A vssd1 vssd1 vccd1 vccd1 _09694_/A sky130_fd_sc_hd__nor2_1
X_08514_ _09478_/B2 _09618_/B2 _09618_/A1 _09476_/A vssd1 vssd1 vccd1 vccd1 _08515_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12642__A2 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09494_ _09495_/A _09495_/B vssd1 vssd1 vccd1 vccd1 _09494_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_93_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08445_ _08445_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08473_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10653__A1 _10551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11850__B1 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08376_ _10064_/B2 _08774_/A2 _08774_/B1 _08837_/B2 vssd1 vssd1 vccd1 vccd1 _08377_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11470__A _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06609__B1 _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07327_ _10565_/A _07327_/B vssd1 vssd1 vccd1 vccd1 _07329_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07258_ _11125_/A _07259_/B vssd1 vssd1 vccd1 vccd1 _07261_/B sky130_fd_sc_hd__or2_1
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07189_ reg1_val[14] _07189_/B vssd1 vssd1 vccd1 vccd1 _07194_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_60_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11905__A1 _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07395__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12910_ _12946_/A hold188/X vssd1 vssd1 vccd1 vccd1 _13225_/D sky130_fd_sc_hd__and2_1
X_12841_ hold56/X hold266/X vssd1 vssd1 vccd1 vccd1 _13052_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09115__A _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12772_ _12772_/A _12778_/B vssd1 vssd1 vccd1 vccd1 _12772_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08837__B2 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08837__A1 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10644__A1 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11723_ _11723_/A _11723_/B vssd1 vssd1 vccd1 vccd1 _11892_/A sky130_fd_sc_hd__nor2_2
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11654_ _11654_/A _11654_/B vssd1 vssd1 vccd1 vccd1 _11655_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout92 _07197_/Y vssd1 vssd1 vccd1 vccd1 _12752_/A sky130_fd_sc_hd__buf_6
Xfanout70 _07078_/X vssd1 vssd1 vccd1 vccd1 fanout70/X sky130_fd_sc_hd__buf_8
Xfanout81 _07312_/X vssd1 vssd1 vccd1 vccd1 fanout81/X sky130_fd_sc_hd__buf_6
XFILLER_0_52_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10605_ _10606_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _10605_/X sky130_fd_sc_hd__and2_1
XFILLER_0_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11585_ _12382_/S _11582_/X _11583_/X _11584_/Y vssd1 vssd1 vccd1 vccd1 dest_val[19]
+ sky130_fd_sc_hd__a22o_4
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09262__B2 _10553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09262__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13324_ instruction[16] vssd1 vssd1 vccd1 vccd1 loadstore_dest[5] sky130_fd_sc_hd__buf_12
XFILLER_0_107_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_26 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12149__A1 _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10536_ fanout32/X _11431_/A _11347_/A fanout29/X vssd1 vssd1 vccd1 vccd1 _10537_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13255_ _13289_/CLK _13255_/D vssd1 vssd1 vccd1 vccd1 hold121/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10467_ _10466_/B _10466_/C _10466_/A vssd1 vssd1 vccd1 vccd1 _10468_/B sky130_fd_sc_hd__a21oi_1
X_12206_ _12206_/A _12206_/B vssd1 vssd1 vccd1 vccd1 _12258_/B sky130_fd_sc_hd__xnor2_1
X_13186_ _13280_/CLK _13186_/D vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfxtp_1
X_10398_ curr_PC[7] _10397_/C curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10399_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12137_ curr_PC[26] _12136_/B _10400_/S vssd1 vssd1 vccd1 vccd1 _12137_/X sky130_fd_sc_hd__o21a_1
X_12068_ _12042_/X _12046_/X _12067_/X _12345_/A vssd1 vssd1 vccd1 vccd1 _12068_/X
+ sky130_fd_sc_hd__a31o_1
X_11019_ _12203_/A _10557_/B fanout13/X _12150_/A vssd1 vssd1 vccd1 vccd1 _11020_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06649__A _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06560_ instruction[11] _06552_/X _06559_/X _06678_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[0]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08230_ _08240_/A _08240_/B vssd1 vssd1 vccd1 vccd1 _08230_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09203__A1_N _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08161_ _08161_/A _08161_/B vssd1 vssd1 vccd1 vccd1 _08209_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08092_ _08091_/A _08151_/A _08103_/A vssd1 vssd1 vccd1 vccd1 _08092_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_113_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07112_ _07112_/A _07112_/B _07111_/C vssd1 vssd1 vccd1 vccd1 _07129_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_70_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07043_ reg1_val[6] _07043_/B vssd1 vssd1 vccd1 vccd1 _07046_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout109_A _07023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11899__B1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08994_ _08995_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _08994_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07945_ _08821_/A _09295_/A _08825_/A2 _08681_/A vssd1 vssd1 vccd1 vccd1 _07946_/B
+ sky130_fd_sc_hd__o22a_1
X_07876_ _07874_/Y _07876_/B _07935_/A vssd1 vssd1 vccd1 vccd1 _07935_/B sky130_fd_sc_hd__nand3b_2
XANTENNA__07154__S _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09615_ _09616_/B _09615_/B vssd1 vssd1 vccd1 vccd1 _09736_/D sky130_fd_sc_hd__and2b_1
XFILLER_0_92_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06827_ reg1_val[20] _07068_/A vssd1 vssd1 vccd1 vccd1 _06827_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08819__B2 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08819__A1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06758_ _06758_/A _06758_/B vssd1 vssd1 vccd1 vccd1 _09970_/A sky130_fd_sc_hd__and2_1
X_09546_ _06870_/A _09545_/X _12277_/B1 vssd1 vssd1 vccd1 vccd1 _09546_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12076__B1 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09477_ _09275_/Y _09280_/B _09278_/Y vssd1 vssd1 vccd1 vccd1 _09481_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_93_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06689_ _06687_/Y _06680_/B1 _06752_/A reg2_val[16] vssd1 vssd1 vccd1 vccd1 _07168_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_08428_ _08456_/B _08456_/A vssd1 vssd1 vccd1 vccd1 _08428_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08047__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08359_ _08359_/A _08359_/B vssd1 vssd1 vccd1 vccd1 _08360_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11370_ _11368_/Y _11370_/B vssd1 vssd1 vccd1 vccd1 _11550_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_61_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10321_ _10473_/A _10321_/B vssd1 vssd1 vccd1 vccd1 _10323_/B sky130_fd_sc_hd__nor2_1
X_13040_ hold246/X _13039_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13040_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07007__B1 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10252_ hold228/A _10252_/B vssd1 vssd1 vccd1 vccd1 _10509_/C sky130_fd_sc_hd__or2_1
XANTENNA__07558__A1 _06989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10183_ fanout58/X fanout95/X fanout54/X _10557_/A vssd1 vssd1 vccd1 vccd1 _10184_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07853__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout271 _06537_/A vssd1 vssd1 vccd1 vccd1 _12722_/A sky130_fd_sc_hd__clkbuf_8
Xfanout282 _06569_/X vssd1 vssd1 vccd1 vccd1 _06752_/A sky130_fd_sc_hd__clkbuf_8
Xfanout260 _11831_/S vssd1 vssd1 vccd1 vccd1 _12361_/B sky130_fd_sc_hd__buf_4
XANTENNA__12303__A1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout293 _13028_/A vssd1 vssd1 vccd1 vccd1 _13086_/A sky130_fd_sc_hd__buf_4
XFILLER_0_88_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10314__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12824_ hold246/X hold27/X vssd1 vssd1 vccd1 vccd1 _12825_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12755_ _11012_/A _12781_/A2 hold71/X _13166_/A vssd1 vssd1 vccd1 vccd1 hold72/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _11706_/A _11706_/B _11706_/C vssd1 vssd1 vccd1 vccd1 _11707_/B sky130_fd_sc_hd__or3_1
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12686_ reg1_val[26] _12708_/B vssd1 vssd1 vccd1 vccd1 _12687_/B sky130_fd_sc_hd__or2_1
XANTENNA__08038__A2 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11637_ _11638_/B vssd1 vssd1 vccd1 vccd1 _11637_/Y sky130_fd_sc_hd__inv_2
X_11568_ _11568_/A _11568_/B vssd1 vssd1 vccd1 vccd1 _11568_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__06932__A _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07246__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13307_ _13309_/CLK _13307_/D vssd1 vssd1 vccd1 vccd1 hold264/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10519_ _09184_/X _10507_/Y _10518_/Y _09115_/X _10517_/X vssd1 vssd1 vccd1 vccd1
+ _10519_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_25_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11499_ _11499_/A _11499_/B vssd1 vssd1 vccd1 vccd1 _11500_/B sky130_fd_sc_hd__and2_1
XFILLER_0_122_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13238_ _13305_/CLK hold223/X vssd1 vssd1 vccd1 vccd1 hold221/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11345__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ _13169_/A hold104/X vssd1 vssd1 vccd1 vccd1 _13312_/D sky130_fd_sc_hd__and2_1
XANTENNA__07763__A _07763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11285__A _11285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07730_ _08853_/A _07730_/B vssd1 vssd1 vccd1 vccd1 _07734_/A sky130_fd_sc_hd__xor2_1
XANTENNA__10305__B1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07661_ _07661_/A _07661_/B vssd1 vssd1 vccd1 vccd1 _07662_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06612_ _06610_/Y _06612_/B vssd1 vssd1 vccd1 vccd1 _06843_/A sky130_fd_sc_hd__nand2b_2
X_09400_ curr_PC[0] curr_PC[1] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09712_/B sky130_fd_sc_hd__and3_1
X_07592_ _07591_/A _07282_/B _07591_/Y vssd1 vssd1 vccd1 vccd1 _07593_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09331_ _09331_/A _09331_/B vssd1 vssd1 vccd1 vccd1 _09660_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_48_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06543_ reg1_val[16] vssd1 vssd1 vccd1 vccd1 _12641_/A sky130_fd_sc_hd__inv_2
XANTENNA__06826__B _07052_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09262_ fanout75/X fanout98/X fanout56/X _10553_/B vssd1 vssd1 vccd1 vccd1 _09263_/B
+ sky130_fd_sc_hd__o22a_1
X_08213_ _08213_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08253_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13022__A2 fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09193_ _09200_/A instruction[5] _09202_/A vssd1 vssd1 vccd1 vccd1 _09193_/X sky130_fd_sc_hd__or3_2
XFILLER_0_16_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08144_ _08144_/A _08144_/B vssd1 vssd1 vccd1 vccd1 _08203_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout226_A _07001_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12781__A1 _09252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12563__B _12563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06561__B _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08075_ _09180_/A _07168_/Y _07179_/A _08544_/C vssd1 vssd1 vccd1 vccd1 _08076_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07026_ reg1_val[9] _07026_/B vssd1 vssd1 vccd1 vccd1 _07026_/Y sky130_fd_sc_hd__xnor2_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _08978_/B _08978_/A vssd1 vssd1 vccd1 vccd1 _08977_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__10811__B _12255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07928_ _07928_/A _07928_/B vssd1 vssd1 vccd1 vccd1 _08024_/B sky130_fd_sc_hd__xor2_2
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
X_07859_ _07856_/Y _07932_/B _07854_/X vssd1 vssd1 vccd1 vccd1 _07880_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10870_ _10747_/A _10749_/X _10868_/Y _10869_/X vssd1 vssd1 vccd1 vccd1 _10872_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07712__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07712__A1 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12738__B _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09529_ _09167_/X _09171_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09529_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout41_A _12255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12540_ _12526_/B _12534_/B _12551_/A vssd1 vssd1 vccd1 vccd1 _12541_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12471_ _12471_/A _12471_/B _12471_/C vssd1 vssd1 vccd1 vccd1 _12472_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11422_ _11422_/A _11422_/B vssd1 vssd1 vccd1 vccd1 _11423_/B sky130_fd_sc_hd__or2_1
XANTENNA__07228__B1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06752__A _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11353_ _11221_/A _11221_/B _11224_/A vssd1 vssd1 vccd1 vccd1 _11358_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11284_ _11183_/B _11183_/C _11379_/A vssd1 vssd1 vccd1 vccd1 _11285_/B sky130_fd_sc_hd__a21o_1
X_10304_ _10461_/A _10304_/B vssd1 vssd1 vccd1 vccd1 _10308_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13023_ _06537_/A _13021_/Y _13022_/X _13151_/A2 hold240/X vssd1 vssd1 vccd1 vccd1
+ hold241/A sky130_fd_sc_hd__a32o_1
X_10235_ _10486_/A _10235_/B vssd1 vssd1 vccd1 vccd1 _10235_/Y sky130_fd_sc_hd__xnor2_2
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06754__A2 _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10166_ _10167_/A _10167_/B vssd1 vssd1 vccd1 vccd1 _10320_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10097_ _09812_/X _09956_/X _09957_/X vssd1 vssd1 vccd1 vccd1 _10097_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12807_ hold260/X hold25/X vssd1 vssd1 vccd1 vccd1 _13107_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__06927__A _12487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10999_ _10400_/S _10997_/X _10998_/Y _10996_/Y vssd1 vssd1 vccd1 vccd1 dest_val[13]
+ sky130_fd_sc_hd__a31o_4
XANTENNA__09456__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09456__B2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12738_ hold77/X _12788_/B vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__or2_1
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10066__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_409 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13004__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09208__A1 _09679_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12669_ _12667_/X _12669_/B vssd1 vssd1 vccd1 vccd1 _12678_/C sky130_fd_sc_hd__nand2b_2
XFILLER_0_127_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07758__A _08853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09759__A2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10184__A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08900_ _08950_/A _08900_/B vssd1 vssd1 vccd1 vccd1 _08902_/B sky130_fd_sc_hd__or2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _09881_/A _09881_/B _09879_/Y vssd1 vssd1 vccd1 vccd1 _10018_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__11318__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08831_ _08831_/A _08831_/B vssd1 vssd1 vccd1 vccd1 _08833_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08589__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10912__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08678_/A _08678_/C _08678_/B vssd1 vssd1 vccd1 vccd1 _08764_/B sky130_fd_sc_hd__a21bo_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07713_ _07974_/A _07713_/B vssd1 vssd1 vccd1 vccd1 _07716_/C sky130_fd_sc_hd__xnor2_1
X_08693_ _09622_/A _08693_/B vssd1 vssd1 vccd1 vccd1 _08696_/A sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout176_A _12781_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07644_ _08217_/B _12752_/A fanout84/X fanout55/X vssd1 vssd1 vccd1 vccd1 _07645_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09447__A1 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09447__B2 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07575_ _07576_/A _07576_/B vssd1 vssd1 vccd1 vccd1 _07575_/X sky130_fd_sc_hd__and2_1
XFILLER_0_48_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09314_ _09314_/A _09314_/B vssd1 vssd1 vccd1 vccd1 _09327_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_75_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09245_ _07506_/A _07505_/Y _07501_/Y vssd1 vssd1 vccd1 vccd1 _09247_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_106_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08670__A2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09176_ _09168_/X _09175_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09176_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08127_ _08777_/A _08127_/B vssd1 vssd1 vccd1 vccd1 _08129_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08058_ _08059_/A _08058_/B _08058_/C vssd1 vssd1 vccd1 vccd1 _08120_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_113_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11309__A2 _11308_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07009_ _07010_/A _07010_/B vssd1 vssd1 vccd1 vccd1 _07595_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_12_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08186__B2 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08186__A1 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08499__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout89_A _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10020_ _10020_/A _10020_/B vssd1 vssd1 vccd1 vccd1 _10077_/A sky130_fd_sc_hd__xor2_4
XANTENNA__06736__A2 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ _12102_/A _11971_/B vssd1 vssd1 vccd1 vccd1 _12072_/A sky130_fd_sc_hd__xnor2_2
X_10922_ fanout57/X fanout15/X fanout7/X _07553_/A vssd1 vssd1 vccd1 vccd1 _10923_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10853_ _10610_/Y _10850_/B _10852_/Y vssd1 vssd1 vccd1 vccd1 _10853_/Y sky130_fd_sc_hd__a21oi_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10784_ _12203_/A fanout52/X _10677_/B _12150_/A vssd1 vssd1 vccd1 vccd1 _10785_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11245__B2 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11245__A1 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07449__B1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12523_ _12529_/B _12523_/B vssd1 vssd1 vccd1 vccd1 new_PC[21] sky130_fd_sc_hd__xnor2_4
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08681__B _08681_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08661__A2 _07322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12745__A1 _07325_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12454_ _12614_/B _12454_/B vssd1 vssd1 vccd1 vccd1 _12455_/B sky130_fd_sc_hd__or2_1
XFILLER_0_41_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12385_ _12394_/A _12385_/B vssd1 vssd1 vccd1 vccd1 _12387_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11405_ _11378_/Y _11381_/X _11404_/X _11315_/Y vssd1 vssd1 vccd1 vccd1 dest_val[17]
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11336_ _11336_/A _11336_/B vssd1 vssd1 vccd1 vccd1 _11337_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_22_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08177__A1 _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08177__B2 _08544_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ _07005_/C _13020_/B2 hold131/X vssd1 vssd1 vccd1 vccd1 _13273_/D sky130_fd_sc_hd__o21a_1
X_11267_ _11268_/A _11268_/B vssd1 vssd1 vccd1 vccd1 _11365_/B sky130_fd_sc_hd__nand2b_1
X_11198_ hold282/A hold295/A _11198_/C vssd1 vssd1 vccd1 vccd1 _11296_/B sky130_fd_sc_hd__or3_1
X_10218_ _10218_/A _10218_/B vssd1 vssd1 vccd1 vccd1 _10220_/B sky130_fd_sc_hd__xnor2_1
X_10149_ _10149_/A _11147_/B vssd1 vssd1 vccd1 vccd1 _10150_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10287__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09429__B2 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09429__A1 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09968__A _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07360_ _12143_/A _07360_/B vssd1 vssd1 vccd1 vccd1 _07362_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12984__A1 _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09030_ _09028_/A _09028_/B _09029_/Y vssd1 vssd1 vccd1 vccd1 _09031_/B sky130_fd_sc_hd__a21o_1
X_07291_ _07356_/A _07291_/B vssd1 vssd1 vccd1 vccd1 _07293_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07488__A _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09932_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09935_/A sky130_fd_sc_hd__xor2_2
XANTENNA_fanout293_A _13028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09863_ _09738_/A _09737_/B _09735_/X vssd1 vssd1 vccd1 vccd1 _09875_/A sky130_fd_sc_hd__a21oi_4
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08814_ _08815_/A _08815_/B _08815_/C vssd1 vssd1 vccd1 vccd1 _08919_/A sky130_fd_sc_hd__a21oi_1
X_09794_ _09795_/A _09795_/B vssd1 vssd1 vccd1 vccd1 _09794_/Y sky130_fd_sc_hd__nor2_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07951__A _08853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08745_ _08744_/B _08744_/C _10015_/A vssd1 vssd1 vccd1 vccd1 _08745_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09117__A0 _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08676_ _08677_/B _08677_/C _08677_/A vssd1 vssd1 vccd1 vccd1 _08678_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07679__B1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ _07628_/A _07628_/B vssd1 vssd1 vccd1 vccd1 _07627_/X sky130_fd_sc_hd__and2b_1
X_07558_ _06989_/A _11782_/A _10433_/A vssd1 vssd1 vccd1 vccd1 _07559_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11227__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__A1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07489_ fanout81/X fanout46/X _09295_/B _11603_/A vssd1 vssd1 vccd1 vccd1 _07490_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07398__A _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09228_ _12736_/A _07389_/B fanout26/X _09772_/A vssd1 vssd1 vccd1 vccd1 _09229_/B
+ sky130_fd_sc_hd__o22a_1
X_09159_ _09157_/X _09158_/X _09359_/S vssd1 vssd1 vccd1 vccd1 _09159_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12170_ _06852_/X _12169_/X _12322_/S vssd1 vssd1 vccd1 vccd1 _12170_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10202__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11121_ _11121_/A _11121_/B vssd1 vssd1 vccd1 vccd1 _11131_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11052_ _11052_/A _11052_/B vssd1 vssd1 vccd1 vccd1 _11054_/C sky130_fd_sc_hd__xor2_1
X_10003_ _10617_/A _10003_/B vssd1 vssd1 vccd1 vccd1 _10003_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11954_ _11955_/A _11955_/B _11955_/C vssd1 vssd1 vccd1 vccd1 _12032_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11885_ _11886_/B _11886_/A vssd1 vssd1 vccd1 vccd1 _11964_/B sky130_fd_sc_hd__nand2b_1
X_10905_ fanout35/X _11431_/A fanout70/X fanout37/X vssd1 vssd1 vccd1 vccd1 _10906_/B
+ sky130_fd_sc_hd__o22a_1
X_10836_ _10837_/A _10837_/B vssd1 vssd1 vccd1 vccd1 _10953_/A sky130_fd_sc_hd__or2_1
XANTENNA__12966__A1 _07115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11769__A2 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08095__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10767_ _09184_/X _10752_/X _10754_/X _06918_/X _10766_/X vssd1 vssd1 vccd1 vccd1
+ _10767_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_124_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12506_ _12551_/A _12507_/B vssd1 vssd1 vccd1 vccd1 _12516_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_89_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10698_ _10698_/A _10698_/B vssd1 vssd1 vccd1 vccd1 _10699_/C sky130_fd_sc_hd__or2_1
X_12437_ _12443_/B _12437_/B vssd1 vssd1 vccd1 vccd1 new_PC[8] sky130_fd_sc_hd__and2_4
XANTENNA__07101__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12368_ hold103/A _12368_/B vssd1 vssd1 vccd1 vccd1 _12368_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12299_ _12345_/A _12299_/B vssd1 vssd1 vccd1 vccd1 dest_val[29] sky130_fd_sc_hd__nor2_8
XFILLER_0_38_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11319_ _11695_/A _11319_/B vssd1 vssd1 vccd1 vccd1 _11321_/B sky130_fd_sc_hd__xnor2_1
X_06860_ _09200_/A _06859_/Y _06849_/X vssd1 vssd1 vccd1 vccd1 _06860_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07373__A2 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10901__B1 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06791_ reg1_val[3] _06964_/A vssd1 vssd1 vccd1 vccd1 _06791_/Y sky130_fd_sc_hd__nand2_1
X_08530_ _08521_/A _08520_/C _08520_/B vssd1 vssd1 vccd1 vccd1 _08531_/C sky130_fd_sc_hd__a21o_1
X_08461_ _08461_/A _08461_/B vssd1 vssd1 vccd1 vccd1 _08482_/B sky130_fd_sc_hd__xnor2_2
X_07412_ _08897_/A _07412_/B vssd1 vssd1 vccd1 vccd1 _07625_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_58_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08392_ _08589_/A _08392_/B vssd1 vssd1 vccd1 vccd1 _08421_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10680__A2 _07322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12957__B2 _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10968__B1 _09059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07343_ _10565_/A _07343_/B vssd1 vssd1 vccd1 vccd1 _07344_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout139_A _07004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11090__C1 _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07274_ _07274_/A _07274_/B vssd1 vssd1 vccd1 vccd1 _07295_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09013_ _09010_/Y _09050_/A _08503_/Y vssd1 vssd1 vccd1 vccd1 _09054_/B sky130_fd_sc_hd__o21a_1
Xhold110 hold110/A vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold121 hold121/A vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold132 hold161/X vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 hold143/A vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11393__B1 _12487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold176 hold186/X vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__buf_1
Xhold154 hold154/A vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13159__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11468__A _11468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 hold187/A vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _10006_/A _09915_/B _09900_/Y vssd1 vssd1 vccd1 vccd1 _10006_/B sky130_fd_sc_hd__nor3b_2
XFILLER_0_0_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09846_ _09683_/X _09684_/Y _09686_/B vssd1 vssd1 vccd1 vccd1 _09850_/A sky130_fd_sc_hd__o21a_1
XANTENNA__11696__A1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12893__B1 fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08777__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11696__B2 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06989_ _06989_/A _11782_/A vssd1 vssd1 vccd1 vccd1 _06989_/X sky130_fd_sc_hd__and2_1
XANTENNA__12299__A _12345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09777_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09778_/B sky130_fd_sc_hd__xnor2_2
X_08728_ _08728_/A _08728_/B vssd1 vssd1 vccd1 vccd1 _08731_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _08841_/A1 _08134_/B fanout51/X _08841_/B2 vssd1 vssd1 vccd1 vccd1 _08660_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12746__B _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11670_ _07068_/A _12250_/B _06930_/Y _11669_/X vssd1 vssd1 vccd1 vccd1 _11670_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10671__A2 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08077__B1 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10621_ _10621_/A _10621_/B vssd1 vssd1 vccd1 vccd1 _10621_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10552_ _10552_/A _10552_/B vssd1 vssd1 vccd1 vccd1 _10570_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_91_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13271_ _13277_/CLK _13271_/D vssd1 vssd1 vccd1 vccd1 hold126/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12762__A _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12222_ _11973_/B _12221_/X _11973_/A vssd1 vssd1 vccd1 vccd1 _12222_/X sky130_fd_sc_hd__a21o_1
X_10483_ _10485_/A _10485_/B vssd1 vssd1 vccd1 vccd1 _10483_/X sky130_fd_sc_hd__or2_1
XANTENNA__11384__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13069__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12153_ _12154_/A _12154_/B vssd1 vssd1 vccd1 vccd1 _12213_/A sky130_fd_sc_hd__and2b_1
X_11104_ _12373_/A1 _11391_/B _11102_/X vssd1 vssd1 vccd1 vccd1 _11104_/Y sky130_fd_sc_hd__a21oi_1
X_12084_ _12085_/B _12085_/A vssd1 vssd1 vccd1 vccd1 _12084_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_20_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11136__B1 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11035_ _11121_/A _11035_/B vssd1 vssd1 vccd1 vccd1 _11044_/A sky130_fd_sc_hd__nor2_1
X_12986_ _07194_/C _12744_/B hold99/X vssd1 vssd1 vccd1 vccd1 _13263_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_91_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11937_ _11938_/A _11938_/B _11938_/C vssd1 vssd1 vccd1 vccd1 _11939_/A sky130_fd_sc_hd__o21ai_1
X_11868_ _12772_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _11872_/A sky130_fd_sc_hd__or2_1
XFILLER_0_55_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10819_ _10819_/A _10819_/B vssd1 vssd1 vccd1 vccd1 _10925_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11799_ _11800_/A _11800_/B vssd1 vssd1 vccd1 vccd1 _11849_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06670__A _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07961_ _07034_/Y _08772_/B2 _08772_/A2 _09925_/A1 vssd1 vssd1 vccd1 vccd1 _07962_/B
+ sky130_fd_sc_hd__o22a_1
X_06912_ instruction[21] _06552_/X _06911_/X _06678_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[3]
+ sky130_fd_sc_hd__o211a_4
X_09700_ hold237/A _09698_/X _09699_/Y vssd1 vssd1 vccd1 vccd1 _09707_/C sky130_fd_sc_hd__o21a_1
XANTENNA__11127__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07892_ _07892_/A _07892_/B vssd1 vssd1 vccd1 vccd1 _07897_/A sky130_fd_sc_hd__or2_1
XFILLER_0_65_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06843_ _06843_/A _06843_/B vssd1 vssd1 vccd1 vccd1 _06843_/Y sky130_fd_sc_hd__nand2_1
X_09631_ _11125_/A _09631_/B vssd1 vssd1 vccd1 vccd1 _09632_/B sky130_fd_sc_hd__xnor2_2
X_06774_ _06783_/A _06649_/A _12573_/B _06772_/X vssd1 vssd1 vccd1 vccd1 _07279_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__09205__B _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09562_ _09498_/A _09498_/B _09499_/Y vssd1 vssd1 vccd1 vccd1 _09656_/A sky130_fd_sc_hd__o21ai_4
X_08513_ _09620_/A _08513_/B vssd1 vssd1 vccd1 vccd1 _08540_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_fanout256_A _12487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09493_ _09310_/A _09310_/B _09308_/Y vssd1 vssd1 vccd1 vccd1 _09495_/B sky130_fd_sc_hd__a21boi_4
X_08444_ _08445_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08444_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10653__A2 _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11850__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11850__B2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08375_ _08375_/A _08375_/B vssd1 vssd1 vccd1 vccd1 _08430_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_18_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07326_ fanout46/X _09295_/B _11603_/A _10433_/A vssd1 vssd1 vccd1 vccd1 _07327_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07257_ reg1_val[16] _07257_/B vssd1 vssd1 vccd1 vccd1 _07259_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_14_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07188_ reg1_val[15] _07188_/B vssd1 vssd1 vccd1 vccd1 _07894_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_112_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout71_A _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ _10752_/S _09828_/Y _09214_/A vssd1 vssd1 vccd1 vccd1 _12181_/B sky130_fd_sc_hd__a21boi_1
X_12840_ _13047_/A _13048_/A _13047_/B vssd1 vssd1 vccd1 vccd1 _13053_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_68_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12771_ _11793_/A _12781_/A2 hold87/X _13147_/A vssd1 vssd1 vccd1 vccd1 _13207_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08837__A2 _07322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11722_/A _11722_/B _11722_/C vssd1 vssd1 vccd1 vccd1 _11723_/B sky130_fd_sc_hd__nor3_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ _11568_/A _11568_/B _11566_/A vssd1 vssd1 vccd1 vccd1 _11654_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout82 _07312_/X vssd1 vssd1 vccd1 vccd1 fanout82/X sky130_fd_sc_hd__buf_4
XFILLER_0_92_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout71 _12766_/A vssd1 vssd1 vccd1 vccd1 _11688_/A sky130_fd_sc_hd__buf_6
Xfanout60 _07153_/X vssd1 vssd1 vccd1 vccd1 _12150_/B sky130_fd_sc_hd__clkbuf_8
X_10604_ _10606_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _10604_/X sky130_fd_sc_hd__or2_1
XFILLER_0_119_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ instruction[15] vssd1 vssd1 vccd1 vccd1 loadstore_dest[4] sky130_fd_sc_hd__buf_12
X_11584_ curr_PC[19] _11671_/C _12005_/A vssd1 vssd1 vccd1 vccd1 _11584_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout93 fanout94/X vssd1 vssd1 vccd1 vccd1 _07553_/A sky130_fd_sc_hd__buf_6
XANTENNA__09262__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10535_ _12255_/A _10535_/B vssd1 vssd1 vccd1 vccd1 _10539_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13254_ _13289_/CLK hold148/X vssd1 vssd1 vccd1 vccd1 hold146/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10466_ _10466_/A _10466_/B _10466_/C vssd1 vssd1 vccd1 vccd1 _10468_/A sky130_fd_sc_hd__and3_1
XFILLER_0_122_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08222__B1 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13185_ _13280_/CLK hold37/X vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dfxtp_1
X_12205_ _12205_/A fanout8/X vssd1 vssd1 vccd1 vccd1 _12206_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12136_ curr_PC[26] _12136_/B vssd1 vssd1 vccd1 vccd1 _12139_/B sky130_fd_sc_hd__nand2_1
X_10397_ curr_PC[7] curr_PC[8] _10397_/C vssd1 vssd1 vccd1 vccd1 _10646_/C sky130_fd_sc_hd__and3_1
XFILLER_0_20_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06784__B1 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11109__B1 _11106_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12067_ _09205_/B _12055_/X _12066_/X _12048_/X vssd1 vssd1 vccd1 vccd1 _12067_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10740__A _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09722__B1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ _11158_/B _11018_/B vssd1 vssd1 vccd1 vccd1 _11046_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__06649__B _12583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12969_ hold146/X _12723_/A _13170_/B hold121/X _13066_/A vssd1 vssd1 vccd1 vccd1
+ hold153/A sky130_fd_sc_hd__o221a_1
XFILLER_0_75_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08160_ _08160_/A _08160_/B vssd1 vssd1 vccd1 vccd1 _08209_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_117_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07111_ _07119_/A _07111_/B _07111_/C vssd1 vssd1 vccd1 vccd1 _07128_/C sky130_fd_sc_hd__and3_1
XFILLER_0_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11596__B1 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08091_ _08091_/A _08151_/A vssd1 vssd1 vccd1 vccd1 _08103_/B sky130_fd_sc_hd__and2_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07042_ reg1_val[4] reg1_val[5] _07105_/B _07105_/A vssd1 vssd1 vccd1 vccd1 _07043_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08993_ _08995_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _09509_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_11_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07944_ _07726_/A _07725_/Y _07721_/Y vssd1 vssd1 vccd1 vccd1 _07948_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__11746__A _11746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07875_ _07872_/B _07872_/C _07872_/A vssd1 vssd1 vccd1 vccd1 _07876_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__06559__B _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_2_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06826_ reg1_val[21] _07052_/B vssd1 vssd1 vccd1 vccd1 _06826_/Y sky130_fd_sc_hd__nand2_1
X_09614_ _10458_/A _09614_/B vssd1 vssd1 vccd1 vccd1 _09616_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08819__A2 _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06757_ reg1_val[5] _06972_/C vssd1 vssd1 vccd1 vccd1 _06758_/B sky130_fd_sc_hd__nand2_1
X_09545_ _06788_/X _09544_/Y _12322_/S vssd1 vssd1 vccd1 vccd1 _09545_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12076__A1 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12076__B2 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06688_ reg2_val[16] _06752_/A _06688_/B1 _06687_/Y vssd1 vssd1 vccd1 vccd1 _07167_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_09476_ _09476_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _09482_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08427_ _08427_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08456_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08358_ _08358_/A _08358_/B _08358_/C vssd1 vssd1 vccd1 vccd1 _08390_/A sky130_fd_sc_hd__or3_2
XFILLER_0_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08289_ _08287_/A _08287_/B _08343_/A vssd1 vssd1 vccd1 vccd1 _08299_/A sky130_fd_sc_hd__a21bo_2
X_07309_ _07175_/A _07175_/B _07175_/C _07303_/B vssd1 vssd1 vccd1 vccd1 _07319_/B
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_73_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ _10320_/A _10320_/B _10320_/C vssd1 vssd1 vccd1 vccd1 _10321_/B sky130_fd_sc_hd__and3_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10251_ _10248_/X _10250_/X _10251_/S vssd1 vssd1 vccd1 vccd1 _10251_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07007__A1 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07007__B2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07558__A2 _11782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ _10182_/A _10182_/B vssd1 vssd1 vccd1 vccd1 _10185_/A sky130_fd_sc_hd__xnor2_1
Xfanout272 hold152/X vssd1 vssd1 vccd1 vccd1 _06537_/A sky130_fd_sc_hd__clkbuf_4
Xfanout261 _12284_/A vssd1 vssd1 vccd1 vccd1 _11831_/S sky130_fd_sc_hd__clkbuf_4
Xfanout283 _06898_/A vssd1 vssd1 vccd1 vccd1 _06783_/A sky130_fd_sc_hd__buf_6
Xfanout294 _13028_/A vssd1 vssd1 vccd1 vccd1 _13066_/A sky130_fd_sc_hd__buf_4
XANTENNA__10314__A1 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10314__B2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ hold27/X hold246/X vssd1 vssd1 vccd1 vccd1 _12823_/X sky130_fd_sc_hd__and2b_1
XANTENNA__12067__A1 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12754_ hold70/X _12786_/B vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__or2_1
XFILLER_0_96_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _11706_/A _11706_/B _11706_/C vssd1 vssd1 vccd1 vccd1 _11797_/A sky130_fd_sc_hd__o21a_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12685_ reg1_val[26] _12708_/B vssd1 vssd1 vccd1 vccd1 _12685_/X sky130_fd_sc_hd__and2_1
XFILLER_0_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11636_ _11636_/A _11814_/A vssd1 vssd1 vccd1 vccd1 _11638_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11567_ _11476_/B _11478_/B _11476_/A vssd1 vssd1 vccd1 vccd1 _11568_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__07246__A1 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07246__B2 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_331 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13111__A _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13306_ _13306_/CLK _13306_/D vssd1 vssd1 vccd1 vccd1 hold286/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10518_ _10251_/S _10116_/X _09214_/A vssd1 vssd1 vccd1 vccd1 _10518_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__06932__B _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13237_ _13305_/CLK hold236/X vssd1 vssd1 vccd1 vccd1 hold234/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11498_ _11499_/A _11499_/B vssd1 vssd1 vccd1 vccd1 _11618_/A sky130_fd_sc_hd__nor2_1
X_10449_ _10464_/A vssd1 vssd1 vccd1 vccd1 _10592_/B sky130_fd_sc_hd__inv_2
X_13168_ hold287/X _13168_/A2 _13167_/X _13168_/B1 hold103/X vssd1 vssd1 vccd1 vccd1
+ hold104/A sky130_fd_sc_hd__a32o_1
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13099_ hold258/X _13098_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13099_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11750__B1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ hold286/A _12183_/C _12119_/B1 vssd1 vssd1 vccd1 vccd1 _12119_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_46_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10305__B2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10305__A1 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ _07661_/A _07661_/B vssd1 vssd1 vccd1 vccd1 _07687_/B sky130_fd_sc_hd__and2_1
XANTENNA__12397__A _12573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06611_ reg1_val[27] _07434_/A vssd1 vssd1 vccd1 vccd1 _06612_/B sky130_fd_sc_hd__nand2_2
X_07591_ _07591_/A _09775_/A vssd1 vssd1 vccd1 vccd1 _07591_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06542_ reg1_val[8] vssd1 vssd1 vccd1 vccd1 _06542_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ _09331_/A _09331_/B vssd1 vssd1 vccd1 vccd1 _09330_/X sky130_fd_sc_hd__and2_1
XFILLER_0_62_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09261_ _09261_/A _09261_/B vssd1 vssd1 vccd1 vccd1 _09282_/A sky130_fd_sc_hd__xnor2_2
X_08212_ _08212_/A _08212_/B vssd1 vssd1 vccd1 vccd1 _08253_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08682__B1 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09192_ _09200_/A instruction[5] _09202_/A vssd1 vssd1 vccd1 vccd1 _09192_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_126_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08143_ _08853_/A _08143_/B vssd1 vssd1 vccd1 vccd1 _08203_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08074_ _08080_/A _08080_/B vssd1 vssd1 vccd1 vccd1 _08074_/X sky130_fd_sc_hd__and2_1
XANTENNA__12781__A2 _12781_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07025_ reg1_val[7] reg1_val[8] _07038_/B _07105_/A vssd1 vssd1 vccd1 vccd1 _07026_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__buf_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _08978_/A _08978_/B vssd1 vssd1 vccd1 vccd1 _08976_/X sky130_fd_sc_hd__and2b_1
X_07927_ _08056_/A _08056_/B _07923_/Y vssd1 vssd1 vccd1 vccd1 _08024_/A sky130_fd_sc_hd__a21boi_2
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
X_07858_ _09580_/A _07858_/B vssd1 vssd1 vccd1 vccd1 _07932_/B sky130_fd_sc_hd__xnor2_2
X_07789_ _07789_/A _07789_/B vssd1 vssd1 vccd1 vccd1 _07790_/C sky130_fd_sc_hd__or2_1
X_06809_ _07303_/A reg1_val[12] vssd1 vssd1 vccd1 vccd1 _06809_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07712__A2 _07322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09528_ _09392_/X _09527_/X _10249_/S vssd1 vssd1 vccd1 vccd1 _09528_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08673__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09459_ _10578_/A _09459_/B vssd1 vssd1 vccd1 vccd1 _09461_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12470_ _12471_/A _12471_/B _12471_/C vssd1 vssd1 vccd1 vccd1 _12478_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11421_ _11422_/A _11422_/B vssd1 vssd1 vccd1 vccd1 _11532_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07228__B2 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07228__A1 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11352_ _11257_/A _11257_/B _11255_/Y vssd1 vssd1 vccd1 vccd1 _11362_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_22_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10555__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10303_ _10303_/A _10303_/B vssd1 vssd1 vccd1 vccd1 _10304_/B sky130_fd_sc_hd__and2_1
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11283_ _11216_/X _11316_/B _11282_/Y vssd1 vssd1 vccd1 vccd1 _11283_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07864__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13022_ hold36/X fanout1/X hold38/X vssd1 vssd1 vccd1 vccd1 _13022_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09925__B1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10234_ _09664_/B _10230_/C _10233_/Y vssd1 vssd1 vccd1 vccd1 _10235_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11732__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10165_ _10306_/A _10165_/B vssd1 vssd1 vccd1 vccd1 _10167_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09689__C1 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ _10229_/B _10229_/C vssd1 vssd1 vccd1 vccd1 _10096_/X sky130_fd_sc_hd__or2_1
XANTENNA__08695__A _08695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13106__A _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12806_ hold25/X hold260/X vssd1 vssd1 vccd1 vccd1 _12806_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_57_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10998_ curr_PC[13] _11107_/C vssd1 vssd1 vccd1 vccd1 _10998_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09456__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12737_ hold13/X _12788_/B _12736_/Y _13086_/A vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__o211a_1
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12668_ reg1_val[22] _12714_/A vssd1 vssd1 vccd1 vccd1 _12669_/B sky130_fd_sc_hd__or2_1
XFILLER_0_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11619_ _11619_/A _11619_/B vssd1 vssd1 vccd1 vccd1 _11620_/B sky130_fd_sc_hd__and2_1
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12599_ _12597_/Y _12599_/B vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07774__A _08415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08830_ _08848_/A vssd1 vssd1 vccd1 vccd1 _08830_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _08761_/A _08761_/B vssd1 vssd1 vccd1 vccd1 _08764_/A sky130_fd_sc_hd__xnor2_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07712_ _08748_/B1 _07322_/A _07322_/B _12730_/A fanout46/X vssd1 vssd1 vccd1 vccd1
+ _07713_/B sky130_fd_sc_hd__o32a_1
X_08692_ _11794_/A _08692_/A2 _08692_/B1 _12768_/A vssd1 vssd1 vccd1 vccd1 _08693_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07643_ _08232_/A _07643_/B vssd1 vssd1 vccd1 vccd1 _07648_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07574_ _07585_/A _07585_/B _07570_/X vssd1 vssd1 vccd1 vccd1 _07576_/B sky130_fd_sc_hd__a21o_1
X_09313_ _09311_/Y _09313_/B vssd1 vssd1 vccd1 vccd1 _09314_/B sky130_fd_sc_hd__and2b_1
XANTENNA__09447__A2 _07132_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10057__A3 _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07014__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09244_ _07563_/B _07566_/B _07561_/X vssd1 vssd1 vccd1 vccd1 _09247_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__12739__C1 _13028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09175_ _09171_/X _09174_/X _09676_/S vssd1 vssd1 vccd1 vccd1 _09175_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08126_ _08841_/A1 _08477_/B _08776_/B1 _08841_/B2 vssd1 vssd1 vccd1 vccd1 _08127_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08057_ _08055_/A _08055_/C _08055_/B vssd1 vssd1 vccd1 vccd1 _08058_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_113_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06984__A3 _07001_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09907__B1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07008_ _10306_/A _07008_/B vssd1 vssd1 vccd1 vccd1 _07010_/B sky130_fd_sc_hd__xor2_1
XANTENNA__08186__A2 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10822__B _10925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06736__A3 _12603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07394__B1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ _08959_/A _08959_/B vssd1 vssd1 vccd1 vccd1 _08960_/B sky130_fd_sc_hd__xor2_4
X_11970_ _12216_/A _12216_/B _11968_/Y vssd1 vssd1 vccd1 vccd1 _11971_/B sky130_fd_sc_hd__o21ba_1
X_10921_ _10921_/A _10921_/B vssd1 vssd1 vccd1 vccd1 _10930_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10852_ _10604_/X _10726_/Y _10727_/X vssd1 vssd1 vccd1 vccd1 _10852_/Y sky130_fd_sc_hd__a21oi_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10783_ _10783_/A _10783_/B vssd1 vssd1 vccd1 vccd1 _10795_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11245__A2 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07449__A1 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07449__B2 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12522_ _12529_/A _12518_/Y _12514_/A vssd1 vssd1 vccd1 vccd1 _12523_/B sky130_fd_sc_hd__o21ai_2
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08661__A3 _07322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12453_ _12614_/B _12454_/B vssd1 vssd1 vccd1 vccd1 _12464_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12745__A2 _12980_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11404_ _11404_/A _11404_/B _11404_/C _11404_/D vssd1 vssd1 vccd1 vccd1 _11404_/X
+ sky130_fd_sc_hd__or4_2
X_12384_ _12563_/B _12384_/B vssd1 vssd1 vccd1 vccd1 _12385_/B sky130_fd_sc_hd__or2_1
XFILLER_0_34_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11335_ _11336_/A _11336_/B vssd1 vssd1 vccd1 vccd1 _11337_/A sky130_fd_sc_hd__and2_1
XFILLER_0_104_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11266_ _11266_/A _11266_/B vssd1 vssd1 vccd1 vccd1 _11268_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08177__A2 _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13005_ hold100/X _13013_/A2 _13020_/A2 hold130/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold131/A sky130_fd_sc_hd__o221a_1
X_10217_ _10085_/A _10085_/B _10083_/Y vssd1 vssd1 vccd1 vccd1 _10218_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11197_ _11193_/Y _11196_/Y _11197_/S vssd1 vssd1 vccd1 vccd1 _11197_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12005__A _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ _10148_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _10150_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10079_ _09948_/A _09948_/B _09946_/Y vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09429__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07769__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07290_ _07291_/B _07356_/A vssd1 vssd1 vccd1 vccd1 _07601_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09601__A2 _09472_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11944__B1 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10923__A _12255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09931_ _10559_/A _09931_/B vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09862_ _09881_/B _09749_/B _09771_/B _09769_/Y vssd1 vssd1 vccd1 vccd1 _09876_/A
+ sky130_fd_sc_hd__o31ai_4
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _08813_/A _08813_/B vssd1 vssd1 vccd1 vccd1 _08815_/C sky130_fd_sc_hd__or2_1
X_09793_ _09793_/A _09793_/B vssd1 vssd1 vccd1 vccd1 _09795_/B sky130_fd_sc_hd__xnor2_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ _10015_/A _08744_/B _08744_/C vssd1 vssd1 vccd1 vccd1 _08744_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _08674_/B _08674_/C _08857_/A vssd1 vssd1 vccd1 vccd1 _08677_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__07679__A1 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07679__B2 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06567__B _06567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07626_ _07626_/A _07626_/B vssd1 vssd1 vccd1 vccd1 _07628_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_76_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07557_ _09294_/A _10551_/A vssd1 vssd1 vccd1 vccd1 _07559_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11227__A2 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07488_ _10559_/A _07488_/B vssd1 vssd1 vccd1 vccd1 _07589_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12188__B1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09227_ _09243_/B _07517_/B _07526_/B _07527_/B _07527_/A vssd1 vssd1 vccd1 vccd1
+ _09240_/B sky130_fd_sc_hd__a32o_1
XANTENNA__06643__A2_N _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09158_ reg1_val[31] _09180_/A _09158_/S vssd1 vssd1 vccd1 vccd1 _09158_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09894__A _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08109_ _08109_/A _08109_/B vssd1 vssd1 vccd1 vccd1 _08165_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09089_ _09088_/A _09088_/B _09079_/A _09079_/B _09082_/X vssd1 vssd1 vccd1 vccd1
+ _12230_/B sky130_fd_sc_hd__a2111o_1
XFILLER_0_101_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11120_ _11121_/A _11121_/B vssd1 vssd1 vccd1 vccd1 _11262_/A sky130_fd_sc_hd__and2_1
XFILLER_0_102_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11051_ _10928_/A _10928_/B _10926_/A vssd1 vssd1 vccd1 vccd1 _11052_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__09833__S _10249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ _10002_/A _10002_/B _10002_/C vssd1 vssd1 vccd1 vccd1 _10003_/B sky130_fd_sc_hd__and3_1
XFILLER_0_99_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11953_ _12032_/A _11953_/B vssd1 vssd1 vccd1 vccd1 _11955_/C sky130_fd_sc_hd__and2_1
X_11884_ _11964_/A _11884_/B vssd1 vssd1 vccd1 vccd1 _11886_/B sky130_fd_sc_hd__nand2_1
X_10904_ _10904_/A _10904_/B vssd1 vssd1 vccd1 vccd1 _10908_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_67_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10835_ _10719_/A _10719_/B _10717_/X vssd1 vssd1 vccd1 vccd1 _10837_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12966__A2 _12742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08095__A1 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10426__B1 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08095__B2 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10766_ _10756_/Y _10757_/X _10765_/Y _09115_/X _10764_/X vssd1 vssd1 vccd1 vccd1
+ _10766_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_66_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12505_ reg1_val[19] curr_PC[19] _12524_/S vssd1 vssd1 vccd1 vccd1 _12507_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_82_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10697_ _10698_/A _10698_/B vssd1 vssd1 vccd1 vccd1 _10832_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_124_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12436_ _12436_/A _12436_/B _12436_/C vssd1 vssd1 vccd1 vccd1 _12437_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12367_ hold287/A _12337_/X _09842_/B vssd1 vssd1 vccd1 vccd1 _12368_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12298_ _07243_/A _12250_/B _06930_/Y _12297_/X vssd1 vssd1 vccd1 vccd1 _12299_/B
+ sky130_fd_sc_hd__o22a_2
X_11318_ fanout19/X fanout47/X _11603_/A _12203_/A vssd1 vssd1 vccd1 vccd1 _11319_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11249_ _11250_/A _11250_/B vssd1 vssd1 vccd1 vccd1 _11327_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10901__A1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10901__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06790_ _06870_/A _06788_/X _06789_/X vssd1 vssd1 vccd1 vccd1 _06790_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12249__A4 _12248_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_7_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08460_ _08488_/A _08460_/B vssd1 vssd1 vccd1 vccd1 _08482_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10665__B1 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08391_ _08841_/A1 _08588_/B _09273_/A1 _08841_/B2 vssd1 vssd1 vccd1 vccd1 _08392_/B
+ sky130_fd_sc_hd__o22a_1
X_07411_ _07411_/A _07411_/B vssd1 vssd1 vccd1 vccd1 _07625_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07530__B1 _12713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07342_ _10144_/B2 _11603_/A _10433_/A fanout46/X vssd1 vssd1 vccd1 vccd1 _07343_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10680__A3 _07322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10968__A1 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07273_ _07274_/B vssd1 vssd1 vccd1 vccd1 _07273_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_116_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09012_ _09049_/A _09049_/B _09049_/C vssd1 vssd1 vccd1 vccd1 _09050_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_60_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold100 hold100/A vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold122 hold122/A vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 hold144/A vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 hold133/A vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold111 hold111/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold177 hold177/A vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 hold166/A vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12254__B1_N _12255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold199 hold199/A vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 hold188/A vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _10037_/B _09913_/C _09913_/A vssd1 vssd1 vccd1 vccd1 _09915_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07962__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09845_ _10752_/S _11923_/A2 _12243_/B1 _06764_/B _09844_/X vssd1 vssd1 vccd1 vccd1
+ _09845_/X sky130_fd_sc_hd__o221a_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12893__B2 _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11696__A2 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _09777_/A _09777_/B vssd1 vssd1 vccd1 vccd1 _09776_/X sky130_fd_sc_hd__and2b_1
X_06988_ _10555_/A _11695_/A _06987_/B vssd1 vssd1 vccd1 vccd1 _11782_/A sky130_fd_sc_hd__or3b_4
X_08727_ _08728_/A _08728_/B vssd1 vssd1 vccd1 vccd1 _08727_/Y sky130_fd_sc_hd__nand2_1
X_08658_ _08658_/A _08658_/B vssd1 vssd1 vccd1 vccd1 _08703_/A sky130_fd_sc_hd__xnor2_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10656__B1 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09889__A _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_8_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13280_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07609_ _07593_/A _07593_/B _07596_/A vssd1 vssd1 vccd1 vccd1 _07611_/B sky130_fd_sc_hd__a21oi_4
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _08589_/A _08598_/S vssd1 vssd1 vccd1 vccd1 _08591_/B sky130_fd_sc_hd__xor2_1
XANTENNA__13070__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08077__B2 _08692_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08077__A1 _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10620_ _06804_/X _10619_/X _11738_/S vssd1 vssd1 vccd1 vccd1 _10621_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_64_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06582__A2_N _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07202__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10551_ _10551_/A _10551_/B vssd1 vssd1 vccd1 vccd1 _10552_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_107_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13270_ _13277_/CLK hold109/X vssd1 vssd1 vccd1 vccd1 hold107/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10482_ _10482_/A _10482_/B vssd1 vssd1 vccd1 vccd1 _10485_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_122_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12221_ _12221_/A _12221_/B _12221_/C vssd1 vssd1 vccd1 vccd1 _12221_/X sky130_fd_sc_hd__and3_1
XFILLER_0_44_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12152_ _12152_/A _12152_/B vssd1 vssd1 vccd1 vccd1 _12154_/B sky130_fd_sc_hd__xor2_1
X_11103_ _11195_/A _09369_/X _09214_/A vssd1 vssd1 vccd1 vccd1 _11391_/B sky130_fd_sc_hd__o21a_1
X_12083_ _12083_/A _12083_/B vssd1 vssd1 vccd1 vccd1 _12085_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12333__B1 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11136__A1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11136__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11034_ _11034_/A _11034_/B vssd1 vssd1 vccd1 vccd1 _11035_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07591__B _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10895__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12985_ hold98/X _13013_/A2 _13170_/B hold90/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold99/A sky130_fd_sc_hd__o221a_1
X_11936_ _12011_/A _11936_/B vssd1 vssd1 vccd1 vccd1 _11938_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11867_ _12200_/A _11867_/B vssd1 vssd1 vccd1 vccd1 _11875_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10818_ fanout54/X fanout20/X fanout18/X fanout95/X vssd1 vssd1 vccd1 vccd1 _10819_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10457__B _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11798_ _11849_/A _11798_/B vssd1 vssd1 vccd1 vccd1 _11800_/B sky130_fd_sc_hd__and2_1
XFILLER_0_125_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10749_ _10753_/A _10753_/B vssd1 vssd1 vccd1 vccd1 _10749_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_55_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06951__A _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12419_ _12588_/B _12419_/B vssd1 vssd1 vccd1 vccd1 _12420_/B sky130_fd_sc_hd__or2_1
XANTENNA__06670__B _12573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07960_ _08232_/A _07960_/B vssd1 vssd1 vccd1 vccd1 _07964_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06911_ instruction[28] _06915_/B vssd1 vssd1 vccd1 vccd1 _06911_/X sky130_fd_sc_hd__or2_1
XANTENNA__11127__B2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11127__A1 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07891_ _08855_/A _07891_/B vssd1 vssd1 vccd1 vccd1 _07892_/B sky130_fd_sc_hd__and2_1
XANTENNA__10886__B1 _12345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06842_ _06620_/B _06841_/X _06838_/Y vssd1 vssd1 vccd1 vccd1 _06843_/B sky130_fd_sc_hd__a21o_1
X_09630_ fanout75/X _08217_/B fanout55/X _10553_/B vssd1 vssd1 vccd1 vccd1 _09631_/B
+ sky130_fd_sc_hd__o22a_1
X_06773_ _06783_/A _06649_/A _12573_/B _06772_/X vssd1 vssd1 vccd1 vccd1 _10249_/S
+ sky130_fd_sc_hd__a31oi_4
X_09561_ _09503_/A _09503_/B _09501_/X vssd1 vssd1 vccd1 vccd1 _09659_/A sky130_fd_sc_hd__a21oi_4
X_08512_ _06864_/A _09888_/B2 _12736_/A _08758_/A2 vssd1 vssd1 vccd1 vccd1 _08513_/B
+ sky130_fd_sc_hd__o22a_1
X_09492_ _09292_/A _09292_/B _09290_/X vssd1 vssd1 vccd1 vccd1 _09495_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__07503__B1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08443_ _08443_/A _08443_/B vssd1 vssd1 vccd1 vccd1 _08473_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_81_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout151_A _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout249_A _08695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10648__A _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11850__A2 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08374_ _08375_/A _08375_/B vssd1 vssd1 vccd1 vccd1 _08620_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13024__A _13028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07325_ _07325_/A _07325_/B vssd1 vssd1 vccd1 vccd1 _07325_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__07957__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ _08836_/A vssd1 vssd1 vccd1 vccd1 _10578_/A sky130_fd_sc_hd__inv_4
XFILLER_0_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12582__B _12583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06580__B _06633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07187_ reg1_val[15] _07188_/B vssd1 vssd1 vccd1 vccd1 _10819_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_5_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08231__A1 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08231__B2 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09828_ _10750_/S _09677_/X _11195_/C vssd1 vssd1 vccd1 vccd1 _09828_/Y sky130_fd_sc_hd__o21ai_1
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09759_ _10553_/B _08134_/B fanout51/X fanout69/X vssd1 vssd1 vccd1 vccd1 _09760_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout64_A _12774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12770_ hold86/X _12778_/B vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__or2_1
XFILLER_0_96_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08837__A3 _07322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06848__A2 _06622_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11721_ _11721_/A vssd1 vssd1 vccd1 vccd1 _11723_/A sky130_fd_sc_hd__inv_2
XFILLER_0_126_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08028__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11652_/A _11652_/B vssd1 vssd1 vccd1 vccd1 _11654_/A sky130_fd_sc_hd__nand2_1
Xfanout83 _07305_/Y vssd1 vssd1 vccd1 vccd1 fanout83/X sky130_fd_sc_hd__buf_8
Xfanout61 _07153_/X vssd1 vssd1 vccd1 vccd1 _10677_/A sky130_fd_sc_hd__clkbuf_8
Xfanout50 fanout51/X vssd1 vssd1 vccd1 vccd1 _10677_/B sky130_fd_sc_hd__buf_6
Xfanout72 _12766_/A vssd1 vssd1 vccd1 vccd1 _10553_/B sky130_fd_sc_hd__buf_4
X_10603_ _10603_/A _10603_/B vssd1 vssd1 vccd1 vccd1 _10606_/B sky130_fd_sc_hd__xnor2_4
X_13322_ instruction[14] vssd1 vssd1 vccd1 vccd1 loadstore_dest[3] sky130_fd_sc_hd__buf_12
XANTENNA__07867__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout94 _07192_/Y vssd1 vssd1 vccd1 vccd1 fanout94/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11583_ curr_PC[19] _11671_/C vssd1 vssd1 vccd1 vccd1 _11583_/X sky130_fd_sc_hd__or2_1
XFILLER_0_52_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09558__S _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10534_ fanout27/X _07553_/A _10927_/A fanout26/X vssd1 vssd1 vccd1 vccd1 _10535_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13253_ _13318_/CLK _13253_/D vssd1 vssd1 vccd1 vccd1 hold159/A sky130_fd_sc_hd__dfxtp_1
X_10465_ _10464_/A _10464_/B _10464_/C vssd1 vssd1 vccd1 vccd1 _10466_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08222__B2 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08222__A1 _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13184_ _13305_/CLK hold35/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
X_10396_ _11381_/A _10369_/Y _10370_/X _10395_/X _10368_/X vssd1 vssd1 vccd1 vccd1
+ _10396_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12204_ _12204_/A _12204_/B vssd1 vssd1 vccd1 vccd1 _12208_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12135_ _12223_/B1 _12106_/X _12107_/Y _12111_/X _12134_/X vssd1 vssd1 vccd1 vccd1
+ _12135_/X sky130_fd_sc_hd__a311o_1
XANTENNA__11109__A1 _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12066_ _12060_/Y _12061_/X _12065_/X _12058_/X vssd1 vssd1 vccd1 vccd1 _12066_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09722__B2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09722__A1 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ _11017_/A _11017_/B vssd1 vssd1 vccd1 vccd1 _11018_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12013__A _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07107__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11852__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12968_ _08775_/A _12788_/B hold147/X vssd1 vssd1 vccd1 vccd1 hold148/A sky130_fd_sc_hd__a21boi_1
XANTENNA__06946__A _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ _12187_/A1 _11992_/B hold226/A vssd1 vssd1 vccd1 vccd1 _11919_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12899_ hold297/X _12955_/A2 _13168_/B1 hold217/X vssd1 vssd1 vccd1 vccd1 hold218/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07110_ _09764_/A _07110_/B vssd1 vssd1 vccd1 vccd1 _07110_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11596__A1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11596__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08090_ _08150_/A _08150_/B vssd1 vssd1 vccd1 vccd1 _08151_/A sky130_fd_sc_hd__or2_1
XANTENNA__07777__A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07041_ reg1_val[5] _07041_/B vssd1 vssd1 vccd1 vccd1 _07763_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11348__A1 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07972__B1 _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08992_ _08992_/A _08992_/B vssd1 vssd1 vccd1 vccd1 _08995_/B sky130_fd_sc_hd__xor2_4
X_07943_ _07770_/A _07770_/B _07766_/Y vssd1 vssd1 vccd1 vccd1 _07949_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_76_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07874_ _08443_/A _07874_/B vssd1 vssd1 vccd1 vccd1 _07874_/Y sky130_fd_sc_hd__xnor2_1
X_06825_ _06865_/A _06822_/Y _06823_/Y vssd1 vssd1 vccd1 vccd1 _06825_/Y sky130_fd_sc_hd__o21ai_1
X_09613_ _10156_/B2 fanout22/X _10677_/A _10156_/A1 vssd1 vssd1 vccd1 vccd1 _09614_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06756_ reg1_val[5] _06972_/C vssd1 vssd1 vccd1 vccd1 _06758_/A sky130_fd_sc_hd__or2_1
X_09544_ _09544_/A _09544_/B vssd1 vssd1 vccd1 vccd1 _09544_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12076__A2 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12577__B _12578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__B1 _11379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06687_ _06687_/A _12563_/B vssd1 vssd1 vccd1 vccd1 _06687_/Y sky130_fd_sc_hd__nor2_1
X_09475_ _09475_/A _09475_/B vssd1 vssd1 vccd1 vccd1 _09484_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_108_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08426_ _08419_/A _08419_/B _08425_/Y vssd1 vssd1 vccd1 vccd1 _08456_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_19_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11036__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08357_ _08443_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _08358_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08288_ _08342_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08343_/A sky130_fd_sc_hd__or2_1
X_07308_ _07308_/A _07308_/B vssd1 vssd1 vccd1 vccd1 _07308_/X sky130_fd_sc_hd__and2_1
XFILLER_0_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07239_ _08589_/A _07239_/B vssd1 vssd1 vccd1 vccd1 _07240_/A sky130_fd_sc_hd__xnor2_1
X_10250_ _11195_/B _10249_/X _11089_/A vssd1 vssd1 vccd1 vccd1 _10250_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07007__A2 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10181_ _10182_/A _10182_/B vssd1 vssd1 vccd1 vccd1 _10181_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08311__A _08311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09704__A1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout262 _06687_/A vssd1 vssd1 vccd1 vccd1 _06649_/A sky130_fd_sc_hd__buf_6
Xfanout273 _09197_/B vssd1 vssd1 vccd1 vccd1 _10638_/B sky130_fd_sc_hd__buf_4
Xfanout251 _06929_/X vssd1 vssd1 vccd1 vccd1 _12250_/B sky130_fd_sc_hd__clkbuf_8
Xfanout295 _13028_/A vssd1 vssd1 vccd1 vccd1 _13179_/A sky130_fd_sc_hd__buf_2
Xfanout284 _06568_/X vssd1 vssd1 vccd1 vccd1 _06898_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10314__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12768__A _12768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12822_ _12820_/X _12822_/B vssd1 vssd1 vccd1 vccd1 _13043_/A sky130_fd_sc_hd__nand2b_1
X_12753_ hold9/X _12788_/B _12752_/Y _13086_/A vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__o211a_1
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10288__A _10453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13016__A1 _07090_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11704_ _11704_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _11706_/C sky130_fd_sc_hd__nor2_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12684_ _12684_/A _12688_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[25] sky130_fd_sc_hd__xnor2_4
XFILLER_0_37_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11635_ _11635_/A _11635_/B vssd1 vssd1 vccd1 vccd1 _11814_/A sky130_fd_sc_hd__or2_1
X_11566_ _11566_/A _11566_/B vssd1 vssd1 vccd1 vccd1 _11568_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07246__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13305_ _13305_/CLK _13305_/D vssd1 vssd1 vccd1 vccd1 hold262/A sky130_fd_sc_hd__dfxtp_1
X_10517_ _10498_/A _09383_/B _10511_/X _10513_/X _10516_/X vssd1 vssd1 vccd1 vccd1
+ _10517_/X sky130_fd_sc_hd__o2111a_1
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13236_ _13305_/CLK hold170/X vssd1 vssd1 vccd1 vccd1 _13236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11497_ _11853_/A _11497_/B vssd1 vssd1 vccd1 vccd1 _11499_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_122_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10448_ _10448_/A _10592_/A _10448_/C vssd1 vssd1 vccd1 vccd1 _10464_/A sky130_fd_sc_hd__and3_1
X_10379_ hold292/A _10514_/C _09385_/C vssd1 vssd1 vccd1 vccd1 _10381_/B sky130_fd_sc_hd__o21a_1
X_13167_ _13167_/A _13167_/B _13167_/C vssd1 vssd1 vccd1 vccd1 _13167_/X sky130_fd_sc_hd__or3_1
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13098_ _13098_/A _13098_/B vssd1 vssd1 vccd1 vccd1 _13098_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08221__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12118_ _12361_/B _09972_/Y _12116_/Y _12117_/X vssd1 vssd1 vccd1 vccd1 _12118_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12049_ _11987_/A _11984_/Y _11986_/B vssd1 vssd1 vccd1 vccd1 _12053_/A sky130_fd_sc_hd__o21a_1
XANTENNA__10305__A2 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07182__A1 _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06610_ reg1_val[27] _07434_/A vssd1 vssd1 vccd1 vccd1 _06610_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07590_ _07590_/A _07590_/B vssd1 vssd1 vccd1 vccd1 _07593_/A sky130_fd_sc_hd__nor2_2
X_06541_ instruction[41] vssd1 vssd1 vccd1 vccd1 _06541_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10198__A _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09260_ _10458_/A _09260_/B vssd1 vssd1 vccd1 vccd1 _09261_/B sky130_fd_sc_hd__xnor2_2
X_08211_ _08211_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _08212_/B sky130_fd_sc_hd__or2_1
XANTENNA__08682__A1 _06989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09191_ instruction[3] _09200_/A _09200_/B instruction[4] vssd1 vssd1 vccd1 vccd1
+ _09191_/X sky130_fd_sc_hd__or4b_4
XFILLER_0_16_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08142_ _12734_/A _08348_/B _07181_/Y _08819_/B2 vssd1 vssd1 vccd1 vccd1 _08143_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08073_ _08836_/A _08073_/B vssd1 vssd1 vccd1 vccd1 _08080_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07024_ reg1_val[7] _07038_/B _07105_/A vssd1 vssd1 vccd1 vccd1 _07070_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_43_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout114_A _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08131__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__B1 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _08975_/A _08975_/B vssd1 vssd1 vccd1 vccd1 _08978_/B sky130_fd_sc_hd__xnor2_4
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _11499_/A _07926_/B vssd1 vssd1 vccd1 vccd1 _08056_/B sky130_fd_sc_hd__xnor2_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ _12730_/A _09752_/B fanout14/X _08748_/B1 vssd1 vssd1 vccd1 vccd1 _07858_/B
+ sky130_fd_sc_hd__o22a_1
X_07788_ _07778_/B _07788_/B vssd1 vssd1 vccd1 vccd1 _07789_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07712__A3 _07322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06808_ _10743_/A _06806_/Y _06807_/Y vssd1 vssd1 vccd1 vccd1 _06808_/Y sky130_fd_sc_hd__o21ai_1
X_06739_ _06739_/A _06739_/B vssd1 vssd1 vccd1 vccd1 _10373_/A sky130_fd_sc_hd__and2_1
X_09527_ _09152_/X _09156_/X _09676_/S vssd1 vssd1 vccd1 vccd1 _09527_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout27_A _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ _12762_/A fanout52/X _10677_/B _12760_/A vssd1 vssd1 vccd1 vccd1 _09459_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08409_ _08775_/A _08409_/B vssd1 vssd1 vccd1 vccd1 _08413_/A sky130_fd_sc_hd__xnor2_2
X_09389_ _12563_/A _09392_/S wire201/X _09388_/Y vssd1 vssd1 vccd1 vccd1 _09389_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11420_ _11604_/A _11420_/B vssd1 vssd1 vccd1 vccd1 _11422_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07228__A2 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11351_ _11351_/A _11351_/B vssd1 vssd1 vccd1 vccd1 _11364_/A sky130_fd_sc_hd__xor2_2
X_10302_ _10303_/A _10303_/B vssd1 vssd1 vccd1 vccd1 _10461_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11282_ _11216_/X _11316_/B _09110_/X vssd1 vssd1 vccd1 vccd1 _11282_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13021_ hold38/X hold36/X fanout1/X vssd1 vssd1 vccd1 vccd1 _13021_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__09925__A1 _09925_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09925__B2 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10233_ _09959_/Y _10487_/A _10232_/Y vssd1 vssd1 vccd1 vccd1 _10233_/Y sky130_fd_sc_hd__a21oi_1
X_10164_ _08680_/B fanout57/X _07553_/A fanout29/X vssd1 vssd1 vccd1 vccd1 _10165_/B
+ sky130_fd_sc_hd__o22ai_1
XFILLER_0_30_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10095_ _10229_/B _10229_/C vssd1 vssd1 vccd1 vccd1 _10609_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_89_628 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11496__B1 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12805_ hold289/A hold88/X vssd1 vssd1 vccd1 vccd1 _13112_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10997_ curr_PC[13] _11107_/C vssd1 vssd1 vccd1 vccd1 _10997_/X sky130_fd_sc_hd__or2_1
X_12736_ _12736_/A _12788_/B vssd1 vssd1 vccd1 vccd1 _12736_/Y sky130_fd_sc_hd__nand2_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12667_ reg1_val[22] _12714_/A vssd1 vssd1 vccd1 vccd1 _12667_/X sky130_fd_sc_hd__and2_1
XANTENNA__09600__A _09600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11618_ _11618_/A _11618_/B _11618_/C _11618_/D vssd1 vssd1 vccd1 vccd1 _11619_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__09613__B1 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08216__A _08853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12598_ reg1_val[8] _12598_/B vssd1 vssd1 vccd1 vccd1 _12599_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11549_ _11368_/Y _11456_/Y _11458_/B vssd1 vssd1 vccd1 vccd1 _11549_/X sky130_fd_sc_hd__o21a_1
X_13219_ _13248_/CLK _13219_/D vssd1 vssd1 vccd1 vccd1 hold297/A sky130_fd_sc_hd__dfxtp_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_10_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13277_/CLK sky130_fd_sc_hd__clkbuf_8
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _08761_/A _08761_/B vssd1 vssd1 vccd1 vccd1 _08834_/A sky130_fd_sc_hd__nor2_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08691_ _07988_/Y _07995_/B _07993_/Y vssd1 vssd1 vccd1 vccd1 _08700_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11487__B1 _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07711_ _07710_/B _07710_/C _09580_/A vssd1 vssd1 vccd1 vccd1 _07716_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08352__B1 _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07642_ _10452_/B2 _07034_/Y _08854_/B2 _09925_/A1 vssd1 vssd1 vccd1 vccd1 _07643_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11239__B1 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07573_ _07573_/A _07573_/B vssd1 vssd1 vccd1 vccd1 _07585_/B sky130_fd_sc_hd__xnor2_4
X_09312_ _09312_/A _09312_/B vssd1 vssd1 vccd1 vccd1 _09313_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09243_ _09243_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _09249_/A sky130_fd_sc_hd__and2_1
XFILLER_0_90_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09174_ _09172_/X _09173_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09174_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08125_ _08775_/A _08125_/B vssd1 vssd1 vccd1 vccd1 _08129_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07030__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09080__A1 _09077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08056_ _08056_/A _08056_/B vssd1 vssd1 vccd1 vccd1 _08058_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_114_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09907__B2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09907__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07007_ _09888_/B2 _08680_/B _12736_/A fanout30/X vssd1 vssd1 vccd1 vccd1 _07008_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10517__A2 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07394__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07394__B2 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ _08959_/A _08959_/B vssd1 vssd1 vccd1 vccd1 _08958_/X sky130_fd_sc_hd__and2_1
X_07909_ _07935_/B _07908_/B _07908_/C _07905_/Y vssd1 vssd1 vccd1 vccd1 _07928_/B
+ sky130_fd_sc_hd__a31o_1
X_08889_ _08889_/A _08889_/B vssd1 vssd1 vccd1 vccd1 _08891_/C sky130_fd_sc_hd__and2_1
X_10920_ _10920_/A _10920_/B vssd1 vssd1 vccd1 vccd1 _10921_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_79_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10851_ _10850_/Y _10851_/B vssd1 vssd1 vccd1 vccd1 _10851_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_94_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10782_ _10783_/A _10783_/B vssd1 vssd1 vccd1 vccd1 _10934_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07449__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12521_ _12557_/A _12521_/B vssd1 vssd1 vccd1 vccd1 _12529_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_109_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12452_ reg1_val[11] curr_PC[11] _12524_/S vssd1 vssd1 vccd1 vccd1 _12454_/B sky130_fd_sc_hd__mux2_1
XANTENNA__06763__B _07001_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11403_ _12290_/C1 _11402_/Y _11400_/X vssd1 vssd1 vccd1 vccd1 _11404_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12383_ _12563_/B _12384_/B vssd1 vssd1 vccd1 vccd1 _12394_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07082__B1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11334_ _11853_/A _11334_/B vssd1 vssd1 vccd1 vccd1 _11336_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11265_ _11266_/B _11266_/A vssd1 vssd1 vccd1 vccd1 _11365_/A sky130_fd_sc_hd__nand2b_1
X_13004_ _10015_/A _13020_/B2 hold101/X vssd1 vssd1 vccd1 vccd1 hold102/A sky130_fd_sc_hd__o21a_1
X_10216_ _10216_/A _10216_/B vssd1 vssd1 vccd1 vccd1 _10218_/A sky130_fd_sc_hd__xnor2_2
X_11196_ _10752_/S _11194_/X _11195_/X vssd1 vssd1 vccd1 vccd1 _11196_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_118_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10147_ _10147_/A _10147_/B _10147_/C vssd1 vssd1 vccd1 vccd1 _10148_/B sky130_fd_sc_hd__or3_1
X_10078_ _09940_/A _09940_/B _09939_/A vssd1 vssd1 vccd1 vccd1 _10088_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12130__A1 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07115__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11860__A _11861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12719_ hold31/X _12719_/B vssd1 vssd1 vccd1 vccd1 hold177/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11944__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11944__B2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09930_ fanout69/X _10557_/B fanout13/X _12762_/A vssd1 vssd1 vccd1 vccd1 _09931_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_68_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09861_ _09806_/A _09806_/B _09807_/Y vssd1 vssd1 vccd1 vccd1 _09955_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_0_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08812_ _08812_/A _08812_/B vssd1 vssd1 vccd1 vccd1 _08813_/B sky130_fd_sc_hd__and2_1
X_09792_ _09792_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09793_/B sky130_fd_sc_hd__xor2_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _06989_/A _11782_/A _08681_/B vssd1 vssd1 vccd1 vccd1 _08744_/C sky130_fd_sc_hd__a21o_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout181_A _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08325__B1 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout279_A _12658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08674_ _08857_/A _08674_/B _08674_/C vssd1 vssd1 vccd1 vccd1 _08677_/B sky130_fd_sc_hd__or3_1
XANTENNA__07679__A2 _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07533__D1 _12713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ _07625_/A _07625_/B vssd1 vssd1 vccd1 vccd1 _07628_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06864__A _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11770__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07556_ _07555_/B _07555_/C _10559_/A vssd1 vssd1 vccd1 vccd1 _07562_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09226_ _09226_/A _09226_/B vssd1 vssd1 vccd1 vccd1 _09328_/A sky130_fd_sc_hd__nand2_2
X_07487_ _10927_/A _10557_/B fanout83/X fanout13/X vssd1 vssd1 vccd1 vccd1 _07488_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_63_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09157_ reg1_val[30] _12563_/A _09158_/S vssd1 vssd1 vccd1 vccd1 _09157_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08108_ _08108_/A _08108_/B vssd1 vssd1 vccd1 vccd1 _08165_/A sky130_fd_sc_hd__xnor2_1
X_09088_ _09088_/A _09088_/B vssd1 vssd1 vccd1 vccd1 _12174_/A sky130_fd_sc_hd__and2_2
XFILLER_0_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08039_ _08857_/A _08039_/B vssd1 vssd1 vccd1 vccd1 _08043_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_101_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11050_ _10921_/A _10921_/B _10909_/Y vssd1 vssd1 vccd1 vccd1 _11052_/A sky130_fd_sc_hd__a21o_1
X_10001_ _10002_/B _10002_/C vssd1 vssd1 vccd1 vccd1 _10523_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11945__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09415__A _10301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11952_ _11952_/A _11952_/B _11952_/C vssd1 vssd1 vccd1 vccd1 _11953_/B sky130_fd_sc_hd__or3_1
XANTENNA__12776__A _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11883_ _11883_/A _11883_/B vssd1 vssd1 vccd1 vccd1 _11884_/B sky130_fd_sc_hd__or2_1
X_10903_ _10904_/A _10904_/B vssd1 vssd1 vccd1 vccd1 _11003_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_79_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10834_ _10834_/A _10834_/B vssd1 vssd1 vccd1 vccd1 _10837_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10426__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10426__A1 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08095__A2 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12504_ _12509_/B _12504_/B vssd1 vssd1 vccd1 vccd1 new_PC[18] sky130_fd_sc_hd__and2_4
XFILLER_0_82_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10765_ _10251_/S _09834_/X _09214_/A vssd1 vssd1 vccd1 vccd1 _10765_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_67_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10696_ _10696_/A _10696_/B vssd1 vssd1 vccd1 vccd1 _10698_/B sky130_fd_sc_hd__xor2_1
X_12435_ _12436_/A _12436_/B _12436_/C vssd1 vssd1 vccd1 vccd1 _12443_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12366_ hold149/A _12364_/X _12365_/Y vssd1 vssd1 vccd1 vccd1 _12366_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11317_ _12230_/A _11730_/A vssd1 vssd1 vccd1 vccd1 _11317_/X sky130_fd_sc_hd__and2_1
XFILLER_0_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12297_ _12272_/Y _12273_/X _12276_/Y _12277_/X _12296_/X vssd1 vssd1 vccd1 vccd1
+ _12297_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09309__B _09309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11248_ _07261_/Y _12349_/A _11247_/X vssd1 vssd1 vccd1 vccd1 _11250_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_38_56 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11179_ _11462_/B _11179_/B vssd1 vssd1 vccd1 vccd1 _11215_/D sky130_fd_sc_hd__xnor2_1
XANTENNA__06949__A _11194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10901__A2 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08307__B1 _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07530__A1 _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10665__A1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10665__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08390_ _08390_/A _08390_/B _08390_/C vssd1 vssd1 vccd1 vccd1 _08390_/X sky130_fd_sc_hd__and3_1
XFILLER_0_58_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07410_ _08897_/A _07412_/B vssd1 vssd1 vccd1 vccd1 _07410_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07341_ _10180_/A _07341_/B vssd1 vssd1 vccd1 vccd1 _07344_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07272_ _07272_/A _07272_/B vssd1 vssd1 vccd1 vccd1 _07274_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09011_ _09011_/A _09011_/B vssd1 vssd1 vccd1 vccd1 _09049_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold101 hold101/A vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 hold134/A vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 hold112/A vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold156 hold156/A vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 hold145/A vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 hold167/A vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold178 hold178/A vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 hold189/A vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09338__A2 _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09913_ _09913_/A _10037_/B _09913_/C vssd1 vssd1 vccd1 vccd1 _10006_/A sky130_fd_sc_hd__and3_1
X_09844_ _11400_/A _09842_/X _09843_/Y _11099_/B reg1_val[4] vssd1 vssd1 vccd1 vccd1
+ _09844_/X sky130_fd_sc_hd__o32a_1
XANTENNA__11765__A _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12342__A1 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12893__A2 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _09775_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _09777_/B sky130_fd_sc_hd__xnor2_2
X_06987_ _10565_/A _06987_/B _10555_/A vssd1 vssd1 vccd1 vccd1 _06989_/A sky130_fd_sc_hd__or3b_4
X_08726_ _10565_/A _08726_/B vssd1 vssd1 vccd1 vccd1 _08728_/B sky130_fd_sc_hd__xnor2_1
X_08657_ _08657_/A _08657_/B vssd1 vssd1 vccd1 vccd1 _08658_/B sky130_fd_sc_hd__xnor2_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10656__B2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10656__A1 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07608_ _07588_/A _07588_/B _07586_/Y vssd1 vssd1 vccd1 vccd1 _07611_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__06594__A _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08588_ _08588_/A _08588_/B vssd1 vssd1 vccd1 vccd1 _08598_/S sky130_fd_sc_hd__nor2_1
XFILLER_0_49_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13070__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08077__A2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07539_ _07539_/A _07539_/B vssd1 vssd1 vccd1 vccd1 _07541_/B sky130_fd_sc_hd__xnor2_2
X_10550_ _10550_/A _10550_/B vssd1 vssd1 vccd1 vccd1 _10552_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09209_ _09209_/A vssd1 vssd1 vccd1 vccd1 _09211_/A sky130_fd_sc_hd__inv_2
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10481_ _10481_/A _10481_/B vssd1 vssd1 vccd1 vccd1 _10482_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_106_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12220_ _12312_/A _12220_/B vssd1 vssd1 vccd1 vccd1 _12317_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12151_ _12200_/A _12151_/B _12151_/C vssd1 vssd1 vccd1 vccd1 _12152_/B sky130_fd_sc_hd__and3_1
XFILLER_0_102_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11102_ _09198_/X _11095_/Y _11098_/Y _11101_/X vssd1 vssd1 vccd1 vccd1 _11102_/X
+ sky130_fd_sc_hd__a211o_1
X_12082_ _12152_/A _12082_/B vssd1 vssd1 vccd1 vccd1 _12083_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11136__A2 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11033_ _11034_/A _11034_/B vssd1 vssd1 vccd1 vccd1 _11121_/A sky130_fd_sc_hd__and2_1
XANTENNA__10895__B2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10895__A1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12984_ _08733_/A _12744_/B hold133/X vssd1 vssd1 vccd1 vccd1 _13262_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_87_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11935_ _11935_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _11936_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_39_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11866_ _12776_/A fanout15/X fanout6/X _11935_/A vssd1 vssd1 vccd1 vccd1 _11867_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10817_ _10696_/A _10696_/B _10694_/X vssd1 vssd1 vccd1 vccd1 _10826_/A sky130_fd_sc_hd__a21o_1
X_11797_ _11797_/A _11797_/B _11797_/C vssd1 vssd1 vccd1 vccd1 _11798_/B sky130_fd_sc_hd__or3_1
X_10748_ _10625_/B _10630_/B _10625_/A vssd1 vssd1 vccd1 vccd1 _10753_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_113_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12418_ _12588_/B _12419_/B vssd1 vssd1 vccd1 vccd1 _12429_/A sky130_fd_sc_hd__nand2_1
X_10679_ _10678_/B _10678_/C _11429_/A vssd1 vssd1 vccd1 vccd1 _10683_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12021__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__B1 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12349_ _12349_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _12350_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_10_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06910_ instruction[20] _06552_/X _06909_/X _06678_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[2]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__11127__A2 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07890_ _08855_/A _07891_/B vssd1 vssd1 vccd1 vccd1 _07892_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06679__A _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07306__C_N _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10335__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06841_ _12045_/A _06840_/X _06839_/X vssd1 vssd1 vccd1 vccd1 _06841_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_4_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06772_ reg2_val[2] _06778_/B vssd1 vssd1 vccd1 vccd1 _06772_/X sky130_fd_sc_hd__and2_1
X_09560_ _10617_/A _10273_/D vssd1 vssd1 vccd1 vccd1 _09666_/A sky130_fd_sc_hd__or2_1
XFILLER_0_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08511_ _09622_/A _08511_/B vssd1 vssd1 vccd1 vccd1 _08540_/A sky130_fd_sc_hd__xor2_2
X_09491_ _09237_/A _09237_/B _09239_/B _09242_/A vssd1 vssd1 vccd1 vccd1 _09496_/A
+ sky130_fd_sc_hd__a31o_2
X_08442_ _10149_/A _07149_/Y _07155_/X _10035_/A vssd1 vssd1 vccd1 vccd1 _08443_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07503__B2 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07503__A1 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08373_ _08373_/A _08373_/B vssd1 vssd1 vccd1 vccd1 _08375_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__06657__A2_N _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07303__A _07303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout144_A _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07324_ _07324_/A _07325_/B vssd1 vssd1 vccd1 vccd1 _07324_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_116_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07255_ reg1_val[17] _07255_/B vssd1 vssd1 vccd1 vccd1 _07255_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08134__A _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07186_ reg1_val[13] reg1_val[14] _07165_/B _07105_/A vssd1 vssd1 vccd1 vccd1 _07188_/B
+ sky130_fd_sc_hd__o31a_4
XFILLER_0_14_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08231__A2 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09827_ _06868_/C _09825_/X _09826_/Y vssd1 vssd1 vccd1 vccd1 _09827_/X sky130_fd_sc_hd__o21a_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09758_ _09758_/A _09758_/B vssd1 vssd1 vccd1 vccd1 _09761_/A sky130_fd_sc_hd__or2_1
XFILLER_0_96_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08709_ _07949_/A _07949_/B _07947_/X vssd1 vssd1 vccd1 vccd1 _08712_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_69_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout57_A _07179_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09689_ _12361_/B _09682_/X _09688_/X _09851_/B vssd1 vssd1 vccd1 vccd1 _09707_/A
+ sky130_fd_sc_hd__o211a_1
X_11720_ _11722_/A _11722_/B _11722_/C vssd1 vssd1 vccd1 vccd1 _11721_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11651_ reg1_val[20] curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11652_/B sky130_fd_sc_hd__or2_1
Xfanout40 _07530_/X vssd1 vssd1 vccd1 vccd1 _12349_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout73 _07069_/Y vssd1 vssd1 vccd1 vccd1 _12766_/A sky130_fd_sc_hd__buf_6
X_11582_ _11381_/A _11558_/X _11559_/Y _11581_/Y _11557_/X vssd1 vssd1 vccd1 vccd1
+ _11582_/X sky130_fd_sc_hd__a311o_2
XANTENNA__12251__B1 _12345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout51 _07262_/X vssd1 vssd1 vccd1 vccd1 fanout51/X sky130_fd_sc_hd__buf_8
Xfanout62 _12772_/A vssd1 vssd1 vccd1 vccd1 fanout62/X sky130_fd_sc_hd__buf_6
X_10602_ _10602_/A _10602_/B vssd1 vssd1 vccd1 vccd1 _10603_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout84 _07305_/Y vssd1 vssd1 vccd1 vccd1 fanout84/X sky130_fd_sc_hd__clkbuf_8
Xfanout95 _08217_/B vssd1 vssd1 vccd1 vccd1 fanout95/X sky130_fd_sc_hd__buf_6
X_13321_ instruction[13] vssd1 vssd1 vccd1 vccd1 loadstore_dest[2] sky130_fd_sc_hd__buf_12
X_10533_ _10533_/A _10533_/B vssd1 vssd1 vccd1 vccd1 _10573_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09094__A1_N _08932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13252_ _13318_/CLK _13252_/D vssd1 vssd1 vccd1 vccd1 hold157/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10464_ _10464_/A _10464_/B _10464_/C vssd1 vssd1 vccd1 vccd1 _10466_/B sky130_fd_sc_hd__or3_1
X_13183_ _13318_/CLK _13183_/D vssd1 vssd1 vccd1 vccd1 hold152/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08222__A2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08758__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10395_ _10395_/A _10395_/B _10395_/C vssd1 vssd1 vccd1 vccd1 _10395_/X sky130_fd_sc_hd__or3_1
XFILLER_0_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12203_ _12203_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _12204_/B sky130_fd_sc_hd__or2_1
XFILLER_0_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ _11381_/A _12132_/Y _12133_/X _12130_/X vssd1 vssd1 vccd1 vccd1 _12134_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__06784__A2 _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12065_ _09184_/X _10111_/Y _10118_/Y _09115_/X _12064_/X vssd1 vssd1 vccd1 vccd1
+ _12065_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09722__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ _11017_/A _11017_/B vssd1 vssd1 vccd1 vccd1 _11158_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12013__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07107__B _07115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11817__B1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09603__A _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12967_ hold159/A _12723_/A _13170_/B hold146/X _13066_/A vssd1 vssd1 vccd1 vccd1
+ hold147/A sky130_fd_sc_hd__o221a_1
XFILLER_0_87_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06946__B _12370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11918_ hold200/A _11918_/B vssd1 vssd1 vccd1 vccd1 _11992_/B sky130_fd_sc_hd__or2_1
X_12898_ _13169_/A hold249/X vssd1 vssd1 vccd1 vccd1 _13219_/D sky130_fd_sc_hd__and2_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07497__B1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07123__A _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11849_ _11849_/A _11849_/B vssd1 vssd1 vccd1 vccd1 _11886_/A sky130_fd_sc_hd__nand2_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12242__B1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11596__A2 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07040_ reg1_val[4] _07105_/B _07105_/A vssd1 vssd1 vccd1 vccd1 _07041_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_42_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11348__A2 _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07793__A _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10556__B1 _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08991_ _08984_/A _08984_/B _08985_/Y vssd1 vssd1 vccd1 vccd1 _08995_/A sky130_fd_sc_hd__a21bo_2
X_07942_ _08019_/A _08019_/B _07886_/X vssd1 vssd1 vccd1 vccd1 _08638_/A sky130_fd_sc_hd__a21oi_4
X_07873_ _12760_/A _08692_/A2 _08692_/B1 _09925_/A1 vssd1 vssd1 vccd1 vccd1 _07874_/B
+ sky130_fd_sc_hd__o22a_1
X_06824_ _06865_/A _06822_/Y _06823_/Y vssd1 vssd1 vccd1 vccd1 _06824_/X sky130_fd_sc_hd__o21a_1
X_09612_ _09612_/A _09612_/B vssd1 vssd1 vccd1 vccd1 _09615_/B sky130_fd_sc_hd__xor2_1
X_09543_ _12563_/A _09392_/S _09362_/S _09180_/A vssd1 vssd1 vccd1 vccd1 _09544_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout261_A _12284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06755_ reg1_val[5] _06972_/C vssd1 vssd1 vccd1 vccd1 _06755_/Y sky130_fd_sc_hd__nor2_1
X_06686_ instruction[0] instruction[1] instruction[2] instruction[26] pred_val vssd1
+ vssd1 vccd1 vccd1 _12563_/B sky130_fd_sc_hd__o311a_4
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09474_ _09474_/A _09474_/B vssd1 vssd1 vccd1 vccd1 _09475_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08425_ _08433_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08425_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_65_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08356_ _10144_/B2 _08692_/B1 _08835_/B1 _08692_/A2 vssd1 vssd1 vccd1 vccd1 _08357_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11036__B2 _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11036__A1 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07307_ _10559_/A _11429_/B _10180_/A vssd1 vssd1 vccd1 vccd1 _07308_/B sky130_fd_sc_hd__nand3b_4
XANTENNA__12593__B _12593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08287_ _08287_/A _08287_/B vssd1 vssd1 vccd1 vccd1 _08342_/B sky130_fd_sc_hd__xnor2_1
X_07238_ _12782_/A _08588_/B _09273_/A1 fanout22/X vssd1 vssd1 vccd1 vccd1 _07239_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07169_ reg1_val[10] reg1_val[11] _07027_/B _07105_/A vssd1 vssd1 vccd1 vccd1 _07170_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_42_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10547__B1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06766__A2 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10180_ _10180_/A _10180_/B vssd1 vssd1 vccd1 vccd1 _10182_/B sky130_fd_sc_hd__xnor2_1
Xfanout230 _06579_/Y vssd1 vssd1 vccd1 vccd1 _06680_/B1 sky130_fd_sc_hd__buf_4
Xfanout241 _09193_/X vssd1 vssd1 vccd1 vccd1 _12277_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout263 _06687_/A vssd1 vssd1 vccd1 vccd1 _06641_/A sky130_fd_sc_hd__clkbuf_4
Xfanout252 _06929_/X vssd1 vssd1 vccd1 vccd1 _11923_/A2 sky130_fd_sc_hd__buf_2
Xfanout274 _07105_/A vssd1 vssd1 vccd1 vccd1 _07165_/A sky130_fd_sc_hd__buf_4
Xfanout285 _06633_/B vssd1 vssd1 vccd1 vccd1 _06678_/B sky130_fd_sc_hd__clkbuf_8
Xfanout296 _06547_/Y vssd1 vssd1 vccd1 vccd1 _13028_/A sky130_fd_sc_hd__clkbuf_4
X_12821_ hold288/A hold13/X vssd1 vssd1 vccd1 vccd1 _12822_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_88_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08039__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12752_ _12752_/A _12788_/B vssd1 vssd1 vccd1 vccd1 _12752_/Y sky130_fd_sc_hd__nand2_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ reg1_val[25] _12708_/B vssd1 vssd1 vccd1 vccd1 _12688_/B sky130_fd_sc_hd__xnor2_4
X_11703_ _11620_/A _11619_/B _11619_/A vssd1 vssd1 vccd1 vccd1 _11712_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12784__A _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11456_/Y _11548_/A _11548_/B vssd1 vssd1 vccd1 vccd1 _11634_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__11578__A2 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06782__A _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11565_ reg1_val[19] curr_PC[19] vssd1 vssd1 vccd1 vccd1 _11566_/B sky130_fd_sc_hd__or2_1
XFILLER_0_80_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10508__S _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10786__B1 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10516_ hold272/A _09385_/C _10635_/B _10515_/Y _12339_/B1 vssd1 vssd1 vccd1 vccd1
+ _10516_/X sky130_fd_sc_hd__a311o_1
X_13304_ _13305_/CLK _13304_/D vssd1 vssd1 vccd1 vccd1 hold256/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11496_ fanout33/X _12203_/A fanout19/X _10553_/A vssd1 vssd1 vccd1 vccd1 _11497_/B
+ sky130_fd_sc_hd__o22a_1
X_13235_ _13312_/CLK _13235_/D vssd1 vssd1 vccd1 vccd1 hold168/A sky130_fd_sc_hd__dfxtp_1
X_10447_ _10446_/A _10446_/B _10446_/C vssd1 vssd1 vccd1 vccd1 _10448_/C sky130_fd_sc_hd__o21ai_1
X_13166_ _13166_/A _13166_/B vssd1 vssd1 vccd1 vccd1 _13311_/D sky130_fd_sc_hd__and2_1
XFILLER_0_103_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10378_ _07015_/B _06928_/X _10638_/B _06739_/A _10377_/Y vssd1 vssd1 vccd1 vccd1
+ _10378_/X sky130_fd_sc_hd__a221o_1
X_13097_ _13097_/A _13097_/B vssd1 vssd1 vccd1 vccd1 _13098_/B sky130_fd_sc_hd__nand2_1
X_12117_ _12112_/X _12114_/X _12115_/Y _11197_/S vssd1 vssd1 vccd1 vccd1 _12117_/X
+ sky130_fd_sc_hd__a31o_1
X_12048_ _11820_/A _09079_/A _09079_/B _11184_/A _12047_/Y vssd1 vssd1 vccd1 vccd1
+ _12048_/X sky130_fd_sc_hd__a311o_1
XANTENNA__06957__A _11780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06540_ _09180_/A vssd1 vssd1 vccd1 vccd1 _06540_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08210_ _08630_/A _08630_/B vssd1 vssd1 vccd1 vccd1 _08210_/X sky130_fd_sc_hd__and2_1
XANTENNA__08682__A2 _11782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06692__A _12641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09190_ instruction[3] _09200_/A instruction[5] instruction[4] vssd1 vssd1 vccd1
+ vccd1 _09197_/B sky130_fd_sc_hd__and4bb_2
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08141_ _08144_/A _08144_/B vssd1 vssd1 vccd1 vccd1 _08141_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08072_ _08748_/B1 _08134_/B fanout51/X _08821_/A vssd1 vssd1 vccd1 vccd1 _08073_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13021__C fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07642__B1 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07023_ _07023_/A _07077_/B vssd1 vssd1 vccd1 vccd1 _07023_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout107_A _07031_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07945__A1 _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07945__B2 _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ _08974_/A _08974_/B vssd1 vssd1 vccd1 vccd1 _08975_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07925_ _08748_/B1 _09752_/B fanout14/X _08821_/A vssd1 vssd1 vccd1 vccd1 _07926_/B
+ sky130_fd_sc_hd__o22a_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__buf_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_07856_ _07932_/A vssd1 vssd1 vccd1 vccd1 _07856_/Y sky130_fd_sc_hd__inv_2
XANTENNA__12588__B _12588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06586__B _06633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07787_ _07785_/A _07785_/C _07785_/B vssd1 vssd1 vccd1 vccd1 _07790_/B sky130_fd_sc_hd__a21oi_1
X_06807_ reg1_val[11] _06807_/B vssd1 vssd1 vccd1 vccd1 _06807_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_78_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06738_ reg1_val[8] _07015_/B vssd1 vssd1 vccd1 vccd1 _06739_/B sky130_fd_sc_hd__nand2_1
X_09526_ _09522_/X _09525_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _09526_/X sky130_fd_sc_hd__mux2_1
X_09457_ _10894_/A _09457_/B vssd1 vssd1 vccd1 vccd1 _09461_/A sky130_fd_sc_hd__xnor2_1
X_06669_ instruction[28] _06678_/B vssd1 vssd1 vccd1 vccd1 _12573_/B sky130_fd_sc_hd__and2_4
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08408_ _08837_/B2 _09618_/B2 _09618_/A1 _07969_/A vssd1 vssd1 vccd1 vccd1 _08409_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09388_ _09679_/S _12250_/B _09387_/X vssd1 vssd1 vccd1 vccd1 _09388_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12757__A1 _11147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08339_ _08339_/A _08339_/B vssd1 vssd1 vccd1 vccd1 _08340_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07633__B1 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11350_ _11350_/A _11350_/B vssd1 vssd1 vccd1 vccd1 _11351_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10301_ _10301_/A _10301_/B vssd1 vssd1 vccd1 vccd1 _10303_/B sky130_fd_sc_hd__xnor2_1
X_13020_ hold38/X _13020_/A2 _11147_/B _13020_/B2 _13019_/Y vssd1 vssd1 vccd1 vccd1
+ hold39/A sky130_fd_sc_hd__o221a_1
XANTENNA__12543__S _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11281_ _11460_/A _11281_/B vssd1 vssd1 vccd1 vccd1 _11316_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09925__A2 _07322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10232_ _09956_/X _10092_/X _10093_/X vssd1 vssd1 vccd1 vccd1 _10232_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10163_ _10280_/A _10163_/B vssd1 vssd1 vccd1 vccd1 _10167_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09689__A1 _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11683__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ _10094_/A _10094_/B vssd1 vssd1 vccd1 vccd1 _10361_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_88_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11496__B2 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11496__A1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10299__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12804_ hold23/X hold280/A vssd1 vssd1 vccd1 vccd1 _12804_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_97_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12996__A1 _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10996_ _10967_/X _10995_/X _12345_/A vssd1 vssd1 vccd1 vccd1 _10996_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12735_ hold27/X _12788_/B _12734_/Y _13086_/A vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__o211a_1
XFILLER_0_96_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12678_/B _12666_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[21] sky130_fd_sc_hd__xor2_4
XANTENNA__09600__B _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12597_ reg1_val[8] _12598_/B vssd1 vssd1 vccd1 vccd1 _12597_/Y sky130_fd_sc_hd__nor2_1
X_11617_ _11618_/A _11618_/B _11618_/C _11618_/D vssd1 vssd1 vccd1 vccd1 _11619_/A
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__09613__A1 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09613__B2 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12019__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11548_ _11548_/A _11548_/B vssd1 vssd1 vccd1 vccd1 _11635_/B sky130_fd_sc_hd__or2_1
XFILLER_0_13_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11479_ _10992_/Y _11478_/X _11831_/S vssd1 vssd1 vccd1 vccd1 _11479_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_110_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08232__A _08232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13218_ _13248_/CLK _13218_/D vssd1 vssd1 vccd1 vccd1 _13218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13149_ _13149_/A _13149_/B vssd1 vssd1 vccd1 vccd1 _13149_/Y sky130_fd_sc_hd__xnor2_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ _09580_/A _07710_/B _07710_/C vssd1 vssd1 vccd1 vccd1 _07716_/A sky130_fd_sc_hd__nand3_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11593__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06687__A _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08690_ _08689_/B _08689_/C _08689_/A vssd1 vssd1 vccd1 vccd1 _08701_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07641_ _07637_/A _07637_/B _08907_/A vssd1 vssd1 vccd1 vccd1 _07651_/B sky130_fd_sc_hd__a21bo_1
X_07572_ _09775_/A _07572_/B vssd1 vssd1 vccd1 vccd1 _07585_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11239__A1 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11239__B2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09311_ _09312_/A _09312_/B vssd1 vssd1 vccd1 vccd1 _09311_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_118_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07863__B1 _08672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09242_ _09242_/A _09242_/B vssd1 vssd1 vccd1 vccd1 _09314_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12739__A1 _10035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09173_ reg1_val[23] reg1_val[8] _09173_/S vssd1 vssd1 vccd1 vccd1 _09173_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_113_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08124_ _08774_/A2 fanout84/X fanout82/X _08774_/B1 vssd1 vssd1 vccd1 vccd1 _08125_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout224_A _06964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08055_ _08055_/A _08055_/B _08055_/C vssd1 vssd1 vccd1 vccd1 _08059_/A sky130_fd_sc_hd__or3_1
XFILLER_0_114_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10672__A _11780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07006_ _12019_/A _11933_/A _07005_/Y vssd1 vssd1 vccd1 vccd1 _07006_/Y sky130_fd_sc_hd__a21boi_4
XANTENNA__09907__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07394__A2 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ _08957_/A _08957_/B vssd1 vssd1 vccd1 vccd1 _08959_/B sky130_fd_sc_hd__xnor2_2
X_07908_ _07935_/B _07908_/B _07908_/C vssd1 vssd1 vccd1 vccd1 _08055_/A sky130_fd_sc_hd__and3_1
X_08888_ _08888_/A _08888_/B vssd1 vssd1 vccd1 vccd1 _08889_/B sky130_fd_sc_hd__nand2_1
X_07839_ _07840_/A _07840_/B vssd1 vssd1 vccd1 vccd1 _07839_/Y sky130_fd_sc_hd__nand2b_1
X_10850_ _10850_/A _10850_/B vssd1 vssd1 vccd1 vccd1 _10850_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_94_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _09660_/A _09509_/B _09509_/C _09660_/C vssd1 vssd1 vccd1 vccd1 wire4/A sky130_fd_sc_hd__nor4_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10269__D _10269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10781_ _12255_/B _10781_/B vssd1 vssd1 vccd1 vccd1 _10783_/B sky130_fd_sc_hd__xnor2_1
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ reg1_val[21] curr_PC[21] _12524_/S vssd1 vssd1 vccd1 vccd1 _12521_/B sky130_fd_sc_hd__mux2_4
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12451_ _12457_/B _12451_/B vssd1 vssd1 vccd1 vccd1 new_PC[10] sky130_fd_sc_hd__and2_4
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11402_ hold178/A _11402_/B vssd1 vssd1 vccd1 vccd1 _11402_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12382_ _12563_/A curr_PC[1] _12382_/S vssd1 vssd1 vccd1 vccd1 _12384_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07082__A1 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07082__B2 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11678__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11333_ _10553_/A _12150_/A _12150_/B fanout33/X vssd1 vssd1 vccd1 vccd1 _11334_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11264_ _11264_/A _11264_/B vssd1 vssd1 vccd1 vccd1 _11266_/B sky130_fd_sc_hd__xnor2_1
X_13003_ hold126/A _13013_/A2 _13020_/A2 hold100/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold101/A sky130_fd_sc_hd__o221a_1
XANTENNA__12363__C1 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ _10215_/A _10215_/B vssd1 vssd1 vccd1 vccd1 _10216_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07891__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11195_ _11195_/A _11195_/B _11195_/C vssd1 vssd1 vccd1 vccd1 _11195_/X sky130_fd_sc_hd__and3_1
XANTENNA__10913__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ _10147_/A _10147_/B _10147_/C vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__o21ai_1
X_10077_ _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10090_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_97_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07115__B _07115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10979_ _11089_/A _10979_/B vssd1 vssd1 vccd1 vccd1 _10979_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12718_ _12719_/B vssd1 vssd1 vccd1 vccd1 _12718_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09330__B _09331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12649_ reg1_val[18] _12714_/A vssd1 vssd1 vccd1 vccd1 _12650_/B sky130_fd_sc_hd__or2_1
XFILLER_0_5_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11944__A2 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13146__B2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09860_ _09811_/A _09811_/B _09809_/X vssd1 vssd1 vccd1 vccd1 _09958_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08573__A1 _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _08780_/A _08780_/B _08778_/X vssd1 vssd1 vccd1 vccd1 _08818_/A sky130_fd_sc_hd__o21a_1
X_09791_ _09792_/A _09792_/B vssd1 vssd1 vccd1 vccd1 _09791_/Y sky130_fd_sc_hd__nand2_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _09600_/A _09294_/A vssd1 vssd1 vccd1 vccd1 _08744_/B sky130_fd_sc_hd__nand2_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08325__A1 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08325__B2 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08673_ _07195_/A _07195_/B _08835_/B1 vssd1 vssd1 vccd1 vccd1 _08674_/C sky130_fd_sc_hd__a21oi_2
XANTENNA__07306__A _10180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07624_ _07624_/A _07624_/B vssd1 vssd1 vccd1 vccd1 _07700_/A sky130_fd_sc_hd__xor2_2
XANTENNA_fanout174_A _06963_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07555_ _10559_/A _07555_/B _07555_/C vssd1 vssd1 vccd1 vccd1 _07562_/A sky130_fd_sc_hd__and3_1
XANTENNA__06864__B _12726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07486_ _07451_/A _07451_/B _07448_/A vssd1 vssd1 vccd1 vccd1 _07496_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09225_ _07620_/A _07620_/B _07618_/X vssd1 vssd1 vccd1 vccd1 _09331_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_91_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09156_ _09154_/X _09155_/X _09359_/S vssd1 vssd1 vccd1 vccd1 _09156_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08107_ _08107_/A _08107_/B vssd1 vssd1 vccd1 vccd1 _08108_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_114_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09087_ _09086_/B _09086_/C _09103_/A vssd1 vssd1 vccd1 vccd1 _09088_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11498__A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08038_ _12734_/A _08217_/B fanout55/X _08819_/B2 vssd1 vssd1 vccd1 vccd1 _08039_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13137__B2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10000_ _12005_/A _09996_/X _09997_/X _09999_/Y vssd1 vssd1 vccd1 vccd1 dest_val[5]
+ sky130_fd_sc_hd__a22o_4
XANTENNA_fanout87_A _08842_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ reg1_val[5] curr_PC[5] vssd1 vssd1 vccd1 vccd1 _09989_/Y sky130_fd_sc_hd__nor2_1
X_11951_ _11952_/A _11952_/B _11952_/C vssd1 vssd1 vccd1 vccd1 _12032_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11882_ _11883_/A _11883_/B vssd1 vssd1 vccd1 vccd1 _11964_/A sky130_fd_sc_hd__nand2_1
X_10902_ _11780_/A _10902_/B vssd1 vssd1 vccd1 vccd1 _10904_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10833_ _10831_/Y _10833_/B vssd1 vssd1 vccd1 vccd1 _10834_/B sky130_fd_sc_hd__and2b_1
X_10764_ _06866_/A _09383_/B _10759_/Y _10760_/X _10763_/Y vssd1 vssd1 vccd1 vccd1
+ _10764_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_13_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10426__A2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12503_ _12515_/A _12515_/B _12516_/B vssd1 vssd1 vccd1 vccd1 _12504_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_66_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10695_ _10695_/A _10695_/B vssd1 vssd1 vccd1 vccd1 _10696_/B sky130_fd_sc_hd__xnor2_1
X_12434_ _12443_/A _12434_/B vssd1 vssd1 vccd1 vccd1 _12436_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13099__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12365_ hold149/A _12364_/X _09198_/X vssd1 vssd1 vccd1 vccd1 _12365_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__13128__B2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11316_ _11316_/A _11316_/B _11316_/C _10523_/Y vssd1 vssd1 vccd1 vccd1 _11730_/A
+ sky130_fd_sc_hd__or4b_2
X_12296_ _09205_/B _12283_/X _12284_/Y _12295_/X _12280_/X vssd1 vssd1 vccd1 vccd1
+ _12296_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_50_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11247_ _07260_/B fanout8/X _11429_/A vssd1 vssd1 vccd1 vccd1 _11247_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11178_ _10734_/C _11174_/Y _11177_/X vssd1 vssd1 vccd1 vccd1 _11179_/B sky130_fd_sc_hd__o21ai_4
X_10129_ reg1_val[6] curr_PC[6] vssd1 vssd1 vccd1 vccd1 _10129_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06949__B _07279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07126__A _07157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06965__A _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10665__A2 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07340_ _10927_/A fanout52/X _10677_/B fanout83/X vssd1 vssd1 vccd1 vccd1 _07341_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09010_ _09010_/A _09010_/B vssd1 vssd1 vccd1 vccd1 _09010_/Y sky130_fd_sc_hd__nand2_1
X_07271_ _07272_/A _07272_/B vssd1 vssd1 vccd1 vccd1 _07271_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13119__B2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold113/A vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold157 hold157/A vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 hold146/A vssd1 vssd1 vccd1 vccd1 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12327__C1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold179 hold179/A vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09338__A3 _09283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09912_ _10037_/A _09911_/C _09911_/A vssd1 vssd1 vccd1 vccd1 _09913_/C sky130_fd_sc_hd__a21o_1
X_09843_ _09842_/B _10122_/C hold288/A vssd1 vssd1 vccd1 vccd1 _09843_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_95_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08420__A _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09743__B1 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ _06986_/A _06986_/B vssd1 vssd1 vccd1 vccd1 _10149_/A sky130_fd_sc_hd__xnor2_4
X_09774_ _09888_/B2 _07278_/B fanout7/X _12736_/A vssd1 vssd1 vccd1 vccd1 _09775_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ _07969_/A fanout47/X fanout12/X _12734_/A vssd1 vssd1 vccd1 vccd1 _08726_/B
+ sky130_fd_sc_hd__o22a_1
X_08656_ _08657_/B _08657_/A vssd1 vssd1 vccd1 vccd1 _08656_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_96_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10656__A2 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _08595_/A _08587_/B vssd1 vssd1 vccd1 vccd1 _08592_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09251__A _10453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07607_ _07603_/A _07602_/B _07600_/X vssd1 vssd1 vccd1 vccd1 _07612_/A sky130_fd_sc_hd__a21o_2
XANTENNA__06594__B _12607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07538_ _07538_/A _07538_/B vssd1 vssd1 vccd1 vccd1 _07539_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07469_ _10306_/A _07469_/B vssd1 vssd1 vccd1 vccd1 _07471_/B sky130_fd_sc_hd__xor2_1
X_09208_ _09679_/S _09213_/B _09207_/X vssd1 vssd1 vccd1 vccd1 _09209_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10480_ _10481_/A _10481_/B vssd1 vssd1 vccd1 vccd1 _10480_/X sky130_fd_sc_hd__and2_1
X_09139_ reg1_val[13] reg1_val[18] _09172_/S vssd1 vssd1 vccd1 vccd1 _09139_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10014__A1_N _09295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12150_ _12150_/A _12150_/B _12304_/B _12088_/A vssd1 vssd1 vccd1 vccd1 _12151_/C
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_20_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06752__C_N _12588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ _06704_/B wire201/X _11838_/A2 _06705_/A _11100_/X vssd1 vssd1 vccd1 vccd1
+ _11101_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_20_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10860__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _12081_/A _12081_/B vssd1 vssd1 vccd1 vccd1 _12082_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12333__A2 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09426__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11032_ _12022_/A _11032_/B vssd1 vssd1 vccd1 vccd1 _11034_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06769__B _11194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10895__A2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12983_ hold132/X _12723_/A _13020_/A2 hold98/X _13066_/A vssd1 vssd1 vccd1 vccd1
+ hold133/A sky130_fd_sc_hd__o221a_1
XFILLER_0_87_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11844__A1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11934_ _07005_/Y fanout8/X _11933_/Y _11780_/A vssd1 vssd1 vccd1 vccd1 _12011_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_95_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11865_ _11786_/A _11786_/B _11778_/A vssd1 vssd1 vccd1 vccd1 _11881_/A sky130_fd_sc_hd__o21ai_1
X_10816_ _10816_/A _10816_/B vssd1 vssd1 vccd1 vccd1 _10827_/A sky130_fd_sc_hd__nand2_1
X_11796_ _11797_/A _11797_/B _11797_/C vssd1 vssd1 vccd1 vccd1 _11849_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10747_ _10747_/A _10747_/B vssd1 vssd1 vccd1 vccd1 _10753_/A sky130_fd_sc_hd__or2_1
XFILLER_0_55_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_11_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10678_ _11429_/A _10678_/B _10678_/C vssd1 vssd1 vccd1 vccd1 _10683_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_113_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08225__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12417_ reg1_val[6] curr_PC[6] _12524_/S vssd1 vssd1 vccd1 vccd1 _12419_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12021__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08776__A1 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12021__B2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08776__B2 _09925_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12348_ _12348_/A _12348_/B vssd1 vssd1 vccd1 vccd1 _12350_/A sky130_fd_sc_hd__xnor2_1
X_12279_ _12279_/A _12279_/B vssd1 vssd1 vccd1 vccd1 _12279_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06679__B _12568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06840_ reg1_val[24] _07126_/B vssd1 vssd1 vccd1 vccd1 _06840_/X sky130_fd_sc_hd__and2_1
XANTENNA__10335__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10335__B2 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06771_ _06768_/Y _06771_/B vssd1 vssd1 vccd1 vccd1 _06868_/D sky130_fd_sc_hd__nand2b_1
XFILLER_0_65_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08510_ _09772_/A _08588_/B _09273_/A1 _09478_/B2 vssd1 vssd1 vccd1 vccd1 _08511_/B
+ sky130_fd_sc_hd__o22a_1
X_09490_ _09314_/A _09313_/B _09311_/Y vssd1 vssd1 vccd1 vccd1 _09500_/A sky130_fd_sc_hd__a21o_1
X_08441_ _08445_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08441_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07503__A2 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08372_ _08372_/A _08372_/B vssd1 vssd1 vccd1 vccd1 _08375_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10010__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07323_ _07015_/B _07175_/A _07175_/B _07303_/B vssd1 vssd1 vccd1 vccd1 _07325_/B
+ sky130_fd_sc_hd__o31a_4
XANTENNA_fanout137_A _07057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10271__B1 _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07254_ reg1_val[16] _07087_/B _07165_/A vssd1 vssd1 vccd1 vccd1 _07255_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08415__A _08415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08134__B _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ reg1_val[13] _07165_/B _07105_/A vssd1 vssd1 vccd1 vccd1 _07189_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11771__B1 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11523__B1 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09826_ _06868_/C _09825_/X _12277_/B1 vssd1 vssd1 vccd1 vccd1 _09826_/Y sky130_fd_sc_hd__a21oi_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06969_ _07087_/B _12658_/B _07105_/A vssd1 vssd1 vccd1 vccd1 _07316_/B sky130_fd_sc_hd__o21ai_2
X_09757_ _09757_/A _09757_/B _09757_/C vssd1 vssd1 vccd1 vccd1 _09758_/B sky130_fd_sc_hd__and3_1
XANTENNA__12079__B2 _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08708_ _07998_/A _07998_/B _07996_/X vssd1 vssd1 vccd1 vccd1 _08713_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_68_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06950__B1 _07001_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09688_ _09683_/X _09686_/X _09687_/Y vssd1 vssd1 vccd1 vccd1 _09688_/X sky130_fd_sc_hd__a21o_1
X_08639_ _08641_/A _08641_/B vssd1 vssd1 vccd1 vccd1 _08639_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11650_ reg1_val[20] curr_PC[20] vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout30 _07006_/Y vssd1 vssd1 vccd1 vccd1 fanout30/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_126_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11581_ _09205_/B _11569_/X _11580_/X _11563_/X vssd1 vssd1 vccd1 vccd1 _11581_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_64_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout52 _08134_/B vssd1 vssd1 vccd1 vccd1 fanout52/X sky130_fd_sc_hd__buf_8
Xfanout41 _12255_/B vssd1 vssd1 vccd1 vccd1 _12200_/A sky130_fd_sc_hd__buf_8
Xfanout63 _07119_/Y vssd1 vssd1 vccd1 vccd1 _12772_/A sky130_fd_sc_hd__buf_8
XFILLER_0_37_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout74 _12768_/A vssd1 vssd1 vccd1 vccd1 _11704_/A sky130_fd_sc_hd__buf_6
XFILLER_0_36_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10601_ _10602_/A _10602_/B vssd1 vssd1 vccd1 vccd1 _10601_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout96 _08672_/A vssd1 vssd1 vccd1 vccd1 _08217_/B sky130_fd_sc_hd__buf_8
Xfanout85 _09580_/A vssd1 vssd1 vccd1 vccd1 _10559_/A sky130_fd_sc_hd__buf_6
X_13320_ instruction[12] vssd1 vssd1 vccd1 vccd1 loadstore_dest[1] sky130_fd_sc_hd__buf_12
X_10532_ _10408_/Y _10411_/B _10416_/A vssd1 vssd1 vccd1 vccd1 _10533_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13251_ _13318_/CLK hold85/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08758__A1 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10463_ _10463_/A _10463_/B vssd1 vssd1 vccd1 vccd1 _10464_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10014__B1 _11222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13182_ hold163/X _12721_/C _13179_/A vssd1 vssd1 vccd1 vccd1 hold164/A sky130_fd_sc_hd__o21a_1
XANTENNA__08758__B2 _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10394_ _12361_/B _09851_/B _10392_/X _11913_/B _12373_/A1 vssd1 vssd1 vccd1 vccd1
+ _10395_/C sky130_fd_sc_hd__a32o_1
XFILLER_0_60_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12202_ _12202_/A _12202_/B vssd1 vssd1 vccd1 vccd1 _12204_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12133_ _12133_/A _12133_/B vssd1 vssd1 vccd1 vccd1 _12133_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12064_ _06596_/Y _12243_/B1 _12062_/Y _06597_/X _12063_/X vssd1 vssd1 vccd1 vccd1
+ _12064_/X sky130_fd_sc_hd__o221a_1
X_11015_ _11158_/A _11015_/B vssd1 vssd1 vccd1 vccd1 _11017_/B sky130_fd_sc_hd__or2_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12966_ _07115_/B _12742_/B hold160/X vssd1 vssd1 vccd1 vccd1 _13253_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_59_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11917_ hold256/A _11915_/X _11916_/Y vssd1 vssd1 vccd1 vccd1 _11926_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08694__B1 _07119_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12897_ _13218_/Q _12955_/A2 _13168_/B1 hold248/X vssd1 vssd1 vccd1 vccd1 hold249/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07497__A1 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07497__B2 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11848_ _11972_/A _11972_/B _11972_/C _11973_/A vssd1 vssd1 vccd1 vccd1 _11848_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12547__A2_N _12538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11779_ fanout29/X fanout20/X fanout18/X fanout32/X vssd1 vssd1 vccd1 vccd1 _11780_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08990_ _08990_/A _08990_/B vssd1 vssd1 vccd1 vccd1 _09507_/B sky130_fd_sc_hd__nand2_2
X_07941_ _07941_/A _07941_/B vssd1 vssd1 vccd1 vccd1 _08019_/B sky130_fd_sc_hd__or2_4
X_07872_ _07872_/A _07872_/B _07872_/C vssd1 vssd1 vccd1 vccd1 _07935_/A sky130_fd_sc_hd__or3_2
X_06823_ reg1_val[19] _07077_/A vssd1 vssd1 vccd1 vccd1 _06823_/Y sky130_fd_sc_hd__nand2_1
X_09611_ _09612_/A _09612_/B vssd1 vssd1 vccd1 vccd1 _09736_/C sky130_fd_sc_hd__nor2_1
X_09542_ hold297/A _11820_/A _09540_/X _12290_/C1 vssd1 vssd1 vccd1 vccd1 _09542_/X
+ sky130_fd_sc_hd__a31o_1
X_06754_ reg2_val[5] _06778_/B _12284_/A vssd1 vssd1 vccd1 vccd1 _06972_/C sky130_fd_sc_hd__a21o_2
XANTENNA__11284__A2 _11183_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06685_ _06685_/A _06685_/B vssd1 vssd1 vccd1 vccd1 _06865_/C sky130_fd_sc_hd__nor2_1
XANTENNA_fanout254_A _12382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09473_ _09474_/A _09474_/B vssd1 vssd1 vccd1 vccd1 _09473_/Y sky130_fd_sc_hd__nand2b_1
X_08424_ _08588_/A _08420_/B _08461_/B _08423_/X vssd1 vssd1 vccd1 vccd1 _08433_/B
+ sky130_fd_sc_hd__o31ai_2
XANTENNA__10492__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08355_ _08695_/A _08355_/B _08355_/C vssd1 vssd1 vccd1 vccd1 _08358_/B sky130_fd_sc_hd__and3_1
XANTENNA__08437__B1 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11036__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07306_ _10180_/A _11429_/B _10559_/A vssd1 vssd1 vccd1 vccd1 _07308_/A sky130_fd_sc_hd__or3b_4
X_08286_ _08286_/A vssd1 vssd1 vccd1 vccd1 _08342_/A sky130_fd_sc_hd__inv_2
XFILLER_0_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07237_ _07237_/A _07237_/B vssd1 vssd1 vccd1 vccd1 _07274_/A sky130_fd_sc_hd__xnor2_2
X_07168_ _07168_/A _07168_/B vssd1 vssd1 vccd1 vccd1 _07168_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__10547__A1 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10547__B2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06766__A3 _12578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07099_ _07098_/A _07098_/B _10280_/A vssd1 vssd1 vccd1 vccd1 _07099_/X sky130_fd_sc_hd__mux2_2
Xfanout231 _06579_/Y vssd1 vssd1 vccd1 vccd1 _06688_/B1 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout220 _10246_/S vssd1 vssd1 vccd1 vccd1 _10247_/S sky130_fd_sc_hd__clkbuf_8
Xfanout264 _06577_/Y vssd1 vssd1 vccd1 vccd1 _06687_/A sky130_fd_sc_hd__buf_4
Xfanout253 _12556_/S vssd1 vssd1 vccd1 vccd1 _12005_/A sky130_fd_sc_hd__buf_6
Xfanout286 _06550_/X vssd1 vssd1 vccd1 vccd1 _06633_/B sky130_fd_sc_hd__buf_4
Xfanout297 _11647_/S vssd1 vssd1 vccd1 vccd1 _11738_/S sky130_fd_sc_hd__clkbuf_8
Xfanout275 _06931_/X vssd1 vssd1 vccd1 vccd1 _07105_/A sky130_fd_sc_hd__clkbuf_8
X_09809_ _09810_/A _09810_/B vssd1 vssd1 vccd1 vccd1 _09809_/X sky130_fd_sc_hd__and2_1
X_12820_ hold13/X hold288/A vssd1 vssd1 vccd1 vccd1 _12820_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_69_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12751_ _10811_/A _12980_/A2 hold62/X _13086_/A vssd1 vssd1 vccd1 vccd1 _13197_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ _12682_/A _12688_/A vssd1 vssd1 vccd1 vccd1 _12684_/A sky130_fd_sc_hd__nand2_2
X_11702_ _11614_/A _11614_/B _11613_/A vssd1 vssd1 vccd1 vccd1 _11713_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11633_ _11633_/A _11633_/B vssd1 vssd1 vccd1 vccd1 _11812_/A sky130_fd_sc_hd__and2_1
XFILLER_0_126_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06782__B _09392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11564_ reg1_val[19] curr_PC[19] vssd1 vssd1 vccd1 vccd1 _11566_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07100__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10786__A1 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10786__B2 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10515_ _09385_/C _10635_/B hold272/A vssd1 vssd1 vccd1 vccd1 _10515_/Y sky130_fd_sc_hd__a21oi_1
X_13303_ _13303_/CLK _13303_/D vssd1 vssd1 vccd1 vccd1 hold293/A sky130_fd_sc_hd__dfxtp_1
X_11495_ _10400_/S _11492_/X _11671_/C _11494_/Y vssd1 vssd1 vccd1 vccd1 dest_val[18]
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_24_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07894__A _07894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13234_ _13306_/CLK _13234_/D vssd1 vssd1 vccd1 vccd1 hold178/A sky130_fd_sc_hd__dfxtp_1
X_10446_ _10446_/A _10446_/B _10446_/C vssd1 vssd1 vccd1 vccd1 _10592_/A sky130_fd_sc_hd__or3_2
XANTENNA__11735__B1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13165_ hold242/X _13165_/A2 _13164_/X _13168_/A2 vssd1 vssd1 vccd1 vccd1 _13166_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11204__A1_N _07178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap99_A _07168_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10377_ reg1_val[8] _10377_/B vssd1 vssd1 vccd1 vccd1 _10377_/Y sky130_fd_sc_hd__nor2_1
X_13096_ _13166_/A hold259/X vssd1 vssd1 vccd1 vccd1 _13296_/D sky130_fd_sc_hd__and2_1
X_12116_ _12114_/X _12115_/Y _12112_/X vssd1 vssd1 vccd1 vccd1 _12116_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12047_ _11820_/A _09079_/B _09079_/A vssd1 vssd1 vccd1 vccd1 _12047_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09614__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06957__B _06965_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12949_ hold213/X _12955_/A2 _13168_/B1 hold165/X vssd1 vssd1 vccd1 vccd1 hold214/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07134__A _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08140_ _08857_/A _08140_/B vssd1 vssd1 vccd1 vccd1 _08144_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_7_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08071_ _08071_/A _08071_/B vssd1 vssd1 vccd1 vccd1 _08080_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_71_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07642__B2 _09925_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07642__A1 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07022_ _06684_/B _07168_/A _07051_/A _07051_/B _07303_/B vssd1 vssd1 vccd1 vccd1
+ _07077_/B sky130_fd_sc_hd__o41a_4
XANTENNA__06609__A2_N _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07945__A2 _09295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08973_ _08974_/A _08974_/B vssd1 vssd1 vccd1 vccd1 _08973_/X sky130_fd_sc_hd__and2_1
X_07924_ _07924_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _08056_/A sky130_fd_sc_hd__xnor2_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__B1 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ _07855_/A _07855_/B vssd1 vssd1 vccd1 vccd1 _07932_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_127_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07786_ _07790_/A vssd1 vssd1 vccd1 vccd1 _07786_/Y sky130_fd_sc_hd__inv_2
X_06806_ _10621_/A _06804_/X _06805_/X vssd1 vssd1 vccd1 vccd1 _06806_/Y sky130_fd_sc_hd__a21oi_1
X_06737_ reg1_val[8] _07015_/B vssd1 vssd1 vccd1 vccd1 _06739_/A sky130_fd_sc_hd__or2_1
XANTENNA__07044__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09525_ _10112_/B _09524_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09525_/X sky130_fd_sc_hd__mux2_1
X_06668_ _06668_/A _06668_/B vssd1 vssd1 vccd1 vccd1 _06865_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_78_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09456_ fanout77/X fanout98/X fanout56/X fanout75/X vssd1 vssd1 vccd1 vccd1 _09457_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08407_ _08407_/A _08407_/B vssd1 vssd1 vccd1 vccd1 _08427_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06599_ instruction[34] _06633_/B vssd1 vssd1 vccd1 vccd1 _12603_/B sky130_fd_sc_hd__and2_4
X_09387_ _11400_/A _09385_/X _09386_/Y _11099_/B reg1_val[1] vssd1 vssd1 vccd1 vccd1
+ _09387_/X sky130_fd_sc_hd__o32a_1
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08338_ _08339_/A _08339_/B vssd1 vssd1 vccd1 vccd1 _08338_/X sky130_fd_sc_hd__or2_1
XANTENNA__12757__A2 _12781_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08269_ _08328_/A _08328_/B vssd1 vssd1 vccd1 vccd1 _08329_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07633__A1 _07260_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07633__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11013__B _11014_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11280_ _10855_/B _11279_/Y _11638_/A vssd1 vssd1 vccd1 vccd1 _11281_/B sky130_fd_sc_hd__o21bai_1
X_10300_ fanout37/X _07553_/A _10927_/A fanout35/X vssd1 vssd1 vccd1 vccd1 _10301_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10231_ _09661_/X _09662_/X _10230_/C vssd1 vssd1 vccd1 vccd1 _10231_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07397__B1 _07157_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09925__A3 _07322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07219__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10162_ _07389_/B fanout81/X _09295_/B fanout26/X vssd1 vssd1 vccd1 vccd1 _10163_/B
+ sky130_fd_sc_hd__o22a_1
X_10093_ _10094_/A _10094_/B vssd1 vssd1 vccd1 vccd1 _10093_/X sky130_fd_sc_hd__and2_1
XFILLER_0_89_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11496__A2 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12803_ hold277/X hold5/X vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__11248__A2 _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12734_ _12734_/A _12788_/B vssd1 vssd1 vccd1 vccd1 _12734_/Y sky130_fd_sc_hd__nand2_1
X_10995_ _10968_/X _10969_/Y _10973_/X _10994_/X vssd1 vssd1 vccd1 vccd1 _10995_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12996__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07321__B1 _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ reg1_val[20] _12714_/A _12661_/A vssd1 vssd1 vccd1 vccd1 _12666_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_37_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12596_ _12595_/A _12592_/Y _12594_/B vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__o21a_2
X_11616_ _11616_/A _11616_/B vssd1 vssd1 vccd1 vccd1 _11620_/A sky130_fd_sc_hd__or2_1
XANTENNA__09613__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11547_ _11547_/A _11547_/B _11547_/C vssd1 vssd1 vccd1 vccd1 _11548_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_25_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11478_ _11478_/A _11478_/B vssd1 vssd1 vccd1 vccd1 _11478_/X sky130_fd_sc_hd__xor2_1
XANTENNA__08513__A _09620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13217_ _13312_/CLK _13217_/D vssd1 vssd1 vccd1 vccd1 hold211/A sky130_fd_sc_hd__dfxtp_1
X_10429_ _10429_/A _10429_/B vssd1 vssd1 vccd1 vccd1 _10430_/B sky130_fd_sc_hd__or2_1
X_13148_ _13148_/A _13148_/B vssd1 vssd1 vccd1 vccd1 _13149_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06595__A2_N _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07129__A _07153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ hold291/A _13078_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13079_/X sky130_fd_sc_hd__mux2_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06968__A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06687__B _12563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07640_ _08906_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08907_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07571_ _08825_/A2 _07278_/B fanout7/X _08588_/A vssd1 vssd1 vccd1 vccd1 _07572_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__07560__B1 _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11239__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09310_ _09310_/A _09310_/B vssd1 vssd1 vccd1 vccd1 _09312_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09852__A2 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07863__A1 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07863__B2 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09241_ _09240_/B _09241_/B vssd1 vssd1 vccd1 vccd1 _09242_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_28_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12739__A2 _12980_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09172_ reg1_val[22] reg1_val[9] _09172_/S vssd1 vssd1 vccd1 vccd1 _09172_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11114__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08123_ _08123_/A _08123_/B vssd1 vssd1 vccd1 vccd1 _08158_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_44_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08054_ _07935_/B _07908_/B _07908_/C vssd1 vssd1 vccd1 vccd1 _08055_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_114_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout217_A _09392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08423__A _10453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07005_ _12019_/A _11853_/A _07005_/C vssd1 vssd1 vccd1 vccd1 _07005_/Y sky130_fd_sc_hd__nand3b_1
XANTENNA__13164__A2 fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07128__A_N _07153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__B2 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _08957_/B _08957_/A vssd1 vssd1 vccd1 vccd1 _08956_/Y sky130_fd_sc_hd__nand2b_1
X_07907_ _07907_/A _07907_/B vssd1 vssd1 vccd1 vccd1 _07908_/C sky130_fd_sc_hd__xor2_1
X_08887_ _08761_/A _08761_/B _08834_/B _08832_/Y vssd1 vssd1 vccd1 vccd1 _08894_/A
+ sky130_fd_sc_hd__o31a_1
XANTENNA__06597__B _07157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ _07786_/Y _07802_/A _07840_/B vssd1 vssd1 vccd1 vccd1 _07838_/X sky130_fd_sc_hd__a21o_1
X_07769_ _08443_/A _07769_/B vssd1 vssd1 vccd1 vccd1 _07770_/B sky130_fd_sc_hd__xor2_4
X_09508_ _07705_/X _09329_/X _09330_/X vssd1 vssd1 vccd1 vccd1 _09508_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_2_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout32_A _07000_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10780_ _07553_/A _07278_/B fanout6/X _10927_/A vssd1 vssd1 vccd1 vccd1 _10781_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09439_ _09303_/B _09306_/B _09301_/X vssd1 vssd1 vccd1 vccd1 _09442_/A sky130_fd_sc_hd__a21oi_1
X_12450_ _12450_/A _12450_/B _12450_/C vssd1 vssd1 vccd1 vccd1 _12451_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_93_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11401_ hold207/A _11480_/C _12187_/A1 vssd1 vssd1 vccd1 vccd1 _11402_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12381_ _12387_/A _12381_/B vssd1 vssd1 vccd1 vccd1 new_PC[0] sky130_fd_sc_hd__and2_4
XFILLER_0_62_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_80 _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07082__A2 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11332_ _12022_/A _11332_/B vssd1 vssd1 vccd1 vccd1 _11336_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13155__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11263_ _11261_/X _11263_/B vssd1 vssd1 vccd1 vccd1 _11264_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_120_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13002_ _06987_/B _13020_/B2 hold127/X vssd1 vssd1 vccd1 vccd1 _13271_/D sky130_fd_sc_hd__o21a_1
X_11194_ _10247_/X _10249_/X _11194_/S vssd1 vssd1 vccd1 vccd1 _11194_/X sky130_fd_sc_hd__mux2_1
X_10214_ _10212_/A _10212_/B _10215_/B vssd1 vssd1 vccd1 vccd1 _10214_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10374__C1 _12228_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11694__A _11695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ _10551_/B _10145_/B vssd1 vssd1 vccd1 vccd1 _10147_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10913__B2 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10913__A1 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10076_ _10074_/Y _10076_/B vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_69_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10978_ _10978_/A _10978_/B vssd1 vssd1 vccd1 vccd1 _10978_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12717_ hold154/X hold176/X hold171/X hold137/X vssd1 vssd1 vccd1 vccd1 _12719_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_85_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10249__S _10249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12648_ reg1_val[18] _12714_/A vssd1 vssd1 vccd1 vccd1 _12648_/X sky130_fd_sc_hd__and2_1
XFILLER_0_108_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12579_ _12577_/Y _12579_/B vssd1 vssd1 vccd1 vccd1 _12580_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13146__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08810_ _08794_/A _08794_/B _08795_/Y vssd1 vssd1 vccd1 vccd1 _08881_/A sky130_fd_sc_hd__o21ai_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _09600_/A _09775_/A _09606_/B _09604_/X vssd1 vssd1 vccd1 vccd1 _09792_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _08741_/A _08741_/B vssd1 vssd1 vccd1 vccd1 _08752_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_84_54 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08325__A2 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08672_ _08672_/A _08672_/B vssd1 vssd1 vccd1 vccd1 _08674_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_84_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07306__B _11429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07623_ _07703_/A _07703_/B vssd1 vssd1 vccd1 vccd1 _07623_/X sky130_fd_sc_hd__and2_1
XANTENNA_fanout167_A _07110_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07554_ _07308_/A _07308_/B _10927_/A vssd1 vssd1 vccd1 vccd1 _07555_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_91_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12290__C1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07322__A _07322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07485_ _07485_/A _07485_/B vssd1 vssd1 vccd1 vccd1 _07581_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09224_ _09559_/A wire3/X _12131_/A vssd1 vssd1 vccd1 vccd1 _09224_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_106_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11396__A1 _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__B2 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09155_ reg1_val[29] reg1_val[2] _09158_/S vssd1 vssd1 vccd1 vccd1 _09155_/X sky130_fd_sc_hd__mux2_1
X_08106_ _08106_/A _08106_/B vssd1 vssd1 vccd1 vccd1 _08108_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09086_ _09103_/A _09086_/B _09086_/C vssd1 vssd1 vccd1 vccd1 _09088_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08037_ _08855_/A _08037_/B vssd1 vssd1 vccd1 vccd1 _08043_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__13137__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07992__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09988_ _09850_/A _09847_/Y _09849_/B vssd1 vssd1 vccd1 vccd1 _09992_/A sky130_fd_sc_hd__o21a_1
X_08939_ _08925_/A _08925_/B _08926_/Y vssd1 vssd1 vccd1 vccd1 _08960_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_98_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11950_ _11950_/A _11950_/B vssd1 vssd1 vccd1 vccd1 _11952_/C sky130_fd_sc_hd__xnor2_1
X_10901_ fanout32/X _11704_/A _11688_/A fanout29/X vssd1 vssd1 vccd1 vccd1 _10902_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12549__S _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11881_ _11881_/A _11881_/B vssd1 vssd1 vccd1 vccd1 _11883_/B sky130_fd_sc_hd__xnor2_1
X_10832_ _10832_/A _10832_/B _10832_/C vssd1 vssd1 vccd1 vccd1 _10833_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_94_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10763_ _06722_/B wire201/X _10762_/X vssd1 vssd1 vccd1 vccd1 _10763_/Y sky130_fd_sc_hd__a21boi_1
X_12502_ _12515_/B _12516_/B _12515_/A vssd1 vssd1 vccd1 vccd1 _12509_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10694_ _10694_/A _12255_/B _10695_/A vssd1 vssd1 vccd1 vccd1 _10694_/X sky130_fd_sc_hd__and3_1
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12433_ _12598_/B _12433_/B vssd1 vssd1 vccd1 vccd1 _12434_/B sky130_fd_sc_hd__or2_1
XFILLER_0_50_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12364_ hold231/A _12332_/C _12332_/B vssd1 vssd1 vccd1 vccd1 _12364_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_50_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13128__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11315_ _11313_/Y _11493_/B _10400_/S vssd1 vssd1 vccd1 vccd1 _11315_/Y sky130_fd_sc_hd__o21ai_1
X_12295_ _12295_/A _12295_/B _12295_/C vssd1 vssd1 vccd1 vccd1 _12295_/X sky130_fd_sc_hd__and3_1
XFILLER_0_120_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11246_ _11499_/A _11246_/B vssd1 vssd1 vccd1 vccd1 _11250_/A sky130_fd_sc_hd__xnor2_1
X_11177_ _10734_/B _11174_/Y _11176_/Y vssd1 vssd1 vccd1 vccd1 _11177_/X sky130_fd_sc_hd__o21a_1
X_10128_ _09992_/A _09989_/Y _09991_/B vssd1 vssd1 vccd1 vccd1 _10132_/A sky130_fd_sc_hd__o21a_1
XANTENNA__07407__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06949__C _09392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07126__B _07126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10059_ _10061_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _10194_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09622__A _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12459__S _12487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06965__B _11780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09268__B1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11075__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07270_ _07270_/A _07270_/B vssd1 vssd1 vccd1 vccd1 _07272_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06981__A _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13119__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold103 hold103/A vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 hold114/A vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 hold158/A vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 hold147/A vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _09911_/A _10037_/A _09911_/C vssd1 vssd1 vccd1 vccd1 _10037_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10008__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold169 hold169/A vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09338__A4 _09620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09842_ hold288/A _09842_/B _10122_/C vssd1 vssd1 vccd1 vccd1 _09842_/X sky130_fd_sc_hd__and3_1
XANTENNA__10889__B1 _10886_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09743__A1 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09743__B2 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08420__B _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07317__A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09773_ _08589_/A _09622_/B _09620_/Y vssd1 vssd1 vccd1 vccd1 _09777_/A sky130_fd_sc_hd__a21oi_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08724_ _08836_/A _08724_/B vssd1 vssd1 vccd1 vccd1 _08728_/A sky130_fd_sc_hd__xnor2_1
X_06985_ _06986_/A _06986_/B vssd1 vssd1 vccd1 vccd1 _06985_/X sky130_fd_sc_hd__xor2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _07958_/A _07958_/B _07954_/X vssd1 vssd1 vccd1 vccd1 _08657_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_96_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10678__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13055__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _08825_/A2 _08758_/A2 _09476_/A _06864_/A vssd1 vssd1 vccd1 vccd1 _08587_/B
+ sky130_fd_sc_hd__o22a_1
X_07606_ _07604_/A _07597_/Y _07605_/X vssd1 vssd1 vccd1 vccd1 _07617_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__09259__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07052__A _07068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07537_ _07538_/A _07538_/B vssd1 vssd1 vccd1 vccd1 _07537_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07987__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06891__A _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07468_ _10144_/B2 _08680_/B fanout30/X _10064_/B2 vssd1 vssd1 vccd1 vccd1 _07469_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07399_ _07396_/A _07396_/B _07396_/C vssd1 vssd1 vccd1 vccd1 _07400_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_63_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09207_ _09158_/X _09213_/B _09359_/S vssd1 vssd1 vccd1 vccd1 _09207_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09138_ reg1_val[12] reg1_val[19] _09172_/S vssd1 vssd1 vccd1 vccd1 _09138_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09069_ _09069_/A _09073_/C vssd1 vssd1 vccd1 vccd1 _09069_/X sky130_fd_sc_hd__or2_1
X_11100_ _07192_/A _06928_/X _10638_/B _06702_/X _11099_/Y vssd1 vssd1 vccd1 vccd1
+ _11100_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_32_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12080_ _12081_/A _12081_/B vssd1 vssd1 vccd1 vccd1 _12152_/A sky130_fd_sc_hd__or2_1
XFILLER_0_12_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12133__A _12133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11031_ fanout37/X _11688_/A fanout70/X fanout35/X vssd1 vssd1 vccd1 vccd1 _11032_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07745__B1 _08774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ _07172_/B _12744_/B hold162/X vssd1 vssd1 vccd1 vccd1 _13261_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_99_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11933_ _11933_/A _12349_/A vssd1 vssd1 vccd1 vccd1 _11933_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08170__B1 _07181_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11864_ _11864_/A _11864_/B vssd1 vssd1 vccd1 vccd1 _11883_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10815_ _10815_/A _10815_/B vssd1 vssd1 vccd1 vccd1 _10816_/B sky130_fd_sc_hd__or2_1
XFILLER_0_95_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11795_ _11795_/A _11795_/B vssd1 vssd1 vccd1 vccd1 _11797_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10746_ reg1_val[11] curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10747_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_55_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10677_ _10677_/A _10677_/B vssd1 vssd1 vccd1 vccd1 _10678_/C sky130_fd_sc_hd__or2_1
XFILLER_0_40_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08225__A1 _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12416_ _12422_/B _12416_/B vssd1 vssd1 vccd1 vccd1 new_PC[5] sky130_fd_sc_hd__and2_4
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12021__A2 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08225__B2 _08692_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08776__A2 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12347_ _12307_/A _12305_/Y _12301_/X vssd1 vssd1 vccd1 vccd1 _12348_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_11_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12278_ _12278_/A _12278_/B vssd1 vssd1 vccd1 vccd1 _12279_/B sky130_fd_sc_hd__and2_1
XFILLER_0_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11229_ _11230_/B _11229_/B vssd1 vssd1 vccd1 vccd1 _11354_/A sky130_fd_sc_hd__and2b_1
XANTENNA__10335__A2 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ _06768_/Y _06771_/B vssd1 vssd1 vccd1 vccd1 _06770_/X sky130_fd_sc_hd__and2b_1
XANTENNA__12697__B _12697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10099__A1 _09511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11093__S _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08440_ _09621_/A _08440_/B vssd1 vssd1 vccd1 vccd1 _08445_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__13037__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08371_ _08371_/A _08371_/B vssd1 vssd1 vccd1 vccd1 _08372_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07322_ _07322_/A _07322_/B vssd1 vssd1 vccd1 vccd1 _07322_/X sky130_fd_sc_hd__or2_2
XFILLER_0_46_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07253_ reg1_val[13] reg1_val[14] reg1_val[15] _07165_/B _07165_/A vssd1 vssd1 vccd1
+ vccd1 _07257_/B sky130_fd_sc_hd__o41a_2
XFILLER_0_45_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07184_ _08733_/A _07184_/B vssd1 vssd1 vccd1 vccd1 _07631_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11771__A1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11771__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09825_ _06792_/Y _09824_/X _12322_/S vssd1 vssd1 vccd1 vccd1 _09825_/X sky130_fd_sc_hd__mux2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11523__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11523__B2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09756_ _09757_/B _09757_/C _09757_/A vssd1 vssd1 vccd1 vccd1 _09758_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__12079__A2 _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ _10169_/A _06968_/B vssd1 vssd1 vccd1 vccd1 _06993_/A sky130_fd_sc_hd__xnor2_1
X_08707_ _08008_/A _08008_/B _08006_/Y vssd1 vssd1 vccd1 vccd1 _08715_/A sky130_fd_sc_hd__a21o_1
X_09687_ _09683_/X _09686_/X _12361_/B vssd1 vssd1 vccd1 vccd1 _09687_/Y sky130_fd_sc_hd__o21ai_1
X_08638_ _08638_/A _08638_/B vssd1 vssd1 vccd1 vccd1 _09076_/A sky130_fd_sc_hd__xnor2_4
X_06899_ instruction[11] _06904_/B vssd1 vssd1 vccd1 vccd1 dest_idx[0] sky130_fd_sc_hd__and2_4
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12236__C1 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ _08568_/B _08568_/C _08568_/A vssd1 vssd1 vccd1 vccd1 _08605_/B sky130_fd_sc_hd__o21ai_1
Xfanout20 _12784_/A vssd1 vssd1 vccd1 vccd1 fanout20/X sky130_fd_sc_hd__clkbuf_8
Xfanout31 fanout32/X vssd1 vssd1 vccd1 vccd1 _08680_/B sky130_fd_sc_hd__buf_6
X_11580_ _11574_/Y _11575_/X _11579_/X _11572_/X vssd1 vssd1 vccd1 vccd1 _11580_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout53 _07260_/Y vssd1 vssd1 vccd1 vccd1 _08134_/B sky130_fd_sc_hd__buf_8
Xfanout64 _12774_/A vssd1 vssd1 vccd1 vccd1 _11935_/A sky130_fd_sc_hd__buf_6
X_10600_ _10600_/A _10600_/B vssd1 vssd1 vccd1 vccd1 _10602_/B sky130_fd_sc_hd__xnor2_4
Xfanout42 _11147_/B vssd1 vssd1 vccd1 vccd1 _12255_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout75 _12768_/A vssd1 vssd1 vccd1 vccd1 fanout75/X sky130_fd_sc_hd__clkbuf_4
Xfanout86 _11499_/A vssd1 vssd1 vccd1 vccd1 _09580_/A sky130_fd_sc_hd__buf_12
XANTENNA__07510__A _10180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10531_ _10705_/A _10531_/B vssd1 vssd1 vccd1 vccd1 _10533_/A sky130_fd_sc_hd__xnor2_4
X_13250_ _13289_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11032__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10462_ _10462_/A _10462_/B vssd1 vssd1 vccd1 vccd1 _10463_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12201_ _12202_/A _12202_/B vssd1 vssd1 vccd1 vccd1 _12201_/Y sky130_fd_sc_hd__nand2_1
X_13181_ hold31/X _12719_/B _13180_/X _13179_/A vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__o211a_1
XFILLER_0_103_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11211__B1 _06898_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11762__A1 _07052_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08758__A2 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10393_ _10251_/S _10250_/X _09214_/A vssd1 vssd1 vccd1 vccd1 _11913_/B sky130_fd_sc_hd__o21a_1
XANTENNA__10014__B2 _09294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12132_ _12133_/A _12133_/B vssd1 vssd1 vccd1 vccd1 _12132_/Y sky130_fd_sc_hd__nand2_1
X_12063_ _07157_/A _12250_/B _10377_/B reg1_val[25] vssd1 vssd1 vccd1 vccd1 _12063_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11014_ _11014_/A _11014_/B vssd1 vssd1 vccd1 vccd1 _11015_/B sky130_fd_sc_hd__and2_1
XFILLER_0_19_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08391__B1 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12965_ hold157/X _12723_/A _13170_/B hold159/X _13066_/A vssd1 vssd1 vccd1 vccd1
+ hold160/A sky130_fd_sc_hd__o221a_1
XFILLER_0_35_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11916_ hold256/A _11915_/X _09200_/X vssd1 vssd1 vccd1 vccd1 _11916_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09340__C1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08694__A1 _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12896_ _13169_/A hold212/X vssd1 vssd1 vccd1 vccd1 _13218_/D sky130_fd_sc_hd__and2_1
XANTENNA__08694__B2 _07869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07497__A2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11847_ _10400_/S _11844_/X _11846_/Y vssd1 vssd1 vccd1 vccd1 dest_val[22] sky130_fd_sc_hd__o21ai_4
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11778_ _11778_/A _11778_/B vssd1 vssd1 vccd1 vccd1 _11786_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10729_ _10483_/X _10604_/X _10605_/X vssd1 vssd1 vccd1 vccd1 _10729_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10781__A _12255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_7_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13309_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07940_ _08021_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _07941_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_76_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07709__B1 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07871_ _09621_/A _07871_/B _07871_/C vssd1 vssd1 vccd1 vccd1 _07872_/C sky130_fd_sc_hd__and3_1
X_06822_ _06677_/Y _06820_/Y _06821_/X vssd1 vssd1 vccd1 vccd1 _06822_/Y sky130_fd_sc_hd__a21oi_2
X_09610_ _09610_/A _09610_/B vssd1 vssd1 vccd1 vccd1 _09612_/B sky130_fd_sc_hd__xnor2_1
X_09541_ _11820_/A _09540_/X hold297/A vssd1 vssd1 vccd1 vccd1 _09541_/Y sky130_fd_sc_hd__a21oi_1
X_06753_ reg2_val[5] _06778_/B _12284_/A vssd1 vssd1 vccd1 vccd1 _06795_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06684_ reg1_val[17] _06684_/B vssd1 vssd1 vccd1 vccd1 _06685_/B sky130_fd_sc_hd__and2_1
XFILLER_0_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09472_ _09472_/A _09472_/B vssd1 vssd1 vccd1 vccd1 _09474_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_93_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08423_ _10453_/A _08461_/A vssd1 vssd1 vccd1 vccd1 _08423_/X sky130_fd_sc_hd__or2_1
XFILLER_0_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08354_ _08355_/B _08355_/C _08695_/A vssd1 vssd1 vccd1 vccd1 _08358_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08437__B2 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08437__A1 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout247_A _07869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07305_ _08305_/B _08305_/C vssd1 vssd1 vccd1 vccd1 _07305_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08285_ _08285_/A _08285_/B vssd1 vssd1 vccd1 vccd1 _08286_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07236_ _09452_/A _07236_/B vssd1 vssd1 vccd1 vccd1 _07237_/B sky130_fd_sc_hd__xnor2_2
X_07167_ _07167_/A _07168_/B vssd1 vssd1 vccd1 vccd1 _07167_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12382__S _12382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12941__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10547__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07098_ _07098_/A _07098_/B vssd1 vssd1 vccd1 vccd1 _07098_/Y sky130_fd_sc_hd__nand2_4
Xfanout232 _09384_/X vssd1 vssd1 vccd1 vccd1 _12119_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_100_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout221 _07279_/A vssd1 vssd1 vccd1 vccd1 _10246_/S sky130_fd_sc_hd__clkbuf_4
Xfanout210 _06917_/Y vssd1 vssd1 vccd1 vccd1 _09851_/B sky130_fd_sc_hd__buf_4
Xfanout265 _12723_/A vssd1 vssd1 vccd1 vccd1 _13013_/A2 sky130_fd_sc_hd__buf_4
XANTENNA__07176__A1 _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout254 _12382_/S vssd1 vssd1 vccd1 vccd1 _12556_/S sky130_fd_sc_hd__buf_6
Xfanout243 _09173_/S vssd1 vssd1 vccd1 vccd1 _09172_/S sky130_fd_sc_hd__clkbuf_8
Xfanout276 _12557_/A vssd1 vssd1 vccd1 vccd1 _12551_/A sky130_fd_sc_hd__buf_6
Xfanout287 _13169_/A vssd1 vssd1 vccd1 vccd1 _12946_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__12411__A _12583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout298 _11647_/S vssd1 vssd1 vccd1 vccd1 _12322_/S sky130_fd_sc_hd__clkbuf_8
X_09808_ _09808_/A _09808_/B vssd1 vssd1 vccd1 vccd1 _09810_/B sky130_fd_sc_hd__xnor2_4
X_09739_ _10452_/B2 _10677_/A fanout58/X _10527_/A vssd1 vssd1 vccd1 vccd1 _09740_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout62_A _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11027__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12750_ hold61/X _12788_/B vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__or2_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12681_/A _12681_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[24] sky130_fd_sc_hd__xnor2_4
X_11701_ _11701_/A _11701_/B vssd1 vssd1 vccd1 vccd1 _11715_/A sky130_fd_sc_hd__xnor2_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11632_/A _11632_/B _11632_/C vssd1 vssd1 vccd1 vccd1 _11633_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_92_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09625__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13302_ _13303_/CLK _13302_/D vssd1 vssd1 vccd1 vccd1 hold252/A sky130_fd_sc_hd__dfxtp_1
X_11563_ _06865_/A _11561_/X _11562_/Y vssd1 vssd1 vccd1 vccd1 _11563_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07100__A1 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07100__B2 _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10786__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10514_ hold268/A hold292/A _10514_/C vssd1 vssd1 vccd1 vccd1 _10635_/B sky130_fd_sc_hd__or3_1
X_11494_ curr_PC[18] _11493_/B _10400_/S vssd1 vssd1 vccd1 vccd1 _11494_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_122_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13233_ _13312_/CLK _13233_/D vssd1 vssd1 vccd1 vccd1 hold207/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11697__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10445_ _10445_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _10446_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13164_ _12891_/C fanout1/X _13162_/Y _13163_/Y vssd1 vssd1 vccd1 vccd1 _13164_/X
+ sky130_fd_sc_hd__a31o_1
X_10376_ hold187/A _10376_/B vssd1 vssd1 vccd1 vccd1 _10376_/Y sky130_fd_sc_hd__xnor2_1
X_12115_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12115_/Y sky130_fd_sc_hd__nand2_1
X_13095_ hold258/X _13151_/A2 _13094_/X _13146_/B2 vssd1 vssd1 vccd1 vccd1 hold259/A
+ sky130_fd_sc_hd__a22o_1
X_12046_ _12045_/A _12045_/B _12045_/Y _12277_/B1 vssd1 vssd1 vccd1 vccd1 _12046_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12948_ _13169_/A hold184/X vssd1 vssd1 vccd1 vccd1 hold185/A sky130_fd_sc_hd__and2_1
XANTENNA__09864__B1 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12879_ hold17/X hold262/X vssd1 vssd1 vccd1 vccd1 _13139_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_118_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08070_ _08070_/A _08070_/B vssd1 vssd1 vccd1 vccd1 _08118_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07642__A2 _07034_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07021_ _07175_/D _07021_/B vssd1 vssd1 vccd1 vccd1 _07051_/B sky130_fd_sc_hd__or2_1
XFILLER_0_3_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11400__A _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12923__B1 _13151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09077__A _09077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ _08972_/A _08972_/B vssd1 vssd1 vccd1 vccd1 _08974_/B sky130_fd_sc_hd__xnor2_2
X_07923_ _07924_/A _07924_/B vssd1 vssd1 vccd1 vccd1 _07923_/Y sky130_fd_sc_hd__nand2b_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07158__A1 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07854_ _07855_/B _07855_/A vssd1 vssd1 vccd1 vccd1 _07854_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09552__C1 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07158__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06805_ reg1_val[10] _07318_/A vssd1 vssd1 vccd1 vccd1 _06805_/X sky130_fd_sc_hd__and2_1
XANTENNA__10162__B1 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07785_ _07785_/A _07785_/B _07785_/C vssd1 vssd1 vccd1 vccd1 _07790_/A sky130_fd_sc_hd__and3_1
X_06736_ _06783_/A _06649_/A _12603_/B _06735_/X vssd1 vssd1 vccd1 vccd1 _07015_/B
+ sky130_fd_sc_hd__a31o_4
XANTENNA__07044__B _07046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09524_ _09143_/X _09164_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09524_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09855__B1 _12382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06667_ reg1_val[19] _07077_/A vssd1 vssd1 vccd1 vccd1 _06668_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_66_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09455_ _09596_/D _09455_/B vssd1 vssd1 vccd1 vccd1 _09475_/A sky130_fd_sc_hd__nor2_1
X_08406_ _08406_/A _08406_/B vssd1 vssd1 vccd1 vccd1 _08427_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_47_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09386_ hold240/A _09385_/C hold279/A vssd1 vssd1 vccd1 vccd1 _09386_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06598_ reg1_val[25] _07157_/A vssd1 vssd1 vccd1 vccd1 _12045_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09607__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08337_ _08341_/A _08341_/B _08300_/Y vssd1 vssd1 vccd1 vccd1 _08339_/B sky130_fd_sc_hd__a21oi_2
X_08268_ _08777_/A _08268_/B vssd1 vssd1 vccd1 vccd1 _08328_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07633__A2 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ _08595_/A _07219_/B vssd1 vssd1 vccd1 vccd1 _07221_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08199_ _08199_/A _08199_/B vssd1 vssd1 vccd1 vccd1 _08201_/B sky130_fd_sc_hd__xnor2_1
X_10230_ _10230_/A _10230_/B _10230_/C vssd1 vssd1 vccd1 vccd1 _10230_/X sky130_fd_sc_hd__or3_1
XFILLER_0_14_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07397__A1 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07397__B2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10161_ _10161_/A _10161_/B vssd1 vssd1 vccd1 vccd1 _10174_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_100_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10092_ _10094_/A _10094_/B vssd1 vssd1 vccd1 vccd1 _10092_/X sky130_fd_sc_hd__or2_1
XANTENNA__08346__B1 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12141__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12802_ hold86/X hold252/X vssd1 vssd1 vccd1 vccd1 _12802_/X sky130_fd_sc_hd__and2b_1
X_10994_ _09184_/X _10981_/Y _10982_/X _09205_/B _10993_/X vssd1 vssd1 vccd1 vccd1
+ _10994_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_69_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12733_ _09600_/A _12980_/A2 hold106/X _13066_/A vssd1 vssd1 vccd1 vccd1 _13188_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06793__B _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07321__A1 _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12664_ _12662_/Y _12664_/B vssd1 vssd1 vccd1 vccd1 _12678_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_53_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12595_ _12595_/A _12595_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[7] sky130_fd_sc_hd__xor2_4
X_11615_ _11529_/A _11529_/B _11515_/X vssd1 vssd1 vccd1 vccd1 _11624_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11546_ _11547_/A _11547_/B _11547_/C vssd1 vssd1 vccd1 vccd1 _11548_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_122_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13216_ _13311_/CLK _13216_/D vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__dfxtp_1
X_11477_ _11390_/A _11387_/Y _11389_/B vssd1 vssd1 vccd1 vccd1 _11478_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11220__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10428_ _10429_/A _10429_/B vssd1 vssd1 vccd1 vccd1 _10586_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13147_ _13147_/A hold265/X vssd1 vssd1 vccd1 vccd1 _13307_/D sky130_fd_sc_hd__and2_1
XFILLER_0_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _10360_/A _10360_/B vssd1 vssd1 vccd1 vccd1 _10359_/X sky130_fd_sc_hd__and2_1
X_13078_ _13078_/A _13078_/B vssd1 vssd1 vccd1 vccd1 _13078_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12029_ _12029_/A _12029_/B vssd1 vssd1 vccd1 vccd1 _12030_/B sky130_fd_sc_hd__or2_1
XANTENNA__07145__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10144__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07570_ _07573_/A _07573_/B vssd1 vssd1 vccd1 vccd1 _07570_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11644__B1 _09073_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09240_ _09241_/B _09240_/B vssd1 vssd1 vccd1 vccd1 _09242_/A sky130_fd_sc_hd__and2b_1
XANTENNA__07863__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09171_ _09169_/X _09170_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09171_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08122_ _08161_/A _08161_/B vssd1 vssd1 vccd1 vccd1 _08122_/X sky130_fd_sc_hd__and2_1
XFILLER_0_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08053_ _08053_/A _08053_/B vssd1 vssd1 vccd1 vccd1 _08055_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07004_ _07004_/A _07004_/B vssd1 vssd1 vccd1 vccd1 _07004_/X sky130_fd_sc_hd__and2_2
XFILLER_0_3_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12372__B2 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08955_ _08955_/A _08955_/B vssd1 vssd1 vccd1 vccd1 _08957_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10922__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07906_ _07935_/A _07876_/B _07874_/Y vssd1 vssd1 vccd1 vccd1 _07908_/B sky130_fd_sc_hd__a21bo_1
X_08886_ _08886_/A _08886_/B vssd1 vssd1 vccd1 vccd1 _08930_/A sky130_fd_sc_hd__nand2_4
X_07837_ _07801_/A _07801_/B _07798_/A vssd1 vssd1 vccd1 vccd1 _07840_/B sky130_fd_sc_hd__a21oi_2
X_07768_ _12766_/A _08692_/A2 _08692_/B1 fanout70/X vssd1 vssd1 vccd1 vccd1 _07769_/B
+ sky130_fd_sc_hd__o22a_2
X_06719_ reg1_val[11] _07018_/A vssd1 vssd1 vccd1 vccd1 _06722_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09507_ _09660_/A _09507_/B _09660_/B _09660_/C vssd1 vssd1 vccd1 vccd1 wire5/A sky130_fd_sc_hd__nor4_1
XFILLER_0_2_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ _08966_/A _07698_/B _07695_/Y vssd1 vssd1 vccd1 vccd1 _08983_/A sky130_fd_sc_hd__a21o_1
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout25_A fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09438_ _09438_/A _09438_/B vssd1 vssd1 vccd1 vccd1 _09444_/A sky130_fd_sc_hd__and2_1
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09369_ _09361_/X _09368_/X _11089_/A vssd1 vssd1 vccd1 vccd1 _09369_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11400_ _11400_/A _11400_/B _11400_/C vssd1 vssd1 vccd1 vccd1 _11400_/X sky130_fd_sc_hd__or3_1
XANTENNA__07067__B1 _06653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ _12560_/B _12380_/B vssd1 vssd1 vccd1 vccd1 _12381_/B sky130_fd_sc_hd__or2_1
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_70 instruction[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_81 _12588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11331_ fanout35/X _11794_/A _12772_/A fanout37/X vssd1 vssd1 vccd1 vccd1 _11332_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ _11262_/A _11262_/B _11262_/C _11262_/D vssd1 vssd1 vccd1 vccd1 _11263_/B
+ sky130_fd_sc_hd__or4_1
X_11193_ _11193_/A _11193_/B vssd1 vssd1 vccd1 vccd1 _11193_/Y sky130_fd_sc_hd__xnor2_1
X_13001_ hold107/X _13013_/A2 _13020_/A2 hold126/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold127/A sky130_fd_sc_hd__o221a_1
X_10213_ _10194_/B _10060_/X _10072_/B _10073_/B _10073_/A vssd1 vssd1 vccd1 vccd1
+ _10215_/B sky130_fd_sc_hd__a32oi_4
XFILLER_0_30_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10144_ _07278_/B _10433_/A fanout7/X _10144_/B2 vssd1 vssd1 vccd1 vccd1 _10145_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10913__A2 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11186__S _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10126__B1 wire201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10075_ _10075_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10076_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06608__A2_N _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09180__A _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09819__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10977_ reg1_val[12] curr_PC[12] _10872_/B vssd1 vssd1 vccd1 vccd1 _10978_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12716_ hold176/X hold171/X hold137/X vssd1 vssd1 vccd1 vccd1 _12716_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_57_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12647_ _12647_/A _12657_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[17] sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12578_ reg1_val[4] _12578_/B vssd1 vssd1 vccd1 vccd1 _12579_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11529_ _11529_/A _11529_/B vssd1 vssd1 vccd1 vccd1 _11542_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07230__B1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _08741_/A _08741_/B vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__or2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08671_ _08855_/A _08671_/B vssd1 vssd1 vccd1 vccd1 _08677_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07622_ _07622_/A _07622_/B vssd1 vssd1 vccd1 vccd1 _07703_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07533__A1 _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07553_ _07553_/A _09752_/B vssd1 vssd1 vccd1 vccd1 _07555_/B sky130_fd_sc_hd__or2_1
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07322__B _07322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11125__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07484_ _07485_/B _07485_/A vssd1 vssd1 vccd1 vccd1 _09316_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_118_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09223_ curr_PC[0] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09223_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09154_ reg1_val[28] reg1_val[3] _09158_/S vssd1 vssd1 vccd1 vccd1 _09154_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08105_ _08105_/A _08105_/B vssd1 vssd1 vccd1 vccd1 _08112_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09085_ _09086_/B _09086_/C vssd1 vssd1 vccd1 vccd1 _09085_/X sky130_fd_sc_hd__and2_1
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08036_ _08841_/A1 _08420_/B _08854_/B2 _08841_/B2 vssd1 vssd1 vccd1 vccd1 _08037_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09265__A _10180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09987_ _06758_/A _10638_/B _11838_/A2 _09970_/A _09986_/Y vssd1 vssd1 vccd1 vccd1
+ _09987_/X sky130_fd_sc_hd__a221o_1
X_08938_ _09098_/A _09103_/A _08937_/Y _08935_/B _08935_/A vssd1 vssd1 vccd1 vccd1
+ _09090_/B sky130_fd_sc_hd__o32a_1
XFILLER_0_99_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08869_ _08754_/A _08754_/C _08754_/B vssd1 vssd1 vccd1 vccd1 _08872_/A sky130_fd_sc_hd__a21bo_2
X_10900_ _12255_/A _10900_/B vssd1 vssd1 vccd1 vccd1 _10904_/A sky130_fd_sc_hd__xnor2_1
X_11880_ _11881_/B _11881_/A vssd1 vssd1 vccd1 vccd1 _11932_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_79_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11608__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10831_ _10832_/A _10832_/B _10832_/C vssd1 vssd1 vccd1 vccd1 _10831_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10762_ _06807_/B _11923_/A2 _11099_/B reg1_val[11] _10761_/Y vssd1 vssd1 vccd1 vccd1
+ _10762_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_67_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12501_ _12488_/B _12493_/B _12551_/A vssd1 vssd1 vccd1 vccd1 _12516_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12432_ _12598_/B _12433_/B vssd1 vssd1 vccd1 vccd1 _12443_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10693_ _10694_/A _12255_/B vssd1 vssd1 vccd1 vccd1 _10695_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12363_ _12362_/A _12362_/B _12362_/Y _09851_/B vssd1 vssd1 vccd1 vccd1 _12363_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12294_ _09158_/S _09533_/X _12293_/X vssd1 vssd1 vccd1 vccd1 _12295_/C sky130_fd_sc_hd__a21oi_1
X_11314_ curr_PC[16] curr_PC[17] _11314_/C vssd1 vssd1 vccd1 vccd1 _11493_/B sky130_fd_sc_hd__and3_1
XANTENNA__07460__B1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12336__B2 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12336__A1 _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11245_ _12301_/A _10557_/B fanout13/X fanout19/X vssd1 vssd1 vccd1 vccd1 _11246_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11176_ _10962_/Y _11374_/A _11175_/Y vssd1 vssd1 vccd1 vccd1 _11176_/Y sky130_fd_sc_hd__a21oi_1
X_10127_ _06750_/A _10638_/B _11838_/A2 _10108_/A _10126_/X vssd1 vssd1 vccd1 vccd1
+ _10127_/X sky130_fd_sc_hd__a221o_1
XANTENNA__06949__D _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10058_ _10058_/A _10147_/B vssd1 vssd1 vccd1 vccd1 _10061_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_54_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06965__C _06965_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09268__B2 _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09268__A1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11075__A1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06981__B _06987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09069__B _09073_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold104 hold104/A vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 hold126/A vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__clkbuf_2
Xhold159 hold159/A vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 hold148/A vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09910_ _09909_/A _09909_/B _09909_/C vssd1 vssd1 vccd1 vccd1 _09911_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09841_ hold246/A _09841_/B vssd1 vssd1 vccd1 vccd1 _10122_/C sky130_fd_sc_hd__or2_1
XANTENNA__07203__B1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09743__A2 _07132_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07317__B _07317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06984_ _06996_/A _06972_/C _07001_/C _07175_/A _07303_/B vssd1 vssd1 vccd1 vccd1
+ _06986_/B sky130_fd_sc_hd__o41ai_4
X_09772_ _09772_/A _12349_/B vssd1 vssd1 vccd1 vccd1 _09778_/A sky130_fd_sc_hd__or2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _08841_/A1 fanout51/X _08835_/B1 _08134_/B vssd1 vssd1 vccd1 vccd1 _08724_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11838__B1 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06962__C1 _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout277_A _12658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08654_ _08654_/A _08654_/B vssd1 vssd1 vccd1 vccd1 _08657_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_68_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13055__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08585_ _08585_/A _08585_/B vssd1 vssd1 vccd1 vccd1 _09039_/A sky130_fd_sc_hd__xnor2_2
X_07605_ _07621_/A _07621_/B vssd1 vssd1 vccd1 vccd1 _07605_/X sky130_fd_sc_hd__and2b_1
XANTENNA__09259__B2 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09259__A1 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07052__B _07052_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07536_ _10551_/B _07536_/B vssd1 vssd1 vccd1 vccd1 _07538_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09206_ _10752_/S _09213_/B vssd1 vssd1 vccd1 vccd1 _09214_/A sky130_fd_sc_hd__or2_4
XFILLER_0_8_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07467_ _10280_/A _07467_/B vssd1 vssd1 vccd1 vccd1 _07471_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10694__A _10694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07398_ _09622_/A _07398_/B vssd1 vssd1 vccd1 vccd1 _07400_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09137_ _09133_/X _09136_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09137_/X sky130_fd_sc_hd__mux2_1
X_09068_ _09068_/A _09070_/D vssd1 vssd1 vccd1 vccd1 _09073_/C sky130_fd_sc_hd__xor2_4
XFILLER_0_102_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10577__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07442__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08019_ _08019_/A _08019_/B vssd1 vssd1 vccd1 vccd1 _08641_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_102_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout92_A _07197_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11030_ _12019_/A _11030_/B vssd1 vssd1 vccd1 vccd1 _11034_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07508__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__B2 _09925_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__A1 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09723__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ hold95/X _13013_/A2 _13020_/A2 hold132/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold162/A sky130_fd_sc_hd__o221a_1
XANTENNA__08170__A1 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11932_ _11932_/A _11932_/B vssd1 vssd1 vccd1 vccd1 _11961_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08170__B2 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07243__A _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11863_ _11864_/A _11864_/B vssd1 vssd1 vccd1 vccd1 _11955_/B sky130_fd_sc_hd__and2b_1
X_10814_ _10815_/A _10815_/B vssd1 vssd1 vccd1 vccd1 _10816_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11794_ _11794_/A _12304_/B _11795_/A vssd1 vssd1 vccd1 vccd1 _11878_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10745_ reg1_val[11] curr_PC[11] vssd1 vssd1 vccd1 vccd1 _10747_/A sky130_fd_sc_hd__and2_1
XFILLER_0_55_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07681__B1 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10676_ _07139_/A _07139_/B fanout52/X vssd1 vssd1 vccd1 vccd1 _10678_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08225__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12415_ _12415_/A _12415_/B _12415_/C vssd1 vssd1 vccd1 vccd1 _12416_/B sky130_fd_sc_hd__nand3_1
X_12346_ _11973_/B _12221_/X _12319_/A _12317_/X _11973_/A vssd1 vssd1 vccd1 vccd1
+ _12353_/A sky130_fd_sc_hd__a41oi_2
XFILLER_0_121_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12277_ _12276_/A _12276_/B _12277_/B1 vssd1 vssd1 vccd1 vccd1 _12277_/X sky130_fd_sc_hd__a21o_1
X_11228_ _12019_/A _11228_/B vssd1 vssd1 vccd1 vccd1 _11229_/B sky130_fd_sc_hd__xnor2_1
X_11159_ _11159_/A _11159_/B vssd1 vssd1 vccd1 vccd1 _11160_/B sky130_fd_sc_hd__and2_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10779__A _12255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07153__A _07153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08370_ _08619_/A _08619_/B vssd1 vssd1 vccd1 vccd1 _08370_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13037__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07321_ _09580_/A _07317_/B _11604_/A vssd1 vssd1 vccd1 vccd1 _07322_/B sky130_fd_sc_hd__o21a_4
XFILLER_0_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07252_ _10894_/A _07252_/B vssd1 vssd1 vccd1 vccd1 _07266_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07183_ _11222_/A _07173_/Y _07179_/A _07182_/X vssd1 vssd1 vccd1 vccd1 _07184_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06658__A_N _07052_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11771__A2 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09824_ _06768_/Y _09694_/A _09694_/B _06771_/B vssd1 vssd1 vccd1 vccd1 _09824_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__11523__A2 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _09754_/B _09754_/C _10559_/A vssd1 vssd1 vccd1 vccd1 _09757_/C sky130_fd_sc_hd__a21o_1
X_06967_ _09772_/A _08821_/B _09478_/B2 fanout36/X vssd1 vssd1 vccd1 vccd1 _06968_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06898_ _06898_/A _06898_/B _06898_/C vssd1 vssd1 vccd1 vccd1 _06904_/B sky130_fd_sc_hd__or3_2
X_08706_ _07984_/B _07999_/B _07984_/A vssd1 vssd1 vccd1 vccd1 _08717_/A sky130_fd_sc_hd__o21ba_1
X_09686_ _09684_/Y _09686_/B vssd1 vssd1 vccd1 vccd1 _09686_/X sky130_fd_sc_hd__and2b_1
X_08637_ _08643_/A _08643_/B _09068_/A _08636_/X vssd1 vssd1 vccd1 vccd1 _09074_/A
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_96_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _08568_/A _08568_/B _08568_/C vssd1 vssd1 vccd1 vccd1 _08568_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout21 _07138_/X vssd1 vssd1 vccd1 vccd1 _12150_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08499_ _10458_/A _08499_/B vssd1 vssd1 vccd1 vccd1 _08507_/B sky130_fd_sc_hd__xnor2_1
X_07519_ _09622_/A _07519_/B vssd1 vssd1 vccd1 vccd1 _07525_/A sky130_fd_sc_hd__xor2_2
Xfanout43 _11147_/B vssd1 vssd1 vccd1 vccd1 _10551_/B sky130_fd_sc_hd__buf_12
Xfanout54 fanout55/X vssd1 vssd1 vccd1 vccd1 fanout54/X sky130_fd_sc_hd__buf_6
Xfanout65 _12774_/A vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__buf_6
Xfanout32 _07000_/X vssd1 vssd1 vccd1 vccd1 fanout32/X sky130_fd_sc_hd__buf_6
XANTENNA__10798__B1 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout76 _07062_/X vssd1 vssd1 vccd1 vccd1 _12768_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__07663__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout98 _08348_/B vssd1 vssd1 vccd1 vccd1 fanout98/X sky130_fd_sc_hd__buf_8
Xfanout87 _08842_/A vssd1 vssd1 vccd1 vccd1 _11499_/A sky130_fd_sc_hd__buf_12
X_10530_ _10705_/A _10531_/B vssd1 vssd1 vccd1 vccd1 _10530_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10461_ _10461_/A _10461_/B _10461_/C vssd1 vssd1 vccd1 vccd1 _10462_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11211__A1 _11181_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11747__C1 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ _12200_/A _12200_/B vssd1 vssd1 vccd1 vccd1 _12202_/B sky130_fd_sc_hd__xnor2_1
X_13180_ hold31/X _12721_/B hold177/A _06537_/A vssd1 vssd1 vccd1 vccd1 _13180_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_115_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10392_ _10392_/A _10392_/B vssd1 vssd1 vccd1 vccd1 _10392_/X sky130_fd_sc_hd__xor2_1
XANTENNA__11762__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12131_ _12131_/A _12131_/B vssd1 vssd1 vccd1 vccd1 _12133_/B sky130_fd_sc_hd__or2_1
X_12062_ _06596_/Y _09194_/Y _10638_/B vssd1 vssd1 vccd1 vccd1 _12062_/Y sky130_fd_sc_hd__a21oi_1
X_11013_ _11014_/A _11014_/B vssd1 vssd1 vccd1 vccd1 _11158_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08391__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08391__B2 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09078__C_N _09076_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11194__S _11194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12964_ _08443_/A _12744_/B hold158/X vssd1 vssd1 vccd1 vccd1 _13252_/D sky130_fd_sc_hd__a21boi_1
X_11915_ hold293/A _11989_/C _12119_/B1 vssd1 vssd1 vccd1 vccd1 _11915_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13019__A2 _06537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08694__A2 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12895_ hold211/X _12955_/A2 _13168_/B1 _13218_/Q vssd1 vssd1 vccd1 vccd1 hold212/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ curr_PC[22] _11929_/C _11845_/Y vssd1 vssd1 vccd1 vccd1 _11846_/Y sky130_fd_sc_hd__o21ai_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _11777_/A _11777_/B _11777_/C vssd1 vssd1 vccd1 vccd1 _11778_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_83_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10728_ _10728_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10959_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_51_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ _10660_/A _10660_/B vssd1 vssd1 vccd1 vccd1 _10659_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07406__B1 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08532__A _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12329_ _09396_/X _12328_/X _12361_/B vssd1 vssd1 vccd1 vccd1 _12329_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07148__A _08695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_45 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07709__A1 _07308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _07871_/B _07871_/C _08695_/A vssd1 vssd1 vccd1 vccd1 _07872_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__06987__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ reg1_val[18] _07075_/A vssd1 vssd1 vccd1 vccd1 _06821_/X sky130_fd_sc_hd__and2_1
X_06752_ _06752_/A _06923_/A _12588_/B vssd1 vssd1 vccd1 vccd1 _11746_/A sky130_fd_sc_hd__or3b_4
XFILLER_0_92_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09540_ _13218_/Q hold211/A vssd1 vssd1 vccd1 vccd1 _09540_/X sky130_fd_sc_hd__or2_1
X_09471_ _08311_/A _07149_/B _07435_/Y _09470_/Y vssd1 vssd1 vccd1 vccd1 _09472_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_78_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06683_ reg1_val[17] _06684_/B vssd1 vssd1 vccd1 vccd1 _06683_/X sky130_fd_sc_hd__or2_1
X_08422_ _08432_/A _08422_/B vssd1 vssd1 vccd1 vccd1 _08461_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07893__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08353_ _08544_/C _10551_/A vssd1 vssd1 vccd1 vccd1 _08355_/C sky130_fd_sc_hd__nand2_1
XANTENNA_fanout142_A _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08437__A2 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08284_ _08284_/A _08284_/B vssd1 vssd1 vccd1 vccd1 _08287_/B sky130_fd_sc_hd__xnor2_1
X_07304_ _08305_/B _08305_/C vssd1 vssd1 vccd1 vccd1 _10811_/A sky130_fd_sc_hd__and2_4
XFILLER_0_74_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11133__A _12255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07235_ fanout77/X _10156_/B2 _10156_/A1 fanout75/X vssd1 vssd1 vccd1 vccd1 _07236_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09398__B1 _12382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07166_ reg1_val[13] _07166_/B vssd1 vssd1 vccd1 vccd1 _09742_/A sky130_fd_sc_hd__xor2_4
X_07097_ _10169_/A _07097_/B vssd1 vssd1 vccd1 vccd1 _07098_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07058__A _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout222 _11194_/S vssd1 vssd1 vccd1 vccd1 _10750_/S sky130_fd_sc_hd__buf_4
Xfanout200 _09188_/X vssd1 vssd1 vccd1 vccd1 _12243_/B1 sky130_fd_sc_hd__buf_6
Xfanout211 _09359_/S vssd1 vssd1 vccd1 vccd1 _09365_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout233 _09384_/X vssd1 vssd1 vccd1 vccd1 _11398_/B sky130_fd_sc_hd__buf_2
XANTENNA__07176__A2 _07303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout244 _12373_/A1 vssd1 vssd1 vccd1 vccd1 _09173_/S sky130_fd_sc_hd__clkbuf_4
Xfanout255 _12487_/S vssd1 vssd1 vccd1 vccd1 _12382_/S sky130_fd_sc_hd__buf_4
Xfanout266 _06537_/Y vssd1 vssd1 vccd1 vccd1 _12723_/A sky130_fd_sc_hd__buf_4
Xfanout277 _12658_/A vssd1 vssd1 vccd1 vccd1 _12557_/A sky130_fd_sc_hd__buf_4
Xfanout288 _13116_/A vssd1 vssd1 vccd1 vccd1 _13169_/A sky130_fd_sc_hd__clkbuf_4
X_07999_ _07999_/A _07999_/B vssd1 vssd1 vccd1 vccd1 _08013_/A sky130_fd_sc_hd__xnor2_4
Xfanout299 _07134_/A vssd1 vssd1 vccd1 vccd1 _06864_/A sky130_fd_sc_hd__buf_6
X_09807_ _09808_/B _09808_/A vssd1 vssd1 vccd1 vccd1 _09807_/Y sky130_fd_sc_hd__nand2b_1
X_09738_ _09738_/A _09738_/B vssd1 vssd1 vccd1 vccd1 _09781_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_96_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _09342_/X _09344_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09669_/X sky130_fd_sc_hd__mux2_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12681_/A _12681_/B vssd1 vssd1 vccd1 vccd1 _12688_/A sky130_fd_sc_hd__nand2b_1
X_11700_ _11791_/B _11700_/B vssd1 vssd1 vccd1 vccd1 _11701_/B sky130_fd_sc_hd__or2_1
XFILLER_0_127_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07521__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09625__A1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11631_ _11633_/A vssd1 vssd1 vccd1 vccd1 _11631_/Y sky130_fd_sc_hd__inv_2
X_11562_ _06865_/A _11561_/X _12228_/B1 vssd1 vssd1 vccd1 vccd1 _11562_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09625__B2 _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13301_ _13303_/CLK _13301_/D vssd1 vssd1 vccd1 vccd1 hold277/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10513_ _06734_/B _12243_/B1 _09191_/X _06732_/Y _10512_/X vssd1 vssd1 vccd1 vccd1
+ _10513_/X sky130_fd_sc_hd__o221a_1
XANTENNA__07100__A2 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11493_ curr_PC[18] _11493_/B vssd1 vssd1 vccd1 vccd1 _11671_/C sky130_fd_sc_hd__and2_2
X_13232_ _13312_/CLK _13232_/D vssd1 vssd1 vccd1 vccd1 hold239/A sky130_fd_sc_hd__dfxtp_1
X_10444_ _11853_/A _10444_/B vssd1 vssd1 vccd1 vccd1 _10445_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09448__A _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13163_ _13163_/A fanout1/X vssd1 vssd1 vccd1 vccd1 _13163_/Y sky130_fd_sc_hd__nor2_1
X_10375_ _13224_/Q _10509_/C _12124_/B vssd1 vssd1 vccd1 vccd1 _10376_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12114_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12114_/X sky130_fd_sc_hd__or2_1
X_13094_ hold282/A _13093_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13094_/X sky130_fd_sc_hd__mux2_1
X_12045_ _12045_/A _12045_/B vssd1 vssd1 vccd1 vccd1 _12045_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06600__A _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09183__A _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12947_ hold183/X _12947_/A2 _12947_/B1 hold213/A vssd1 vssd1 vccd1 vccd1 hold184/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09864__A1 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09864__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12878_ _13135_/A _12877_/B _12800_/X vssd1 vssd1 vccd1 vccd1 _13140_/A sky130_fd_sc_hd__a21o_1
X_11829_ _11743_/B _11745_/B _11743_/A vssd1 vssd1 vccd1 vccd1 _11830_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_56_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07020_ _07175_/D _07021_/B vssd1 vssd1 vccd1 vccd1 _07050_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_101_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08971_ _08972_/B _08972_/A vssd1 vssd1 vccd1 vccd1 _08971_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07922_ _08836_/A _07922_/B vssd1 vssd1 vccd1 vccd1 _07924_/B sky130_fd_sc_hd__xnor2_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_07853_ _10565_/A _07853_/B vssd1 vssd1 vccd1 vccd1 _07855_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07158__A2 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10162__A1 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ _10498_/A _06802_/Y _06803_/X vssd1 vssd1 vccd1 vccd1 _06804_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10162__B2 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11128__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07784_ _07751_/A _07751_/B _07749_/X vssd1 vssd1 vccd1 vccd1 _07785_/C sky130_fd_sc_hd__o21bai_1
XANTENNA__09304__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13100__B2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06735_ reg2_val[8] _06778_/B vssd1 vssd1 vccd1 vccd1 _06735_/X sky130_fd_sc_hd__and2_1
X_09523_ _09136_/X _09140_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _10112_/B sky130_fd_sc_hd__mux2_1
XANTENNA__09821__A _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11111__B1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07866__B1 _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06666_ _06668_/A vssd1 vssd1 vccd1 vccd1 _06666_/Y sky130_fd_sc_hd__inv_2
X_09454_ _09453_/B _09454_/B vssd1 vssd1 vccd1 vccd1 _09455_/B sky130_fd_sc_hd__and2b_1
X_08405_ _08619_/A _08619_/B _08621_/A vssd1 vssd1 vccd1 vccd1 _08405_/Y sky130_fd_sc_hd__a21oi_1
X_09385_ hold279/A hold240/A _09385_/C vssd1 vssd1 vccd1 vccd1 _09385_/X sky130_fd_sc_hd__and3_1
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07341__A _10180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08336_ _08336_/A _08336_/B vssd1 vssd1 vccd1 vccd1 _08341_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_108_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06597_ reg1_val[25] _07157_/A vssd1 vssd1 vccd1 vccd1 _06597_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_47_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09607__A1 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09607__B2 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08267_ _07004_/X _08477_/B _08776_/B1 _12734_/A vssd1 vssd1 vccd1 vccd1 _08268_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10622__C1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08198_ _08198_/A _08198_/B vssd1 vssd1 vccd1 vccd1 _08201_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07218_ _12782_/A _08758_/A2 fanout20/X _06864_/A vssd1 vssd1 vccd1 vccd1 _07219_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07149_ _07149_/A _07149_/B vssd1 vssd1 vccd1 vccd1 _07149_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_42_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07397__A2 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ _10160_/A _10160_/B vssd1 vssd1 vccd1 vccd1 _10161_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_30_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10091_ _10091_/A _10091_/B vssd1 vssd1 vccd1 vccd1 _10094_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_100_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08346__A1 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08346__B2 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__B1 _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12801_ hold293/A hold15/X vssd1 vssd1 vccd1 vccd1 _13130_/A sky130_fd_sc_hd__nand2b_1
X_10993_ _10984_/Y _10985_/X _10992_/Y _09115_/X _10991_/X vssd1 vssd1 vccd1 vccd1
+ _10993_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07857__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12732_ hold105/X _12744_/B vssd1 vssd1 vccd1 vccd1 hold106/A sky130_fd_sc_hd__or2_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08347__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07321__A2 _07317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ reg1_val[21] _12714_/A vssd1 vssd1 vccd1 vccd1 _12664_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_32_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12594_ _12592_/Y _12594_/B vssd1 vssd1 vccd1 vccd1 _12595_/B sky130_fd_sc_hd__nand2b_2
X_11614_ _11614_/A _11614_/B vssd1 vssd1 vccd1 vccd1 _11626_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_108_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11545_ _11632_/B _11545_/B vssd1 vssd1 vccd1 vccd1 _11547_/C sky130_fd_sc_hd__and2_1
X_11476_ _11476_/A _11476_/B vssd1 vssd1 vccd1 vccd1 _11478_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13215_ _13306_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10427_ _12022_/A _10427_/B vssd1 vssd1 vccd1 vccd1 _10429_/B sky130_fd_sc_hd__xnor2_1
X_13146_ hold264/X _13165_/A2 _13145_/X _13146_/B2 vssd1 vssd1 vccd1 vccd1 hold265/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09906__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10358_ _10360_/A _10360_/B vssd1 vssd1 vccd1 vccd1 _10358_/X sky130_fd_sc_hd__or2_1
X_13077_ _13077_/A _13077_/B vssd1 vssd1 vccd1 vccd1 _13078_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11647__S _11647_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10289_ _07073_/B _12349_/A _10458_/A vssd1 vssd1 vccd1 vccd1 _10289_/Y sky130_fd_sc_hd__a21oi_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12028_ _12029_/A _12029_/B vssd1 vssd1 vccd1 vccd1 _12098_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10144__B2 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10144__A1 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07145__B _07148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10787__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09170_ reg1_val[21] reg1_val[10] _09172_/S vssd1 vssd1 vccd1 vccd1 _09170_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08121_ _08121_/A _08121_/B vssd1 vssd1 vccd1 vccd1 _08161_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08273__B1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08052_ _08060_/B _08060_/A vssd1 vssd1 vccd1 vccd1 _08062_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11411__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07003_ _07303_/B _07175_/A _07001_/X _06795_/B vssd1 vssd1 vccd1 vccd1 _07004_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_3_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08025__B1 _07869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout105_A _07034_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09816__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ _08954_/A _08954_/B vssd1 vssd1 vccd1 vccd1 _08955_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07905_ _07907_/A _07907_/B vssd1 vssd1 vccd1 vccd1 _07905_/Y sky130_fd_sc_hd__nor2_1
X_08885_ _08881_/A _08881_/B _08879_/X vssd1 vssd1 vccd1 vccd1 _08932_/A sky130_fd_sc_hd__a21o_2
X_07836_ _07790_/B _07790_/C _07790_/A vssd1 vssd1 vccd1 vccd1 _07840_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_98_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07767_ _07767_/A _07767_/B vssd1 vssd1 vccd1 vccd1 _07770_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_79_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06718_ _07018_/A vssd1 vssd1 vccd1 vccd1 _06807_/B sky130_fd_sc_hd__inv_2
X_09506_ _09506_/A _09506_/B vssd1 vssd1 vccd1 vccd1 _09816_/A sky130_fd_sc_hd__xnor2_4
X_07698_ _07695_/Y _07698_/B vssd1 vssd1 vccd1 vccd1 _08966_/B sky130_fd_sc_hd__and2b_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07071__A _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06649_ _06649_/A _12583_/B vssd1 vssd1 vccd1 vccd1 _06649_/Y sky130_fd_sc_hd__nor2_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09437_ _09437_/A _09437_/B vssd1 vssd1 vccd1 vccd1 _09487_/A sky130_fd_sc_hd__xnor2_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ _09364_/X _09367_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09368_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_35_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08319_ _08733_/A _08319_/B vssd1 vssd1 vccd1 vccd1 _08345_/A sky130_fd_sc_hd__xor2_2
XANTENNA_fanout18_A _12786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09299_ _10559_/A _09300_/B vssd1 vssd1 vccd1 vccd1 _09302_/C sky130_fd_sc_hd__and2_1
XANTENNA_60 reg2_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_82 reg1_val[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_71 reg1_val[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _11444_/B _11330_/B vssd1 vssd1 vccd1 vccd1 _11342_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11321__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12899__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11261_ _11262_/A _11262_/B _11262_/C _11262_/D vssd1 vssd1 vccd1 vccd1 _11261_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11040__B _11041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11192_ _11088_/A _11088_/B _11086_/A vssd1 vssd1 vccd1 vccd1 _11193_/B sky130_fd_sc_hd__o21a_1
X_13000_ _11604_/A _13020_/B2 hold108/X vssd1 vssd1 vccd1 vccd1 hold109/A sky130_fd_sc_hd__o21a_1
X_10212_ _10212_/A _10212_/B vssd1 vssd1 vccd1 vccd1 _10215_/A sky130_fd_sc_hd__nand2_1
X_10143_ _10086_/A _10086_/B _10087_/Y vssd1 vssd1 vccd1 vccd1 _10224_/A sky130_fd_sc_hd__a21bo_1
X_10074_ _10075_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10074_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_89_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10976_ _10976_/A _10976_/B vssd1 vssd1 vccd1 vccd1 _10978_/A sky130_fd_sc_hd__nand2_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12715_ hold171/X hold137/X vssd1 vssd1 vccd1 vccd1 _12715_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12646_ reg1_val[17] _12714_/A vssd1 vssd1 vccd1 vccd1 _12657_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_26_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12577_ reg1_val[4] _12578_/B vssd1 vssd1 vccd1 vccd1 _12577_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10062__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11528_ _11528_/A vssd1 vssd1 vccd1 vccd1 _11529_/B sky130_fd_sc_hd__inv_2
XFILLER_0_40_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11459_ _11275_/A _11368_/Y _11370_/B vssd1 vssd1 vccd1 vccd1 _11459_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09755__B1 _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09636__A _09637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13129_ _13147_/A _13129_/B vssd1 vssd1 vccd1 vccd1 _13303_/D sky130_fd_sc_hd__and2_1
XANTENNA__11562__B1 _12228_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07230__A1 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07230__B2 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10117__A1 _11194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08670_ _08420_/B fanout94/X _12752_/A _08854_/B2 vssd1 vssd1 vccd1 vccd1 _08671_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09371__A _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ _07621_/A _07621_/B vssd1 vssd1 vccd1 vccd1 _07703_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07552_ _07549_/B _07599_/B _07549_/A vssd1 vssd1 vccd1 vccd1 _07577_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_76_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08494__B1 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07483_ _09316_/A _07483_/B vssd1 vssd1 vccd1 vccd1 _07485_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_118_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09222_ curr_PC[0] curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09153_ _09149_/X _09152_/X _09676_/S vssd1 vssd1 vccd1 vccd1 _09153_/X sky130_fd_sc_hd__mux2_1
X_08104_ _08123_/A _08102_/Y _08092_/Y vssd1 vssd1 vccd1 vccd1 _08112_/A sky130_fd_sc_hd__a21o_1
XANTENNA_fanout222_A _11194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10053__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09084_ _09031_/A _09031_/B _09032_/A _09098_/A vssd1 vssd1 vccd1 vccd1 _09086_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08035_ _08032_/Y _08106_/B _08031_/Y vssd1 vssd1 vccd1 vccd1 _08050_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_440 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09986_ _06795_/B _11923_/A2 _12243_/B1 _06758_/B _09985_/X vssd1 vssd1 vccd1 vccd1
+ _09986_/Y sky130_fd_sc_hd__o221ai_1
X_08937_ _08937_/A vssd1 vssd1 vccd1 vccd1 _08937_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_99_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08868_ _08782_/A _08782_/B _08783_/X vssd1 vssd1 vccd1 vccd1 _08873_/A sky130_fd_sc_hd__a21o_1
X_07819_ _08572_/B _07168_/Y _11147_/A _07117_/Y vssd1 vssd1 vccd1 vccd1 _07820_/B
+ sky130_fd_sc_hd__a22o_1
X_08799_ _08800_/B _08800_/A vssd1 vssd1 vccd1 vccd1 _08883_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_79_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10830_ _10707_/A _10707_/B _10706_/A vssd1 vssd1 vccd1 vccd1 _10832_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__11608__A1 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11608__B2 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10761_ reg1_val[11] _07018_/A _10638_/B vssd1 vssd1 vccd1 vccd1 _10761_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12500_ _12500_/A _12500_/B vssd1 vssd1 vccd1 vccd1 _12515_/B sky130_fd_sc_hd__or2_1
XFILLER_0_82_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10692_ _12206_/A _10692_/B vssd1 vssd1 vccd1 vccd1 _10695_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_125_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12431_ reg1_val[8] curr_PC[8] _12524_/S vssd1 vssd1 vccd1 vccd1 _12433_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_35_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10044__B1 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12147__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12362_ _12362_/A _12362_/B vssd1 vssd1 vccd1 vccd1 _12362_/Y sky130_fd_sc_hd__nand2_1
X_12293_ _09183_/Y _12284_/B _12292_/Y _06585_/B _12291_/X vssd1 vssd1 vccd1 vccd1
+ _12293_/X sky130_fd_sc_hd__a221o_1
X_11313_ curr_PC[16] _11314_/C curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11313_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07460__B2 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07460__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11244_ _11244_/A _11244_/B vssd1 vssd1 vccd1 vccd1 _11252_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11197__S _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11175_ _10956_/X _11066_/Y _11068_/B vssd1 vssd1 vccd1 vccd1 _11175_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10126_ _06996_/A _06928_/X wire201/X _06748_/X _10125_/Y vssd1 vssd1 vccd1 vccd1
+ _10126_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11847__A1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ _10155_/A _07056_/B _12349_/A _10056_/Y vssd1 vssd1 vccd1 vccd1 _10147_/B
+ sky130_fd_sc_hd__a31o_2
XANTENNA__11226__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09268__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10959_ _10959_/A _10959_/B _10959_/C vssd1 vssd1 vccd1 vccd1 _11174_/A sky130_fd_sc_hd__and3_1
XFILLER_0_85_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12629_ _12629_/A _12629_/B _12629_/C vssd1 vssd1 vccd1 vccd1 _12630_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 hold116/A vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold138 hold138/A vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 hold149/A vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08270__A _10819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07203__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09840_ hold224/A _11820_/A _10119_/C _09839_/Y _12290_/C1 vssd1 vssd1 vccd1 vccd1
+ _09840_/X sky130_fd_sc_hd__a311o_1
XANTENNA__07203__B2 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06983_ _06795_/B _10752_/S _06951_/C _07135_/B vssd1 vssd1 vccd1 vccd1 _06996_/B
+ sky130_fd_sc_hd__a31o_2
X_09771_ _09771_/A _09771_/B vssd1 vssd1 vccd1 vccd1 _09780_/A sky130_fd_sc_hd__xnor2_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _08722_/A _08722_/B vssd1 vssd1 vccd1 vccd1 _08800_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06962__B1 _12370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08653_ _08654_/A _08654_/B vssd1 vssd1 vccd1 vccd1 _08766_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_96_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout172_A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08584_ _08585_/B _08585_/A vssd1 vssd1 vccd1 vccd1 _08584_/X sky130_fd_sc_hd__and2b_1
X_07604_ _07604_/A _07604_/B vssd1 vssd1 vccd1 vccd1 _07621_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09259__A2 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07535_ _07278_/B _09476_/A fanout7/X _08825_/A2 vssd1 vssd1 vccd1 vccd1 _07536_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10274__B1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07466_ _09772_/A _07389_/B fanout26/X _09478_/B2 vssd1 vssd1 vccd1 vccd1 _07467_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09205_ _12713_/A _09205_/B vssd1 vssd1 vccd1 vccd1 _09213_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10694__B _12255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07397_ _10557_/A _09273_/A1 _07157_/Y _08588_/B vssd1 vssd1 vccd1 vccd1 _07398_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12015__A1 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09136_ _09134_/X _09135_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09136_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10577__A1 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ _11559_/B _11559_/C vssd1 vssd1 vccd1 vccd1 _09069_/A sky130_fd_sc_hd__or2_1
XFILLER_0_71_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10577__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07442__B2 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07442__A1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08018_ _08638_/A _08638_/B vssd1 vssd1 vccd1 vccd1 _08018_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07745__A2 _08774_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ _09968_/A _06794_/Y _09968_/Y vssd1 vssd1 vccd1 vccd1 _09970_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout85_A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12980_ _10453_/A _12980_/A2 hold96/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__o21a_1
XFILLER_0_87_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11931_ _10400_/S _11928_/X _11930_/Y _11927_/X vssd1 vssd1 vccd1 vccd1 dest_val[23]
+ sky130_fd_sc_hd__a31o_4
XANTENNA__08170__A2 _08348_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07243__B _12250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11862_ _11955_/A _11862_/B vssd1 vssd1 vccd1 vccd1 _11864_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12254__A1 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10813_ _10813_/A _10813_/B vssd1 vssd1 vccd1 vccd1 _10815_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11793_ _11793_/A _12255_/B vssd1 vssd1 vccd1 vccd1 _11795_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08355__A _08695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10744_ _10743_/A _10743_/B _12277_/B1 vssd1 vssd1 vccd1 vccd1 _10744_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07681__B2 _07034_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07681__A1 _07023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12006__A1 _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10675_ _10824_/B _10675_/B vssd1 vssd1 vccd1 vccd1 _10699_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_125_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12414_ _12415_/A _12415_/B _12415_/C vssd1 vssd1 vccd1 vccd1 _12422_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_63_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12345_ _12345_/A _12345_/B vssd1 vssd1 vccd1 vccd1 dest_val[30] sky130_fd_sc_hd__nor2_8
XFILLER_0_2_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12276_ _12276_/A _12276_/B vssd1 vssd1 vccd1 vccd1 _12276_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11517__B1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11227_ fanout32/X _11935_/A _12772_/A fanout29/X vssd1 vssd1 vccd1 vccd1 _11228_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12190__B1 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158_ _11158_/A _11158_/B _11156_/Y vssd1 vssd1 vccd1 vccd1 _11159_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_4_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10109_ _10108_/A _10108_/B _12228_/B1 vssd1 vssd1 vccd1 vccd1 _10109_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_65_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11089_ _11089_/A _11089_/B vssd1 vssd1 vccd1 vccd1 _11089_/X sky130_fd_sc_hd__or2_1
XFILLER_0_78_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12245__A1 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07320_ _11499_/A _07317_/B _09926_/A vssd1 vssd1 vccd1 vccd1 _07322_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_116_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07251_ _11431_/A fanout98/X fanout56/X _11347_/A vssd1 vssd1 vccd1 vccd1 _07252_/B
+ sky130_fd_sc_hd__o22a_1
X_07182_ _08733_/A _07174_/B _07180_/X vssd1 vssd1 vccd1 vccd1 _07182_/X sky130_fd_sc_hd__a21o_4
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10035__A _10035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _09040_/B _09821_/X _09822_/Y vssd1 vssd1 vccd1 vccd1 _09823_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12250__A _12250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ _10559_/A _09754_/B _09754_/C vssd1 vssd1 vccd1 vccd1 _09757_/B sky130_fd_sc_hd__nand3_1
X_06966_ _12022_/A _12078_/A _06965_/X vssd1 vssd1 vccd1 vccd1 _06966_/Y sky130_fd_sc_hd__a21oi_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08705_ _08705_/A _08705_/B vssd1 vssd1 vccd1 vccd1 _08720_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_69_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09685_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09686_/B sky130_fd_sc_hd__nand2_1
X_06897_ instruction[13] _06897_/B vssd1 vssd1 vccd1 vccd1 dest_pred[2] sky130_fd_sc_hd__and2_4
X_08636_ _09072_/A _09070_/D vssd1 vssd1 vccd1 vccd1 _08636_/X sky130_fd_sc_hd__and2_2
XFILLER_0_96_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10495__B1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11039__A2 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12236__A1 _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12396__S _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08567_ _08568_/B _08567_/B _08567_/C vssd1 vssd1 vccd1 vccd1 _08577_/A sky130_fd_sc_hd__or3_1
XFILLER_0_49_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout22 _07138_/X vssd1 vssd1 vccd1 vccd1 fanout22/X sky130_fd_sc_hd__clkbuf_8
Xfanout11 _07322_/X vssd1 vssd1 vccd1 vccd1 _11603_/A sky130_fd_sc_hd__buf_8
X_08498_ _08528_/A _08528_/B vssd1 vssd1 vccd1 vccd1 _08529_/A sky130_fd_sc_hd__nor2_1
Xfanout33 _06989_/X vssd1 vssd1 vccd1 vccd1 fanout33/X sky130_fd_sc_hd__buf_8
Xfanout44 _11147_/B vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__clkbuf_8
X_07518_ _09273_/A1 fanout20/X fanout18/X _08588_/B vssd1 vssd1 vccd1 vccd1 _07519_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout55 _07195_/X vssd1 vssd1 vccd1 vccd1 fanout55/X sky130_fd_sc_hd__buf_8
XANTENNA__10798__A1 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07663__B2 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07663__A1 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout66 _10280_/A vssd1 vssd1 vccd1 vccd1 _12206_/A sky130_fd_sc_hd__clkbuf_16
Xfanout88 _08836_/A vssd1 vssd1 vccd1 vccd1 _11429_/A sky130_fd_sc_hd__clkbuf_16
Xfanout77 _11794_/A vssd1 vssd1 vccd1 vccd1 fanout77/X sky130_fd_sc_hd__buf_8
XFILLER_0_36_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10798__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07449_ _11347_/A fanout95/X fanout54/X _11134_/B2 vssd1 vssd1 vccd1 vccd1 _07450_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_107_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06602__A_N _07126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10460_ _10461_/A _10461_/B _10461_/C vssd1 vssd1 vccd1 vccd1 _10462_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_60_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09119_ reg1_val[2] reg1_val[29] _09158_/S vssd1 vssd1 vccd1 vccd1 _09119_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12425__A _12593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10391_ _10389_/Y _10391_/B vssd1 vssd1 vccd1 vccd1 _10392_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_103_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12130_ _09851_/B _12118_/X _12121_/Y _12129_/X vssd1 vssd1 vccd1 vccd1 _12130_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07519__A _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ hold209/A _12124_/B _12122_/B _12290_/C1 vssd1 vssd1 vccd1 vccd1 _12061_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11012_ _11012_/A _11147_/B vssd1 vssd1 vccd1 vccd1 _11014_/B sky130_fd_sc_hd__nand2_2
XANTENNA__08391__A2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12963_ hold83/X _12723_/A _13170_/B hold157/X _13179_/A vssd1 vssd1 vccd1 vccd1
+ hold158/A sky130_fd_sc_hd__o221a_1
XFILLER_0_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11914_ _11197_/S _11912_/Y _11913_/X _09851_/B vssd1 vssd1 vccd1 vccd1 _11926_/A
+ sky130_fd_sc_hd__o211a_1
X_12894_ _13169_/A _12894_/B vssd1 vssd1 vccd1 vccd1 _13217_/D sky130_fd_sc_hd__and2_1
XFILLER_0_87_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11845_ curr_PC[22] _11929_/C _12556_/S vssd1 vssd1 vccd1 vccd1 _11845_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08085__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11776_ _11777_/A _11777_/B _11777_/C vssd1 vssd1 vccd1 vccd1 _11778_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10727_ _10728_/A _10728_/B vssd1 vssd1 vccd1 vccd1 _10727_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_42_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07406__A1 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10658_ _10658_/A _10658_/B vssd1 vssd1 vccd1 vccd1 _10660_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07406__B2 _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08532__B _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10589_ _10589_/A _10589_/B vssd1 vssd1 vccd1 vccd1 _10602_/A sky130_fd_sc_hd__xnor2_4
X_12328_ reg1_val[30] _12361_/C vssd1 vssd1 vccd1 vccd1 _12328_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07148__B _07148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12259_ _12258_/B _12259_/B vssd1 vssd1 vccd1 vccd1 _12260_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_76_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07709__A2 _07308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06987__B _06987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ _06865_/C _06818_/X _06819_/Y vssd1 vssd1 vccd1 vccd1 _06820_/Y sky130_fd_sc_hd__o21ai_1
X_06751_ _06541_/Y _06572_/X _06575_/Y _12588_/B _06898_/A vssd1 vssd1 vccd1 vccd1
+ _12284_/A sky130_fd_sc_hd__o2111a_4
X_06682_ reg1_val[17] _06684_/B vssd1 vssd1 vccd1 vccd1 _06685_/A sky130_fd_sc_hd__nor2_1
X_09470_ _07155_/X _07435_/Y _08443_/A vssd1 vssd1 vccd1 vccd1 _09470_/Y sky130_fd_sc_hd__a21oi_1
X_08421_ _08421_/A _08421_/B vssd1 vssd1 vccd1 vccd1 _08422_/B sky130_fd_sc_hd__and2_1
XFILLER_0_59_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07342__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07893__A1 _07004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__B2 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08352_ _07313_/A _07313_/B _07134_/A vssd1 vssd1 vccd1 vccd1 _08355_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_73_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08283_ _08283_/A _08283_/B vssd1 vssd1 vccd1 vccd1 _08287_/A sky130_fd_sc_hd__xnor2_1
X_07303_ _07303_/A _07303_/B _07303_/C vssd1 vssd1 vccd1 vccd1 _08305_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout135_A _07073_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07234_ _07234_/A _07234_/B vssd1 vssd1 vccd1 vccd1 _07237_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07165_ _07165_/A _07165_/B vssd1 vssd1 vccd1 vccd1 _07166_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12941__A2 _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07096_ _10169_/A _07097_/B vssd1 vssd1 vccd1 vccd1 _07098_/A sky130_fd_sc_hd__or2_1
XFILLER_0_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout223 _06767_/X vssd1 vssd1 vccd1 vccd1 _11194_/S sky130_fd_sc_hd__buf_4
Xfanout212 _09362_/S vssd1 vssd1 vccd1 vccd1 _09359_/S sky130_fd_sc_hd__buf_4
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout234 _09384_/X vssd1 vssd1 vccd1 vccd1 _09842_/B sky130_fd_sc_hd__buf_4
Xfanout256 _12487_/S vssd1 vssd1 vccd1 vccd1 _12524_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__11901__B1 _09076_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout245 _12373_/A1 vssd1 vssd1 vccd1 vccd1 _09158_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06897__B _06897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout289 _13116_/A vssd1 vssd1 vccd1 vccd1 _13147_/A sky130_fd_sc_hd__buf_4
Xfanout267 _12955_/A2 vssd1 vssd1 vccd1 vccd1 _12947_/A2 sky130_fd_sc_hd__buf_4
X_07998_ _07998_/A _07998_/B vssd1 vssd1 vccd1 vccd1 _07999_/B sky130_fd_sc_hd__xnor2_4
Xfanout278 _12658_/A vssd1 vssd1 vccd1 vccd1 _12714_/A sky130_fd_sc_hd__buf_12
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09806_ _09806_/A _09806_/B vssd1 vssd1 vccd1 vccd1 _09808_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07074__A _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06949_ _11194_/S _07279_/A _09392_/S _09362_/S vssd1 vssd1 vccd1 vccd1 _07175_/A
+ sky130_fd_sc_hd__or4_4
X_09737_ _09735_/X _09737_/B vssd1 vssd1 vccd1 vccd1 _09738_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09668_ _10617_/A _09668_/B _09668_/C vssd1 vssd1 vccd1 vccd1 _09668_/X sky130_fd_sc_hd__or3_1
XANTENNA__07333__B1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout48_A _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08619_ _08619_/A _08619_/B vssd1 vssd1 vccd1 vccd1 _09060_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_84_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09599_ _09599_/A _09599_/B vssd1 vssd1 vccd1 vccd1 _09638_/A sky130_fd_sc_hd__or2_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11630_ _11632_/A _11632_/B _11632_/C vssd1 vssd1 vccd1 vccd1 _11633_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_126_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11561_ _06822_/Y _11560_/X _11738_/S vssd1 vssd1 vccd1 vccd1 _11561_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09625__A2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13300_ _13303_/CLK _13300_/D vssd1 vssd1 vccd1 vccd1 hold280/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10640__B1 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10512_ _07325_/A _11923_/A2 _10377_/B reg1_val[9] _12487_/S vssd1 vssd1 vccd1 vccd1
+ _10512_/X sky130_fd_sc_hd__o221a_1
X_11492_ _11184_/A _11468_/Y _11491_/X _11466_/X vssd1 vssd1 vccd1 vccd1 _11492_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_80_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09389__A1 _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13231_ _13312_/CLK hold182/X vssd1 vssd1 vccd1 vccd1 hold180/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11196__A1 _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10443_ fanout33/X _11431_/A fanout70/X _10553_/A vssd1 vssd1 vccd1 vccd1 _10444_/B
+ sky130_fd_sc_hd__o22a_1
X_13162_ _13162_/A _13162_/B vssd1 vssd1 vccd1 vccd1 _13162_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11735__A3 _09073_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10374_ _10373_/A _10373_/B _10373_/Y _12228_/B1 vssd1 vssd1 vccd1 vccd1 _10395_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12113_ reg1_val[26] curr_PC[26] vssd1 vssd1 vccd1 vccd1 _12113_/Y sky130_fd_sc_hd__nor2_1
X_13093_ _13093_/A _13093_/B vssd1 vssd1 vccd1 vccd1 _13093_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09464__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12044_ _06850_/X _12043_/X _12322_/S vssd1 vssd1 vccd1 vccd1 _12045_/B sky130_fd_sc_hd__mux2_1
XANTENNA__12602__B _12603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06600__B _12603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07080__A_N _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11656__C1 _06918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12946_ _12946_/A hold210/X vssd1 vssd1 vccd1 vccd1 _13243_/D sky130_fd_sc_hd__and2_1
XFILLER_0_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09864__A2 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12877_ _12800_/X _12877_/B vssd1 vssd1 vccd1 vccd1 _13135_/B sky130_fd_sc_hd__nand2b_1
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11828_ _11828_/A _11828_/B vssd1 vssd1 vccd1 vccd1 _11830_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11759_ _11749_/Y _11750_/X _11754_/X _11758_/X vssd1 vssd1 vccd1 vccd1 _11759_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_71_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12923__A2 _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07159__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08970_ _08970_/A _08970_/B vssd1 vssd1 vccd1 vccd1 _08972_/B sky130_fd_sc_hd__xnor2_1
X_07921_ _08819_/B2 _08134_/B fanout51/X _12730_/A vssd1 vssd1 vccd1 vccd1 _07922_/B
+ sky130_fd_sc_hd__o22a_1
X_07852_ _08821_/A _07852_/B vssd1 vssd1 vccd1 vccd1 _07853_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09552__A1 _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11409__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06803_ reg1_val[9] _07325_/A vssd1 vssd1 vccd1 vccd1 _06803_/X sky130_fd_sc_hd__and2_1
XANTENNA__10162__A2 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13100__A2 _13151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07783_ _07783_/A _07783_/B vssd1 vssd1 vccd1 vccd1 _07785_/B sky130_fd_sc_hd__xor2_1
X_09522_ _09520_/X _09521_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09522_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_36_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09304__B2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09304__A1 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06734_ _06732_/Y _06734_/B vssd1 vssd1 vccd1 vccd1 _10498_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11111__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11111__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07866__A1 _08572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06665_ _07077_/A reg1_val[19] vssd1 vssd1 vccd1 vccd1 _06668_/A sky130_fd_sc_hd__and2b_1
XANTENNA__11662__A2 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09453_ _09454_/B _09453_/B vssd1 vssd1 vccd1 vccd1 _09596_/D sky130_fd_sc_hd__and2b_1
X_08404_ _08620_/A _08620_/B _08620_/C vssd1 vssd1 vccd1 vccd1 _08621_/A sky130_fd_sc_hd__o21a_1
X_09384_ hold33/A _11823_/S vssd1 vssd1 vccd1 vccd1 _09384_/X sky130_fd_sc_hd__and2_2
XFILLER_0_59_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08335_ _08344_/B _08344_/A vssd1 vssd1 vccd1 vccd1 _08336_/B sky130_fd_sc_hd__nand2b_1
X_06596_ _07157_/A reg1_val[25] vssd1 vssd1 vccd1 vccd1 _06596_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_47_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09607__A2 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08266_ _08773_/A _08266_/B vssd1 vssd1 vccd1 vccd1 _08328_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07094__A2 _07087_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ _08205_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08197_/X sky130_fd_sc_hd__or2_1
X_07217_ _07243_/A _07217_/B vssd1 vssd1 vccd1 vccd1 _12784_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07148_ _08695_/A _07148_/B vssd1 vssd1 vccd1 vccd1 _07150_/B sky130_fd_sc_hd__or2_1
XFILLER_0_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07079_ _07079_/A _07079_/B vssd1 vssd1 vccd1 vccd1 _11511_/A sky130_fd_sc_hd__nand2_4
X_10090_ _10090_/A _10090_/B vssd1 vssd1 vccd1 vccd1 _10091_/B sky130_fd_sc_hd__xor2_4
XANTENNA__08346__A2 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__A1 _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__B2 _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11319__A _11695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10689__B1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__B1 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12800_ hold19/X hold256/X vssd1 vssd1 vccd1 vccd1 _12800_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11102__A1 _09198_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10992_ _11195_/A _09532_/X _09214_/A vssd1 vssd1 vccd1 vccd1 _10992_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__07857__B2 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07857__A1 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12731_ hold29/X _12744_/B _12730_/Y _13066_/A vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__o211a_1
XFILLER_0_97_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12662_ reg1_val[21] _12714_/A vssd1 vssd1 vccd1 vccd1 _12662_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11613_ _11613_/A _11613_/B vssd1 vssd1 vccd1 vccd1 _11614_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11405__A2 _11381_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12593_ reg1_val[7] _12593_/B vssd1 vssd1 vccd1 vccd1 _12594_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10893__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09459__A _10578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11544_ _11544_/A _11544_/B _11544_/C vssd1 vssd1 vccd1 vccd1 _11545_/B sky130_fd_sc_hd__or3_1
XFILLER_0_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11475_ reg1_val[18] curr_PC[18] vssd1 vssd1 vccd1 vccd1 _11476_/B sky130_fd_sc_hd__or2_1
XFILLER_0_122_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13214_ _13306_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
X_10426_ _08821_/B fanout57/X _07553_/A fanout36/X vssd1 vssd1 vccd1 vccd1 _10427_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13145_ hold286/A _13144_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13145_/X sky130_fd_sc_hd__mux2_1
XANTENNA_max_cap97_A _11147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10357_ _10357_/A _10357_/B vssd1 vssd1 vccd1 vccd1 _10360_/B sky130_fd_sc_hd__xnor2_2
X_13076_ _13086_/A _13076_/B vssd1 vssd1 vccd1 vccd1 _13292_/D sky130_fd_sc_hd__and2_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ _10453_/A _10288_/B vssd1 vssd1 vccd1 vccd1 _10292_/A sky130_fd_sc_hd__xnor2_1
X_12027_ _12027_/A _12027_/B vssd1 vssd1 vccd1 vccd1 _12029_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10144__A2 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09298__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13163__B fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12929_ hold178/X _13146_/B2 _12947_/B1 hold168/X vssd1 vssd1 vccd1 vccd1 hold179/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08120_ _08120_/A _08120_/B vssd1 vssd1 vccd1 vccd1 _08161_/A sky130_fd_sc_hd__and2_2
XFILLER_0_113_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08273__A1 _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08273__B2 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09470__B1 _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08051_ _08105_/A _08105_/B _08045_/Y vssd1 vssd1 vccd1 vccd1 _08060_/B sky130_fd_sc_hd__a21boi_2
XANTENNA__08025__A1 _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07002_ _06761_/Y _06951_/C _07135_/B _06972_/C vssd1 vssd1 vccd1 vccd1 _07004_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08025__B2 _09925_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06813__A_N _07192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10742__S _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09773__A1 _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08953_ _08953_/A _08953_/B vssd1 vssd1 vccd1 vccd1 _08954_/B sky130_fd_sc_hd__xnor2_2
X_07904_ _07904_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _07907_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08884_ _08884_/A _08884_/B vssd1 vssd1 vccd1 vccd1 _09098_/A sky130_fd_sc_hd__or2_4
XFILLER_0_47_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10043__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07835_ _07842_/A _07842_/B _07831_/B _07832_/Y vssd1 vssd1 vccd1 vccd1 _07841_/A
+ sky130_fd_sc_hd__o31ai_4
XANTENNA__13085__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07766_ _07767_/A _07767_/B vssd1 vssd1 vccd1 vccd1 _07766_/Y sky130_fd_sc_hd__nor2_1
X_06717_ _06783_/A _06641_/A _12620_/B _06716_/X vssd1 vssd1 vccd1 vccd1 _07018_/A
+ sky130_fd_sc_hd__a31o_2
X_09505_ _09506_/A _09506_/B vssd1 vssd1 vccd1 vccd1 _09505_/X sky130_fd_sc_hd__and2_1
XFILLER_0_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07697_ _07697_/A _07697_/B vssd1 vssd1 vccd1 vccd1 _07698_/B sky130_fd_sc_hd__nand2_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07071__B _07080_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09436_ _09436_/A _09436_/B vssd1 vssd1 vccd1 vccd1 _09437_/B sky130_fd_sc_hd__xor2_1
X_06648_ instruction[30] _06678_/B vssd1 vssd1 vccd1 vccd1 _12583_/B sky130_fd_sc_hd__and2_4
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06579_ _06898_/A _06579_/B vssd1 vssd1 vccd1 vccd1 _06579_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09367_ _09365_/X _09366_/X _09676_/S vssd1 vssd1 vccd1 vccd1 _09367_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_117_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_50 reg2_val[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08318_ _09283_/A _07173_/Y _07182_/X _09362_/S vssd1 vssd1 vccd1 vccd1 _08319_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09279__A _09620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09298_ fanout57/X _09752_/B fanout13/X _07553_/A vssd1 vssd1 vccd1 vccd1 _09300_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11602__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08249_ _08244_/A _08244_/B _08246_/B _08297_/A _08297_/B vssd1 vssd1 vccd1 vccd1
+ _08261_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_105_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_61 reg2_val[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_83 reg1_val[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_72 reg1_val[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11260_ _11148_/A _11148_/B _11151_/A vssd1 vssd1 vccd1 vccd1 _11264_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_120_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11191_ _11191_/A _11191_/B vssd1 vssd1 vccd1 vccd1 _11193_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12433__A _12598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10211_ _10020_/A _10020_/B _10019_/A vssd1 vssd1 vccd1 vccd1 _10216_/A sky130_fd_sc_hd__o21ai_2
X_10142_ _10091_/A _10091_/B _10089_/X vssd1 vssd1 vccd1 vccd1 _10227_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_100_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10073_ _10073_/A _10073_/B vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10126__A2 _06928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09742__A _09742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10975_ reg1_val[13] curr_PC[13] vssd1 vssd1 vccd1 vccd1 _10976_/B sky130_fd_sc_hd__or2_1
XFILLER_0_85_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ _12714_/A _12714_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[31] sky130_fd_sc_hd__xnor2_4
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12645_ reg1_val[16] _12714_/A _12657_/A vssd1 vssd1 vccd1 vccd1 _12647_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_38_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12576_ _12575_/A _12572_/Y _12574_/B vssd1 vssd1 vccd1 vccd1 _12580_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_108_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10062__A1 _07098_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10062__B2 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11527_ _11616_/B _11527_/B vssd1 vssd1 vccd1 vccd1 _11528_/A sky130_fd_sc_hd__or2_1
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13000__A1 _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09204__B1 _09200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08821__A _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11458_ _11456_/Y _11458_/B vssd1 vssd1 vccd1 vccd1 _11635_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_111_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11389_ _11387_/Y _11389_/B vssd1 vssd1 vccd1 vccd1 _11390_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10409_ fanout22/X fanout95/X fanout54/X _12150_/B vssd1 vssd1 vccd1 vccd1 _10410_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13128_ hold293/X _13165_/A2 _13127_/X _13146_/B2 vssd1 vssd1 vccd1 vccd1 _13129_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07230__A2 _10553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_13 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ hold292/A _13058_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13059_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07518__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11865__A2 _11786_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08191__B1 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07620_ _07620_/A _07620_/B vssd1 vssd1 vccd1 vccd1 _07707_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08268__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11078__B1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07172__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07551_ _10306_/A _07551_/B vssd1 vssd1 vccd1 vccd1 _07599_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08494__A1 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08494__B2 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07482_ _07482_/A _07482_/B _07583_/A vssd1 vssd1 vccd1 vccd1 _07483_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07900__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09221_ _10400_/S _09219_/X _09220_/X vssd1 vssd1 vccd1 vccd1 dest_val[0] sky130_fd_sc_hd__o21ai_4
XFILLER_0_33_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09152_ _09150_/X _09151_/X _09359_/S vssd1 vssd1 vccd1 vccd1 _09152_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08103_ _08103_/A _08103_/B vssd1 vssd1 vccd1 vccd1 _08123_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_71_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10053__B2 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10053__A1 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09083_ _08803_/Y _08884_/A _08884_/B vssd1 vssd1 vccd1 vccd1 _09086_/B sky130_fd_sc_hd__o21bai_1
XANTENNA_fanout215_A _12726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08034_ _08034_/A _08034_/B vssd1 vssd1 vccd1 vccd1 _08106_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_4_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12253__A _12255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07757__B1 _07325_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ reg1_val[5] _11099_/B _09983_/Y _09984_/X vssd1 vssd1 vccd1 vccd1 _09985_/X
+ sky130_fd_sc_hd__o22a_1
X_08936_ _08804_/B _09029_/B _08801_/X vssd1 vssd1 vccd1 vccd1 _08937_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07509__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08867_ _08770_/B _08785_/B _08768_/Y vssd1 vssd1 vccd1 vccd1 _08878_/A sky130_fd_sc_hd__a21oi_2
X_07818_ _07842_/A _07842_/B vssd1 vssd1 vccd1 vccd1 _07831_/A sky130_fd_sc_hd__nor2_2
XANTENNA__09281__B _09281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08178__A _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08798_ _08798_/A _08798_/B vssd1 vssd1 vccd1 vccd1 _08800_/B sky130_fd_sc_hd__xnor2_2
X_07749_ _08443_/A _07749_/B vssd1 vssd1 vccd1 vccd1 _07749_/X sky130_fd_sc_hd__xor2_1
XANTENNA__11608__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10760_ hold291/A _09385_/C _10877_/B _12339_/B1 vssd1 vssd1 vccd1 vccd1 _10760_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout30_A _07006_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09419_ _09645_/A _09419_/B vssd1 vssd1 vccd1 vccd1 _09421_/B sky130_fd_sc_hd__nand2_2
X_10691_ fanout27/X fanout57/X _07553_/A fanout26/X vssd1 vssd1 vccd1 vccd1 _10692_/B
+ sky130_fd_sc_hd__o22a_1
X_12430_ _12436_/B _12430_/B vssd1 vssd1 vccd1 vccd1 new_PC[7] sky130_fd_sc_hd__and2_4
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11332__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10044__A1 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12361_ reg1_val[30] _12361_/B _12361_/C vssd1 vssd1 vccd1 vccd1 _12362_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10044__B2 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12292_ _06583_/X _09383_/B _09191_/X vssd1 vssd1 vccd1 vccd1 _12292_/Y sky130_fd_sc_hd__o21ai_1
X_11312_ _10400_/S _11310_/Y _11311_/X _11309_/X vssd1 vssd1 vccd1 vccd1 dest_val[16]
+ sky130_fd_sc_hd__a31o_4
XANTENNA__07460__A2 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11243_ _11244_/B _11244_/A vssd1 vssd1 vccd1 vccd1 _11356_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_120_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07748__B1 _08692_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ _11174_/A _11374_/A vssd1 vssd1 vccd1 vccd1 _11174_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10125_ reg1_val[6] _11099_/B _10123_/Y _10124_/X vssd1 vssd1 vccd1 vccd1 _10125_/Y
+ sky130_fd_sc_hd__o22ai_2
X_10056_ _07047_/A _12349_/A _10155_/A vssd1 vssd1 vccd1 vccd1 _10056_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11507__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08088__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10958_ _10958_/A _10958_/B vssd1 vssd1 vccd1 vccd1 _11173_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07720__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10889_ _11107_/C _10888_/Y _10886_/X vssd1 vssd1 vccd1 vccd1 dest_val[12] sky130_fd_sc_hd__o21ai_4
X_12628_ _12629_/A _12629_/B _12629_/C vssd1 vssd1 vccd1 vccd1 _12635_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09425__B1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11232__B1 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12559_ reg1_val[0] _12560_/B vssd1 vssd1 vccd1 vccd1 _12565_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold106 hold106/A vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 hold117/A vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold139 hold139/A vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10338__A2 _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07203__A2 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06982_ _11604_/A _06987_/B vssd1 vssd1 vccd1 vccd1 _06982_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__06962__A1 _07279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09770_ _09770_/A _09770_/B vssd1 vssd1 vccd1 vccd1 _09771_/B sky130_fd_sc_hd__xnor2_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _08805_/B _08805_/A vssd1 vssd1 vccd1 vccd1 _08801_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__11838__A2 _11838_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09382__A _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08652_ _08773_/A _08652_/B vssd1 vssd1 vccd1 vccd1 _08654_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07911__B1 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07603_ _07603_/A _07603_/B vssd1 vssd1 vccd1 vccd1 _07621_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_95_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout165_A _07116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08583_ _08583_/A _08583_/B vssd1 vssd1 vccd1 vccd1 _08585_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07534_ _07090_/A _07090_/B _07277_/B _10551_/B _12301_/C vssd1 vssd1 vccd1 vccd1
+ fanout7/A sky130_fd_sc_hd__o41a_1
XANTENNA__08726__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07465_ _07584_/A _07584_/B _07452_/X vssd1 vssd1 vccd1 vccd1 _07485_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_107_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09204_ _06864_/Y _09197_/X _09200_/X hold240/A _09203_/X vssd1 vssd1 vccd1 vccd1
+ _09204_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_57_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07396_ _07396_/A _07396_/B _07396_/C vssd1 vssd1 vccd1 vccd1 _07401_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12015__A2 _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09135_ reg1_val[11] reg1_val[20] _09172_/S vssd1 vssd1 vccd1 vccd1 _09135_/X sky130_fd_sc_hd__mux2_1
X_09066_ _09070_/C _09066_/B vssd1 vssd1 vccd1 vccd1 _11559_/C sky130_fd_sc_hd__xor2_4
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10577__A2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07442__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08017_ _08638_/B _08638_/A vssd1 vssd1 vccd1 vccd1 _08017_/X sky130_fd_sc_hd__and2b_1
XANTENNA__06650__B1 _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09968_ _09968_/A _09968_/B vssd1 vssd1 vccd1 vccd1 _09968_/Y sky130_fd_sc_hd__nor2_1
X_08919_ _08919_/A _08919_/B vssd1 vssd1 vccd1 vccd1 _08922_/A sky130_fd_sc_hd__or2_2
XANTENNA_fanout78_A _07055_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ _12070_/C vssd1 vssd1 vccd1 vccd1 _11930_/Y sky130_fd_sc_hd__inv_2
X_09899_ _09900_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09899_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11861_ _11861_/A _11861_/B vssd1 vssd1 vccd1 vccd1 _11862_/B sky130_fd_sc_hd__and2_1
XFILLER_0_79_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11792_ _11878_/A _11792_/B vssd1 vssd1 vccd1 vccd1 _11795_/A sky130_fd_sc_hd__and2_1
XANTENNA__12254__A2 _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10812_ _10812_/A _10812_/B vssd1 vssd1 vccd1 vccd1 _10813_/B sky130_fd_sc_hd__xnor2_1
X_10743_ _10743_/A _10743_/B vssd1 vssd1 vccd1 vccd1 _10743_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07681__A2 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09407__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10674_ _10674_/A _10674_/B vssd1 vssd1 vccd1 vccd1 _10675_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_106_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12413_ _12422_/A _12413_/B vssd1 vssd1 vccd1 vccd1 _12415_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_62_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11214__B1 _11211_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12344_ _06834_/B _12250_/B _06930_/Y _12343_/X vssd1 vssd1 vccd1 vccd1 _12345_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__10973__C1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06603__B _07126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09186__B _09199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12275_ _06854_/Y _12274_/X _12322_/S vssd1 vssd1 vccd1 vccd1 _12276_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11517__B2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11517__A1 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11226_ _12206_/A _11226_/B vssd1 vssd1 vccd1 vccd1 _11230_/B sky130_fd_sc_hd__xnor2_1
X_11157_ _11158_/A _11158_/B _11156_/Y vssd1 vssd1 vccd1 vccd1 _11159_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10108_ _10108_/A _10108_/B vssd1 vssd1 vccd1 vccd1 _10108_/Y sky130_fd_sc_hd__nand2_1
X_11088_ _11088_/A _11088_/B vssd1 vssd1 vccd1 vccd1 _11088_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10039_ _10040_/A _10040_/B vssd1 vssd1 vccd1 vccd1 _10206_/B sky130_fd_sc_hd__and2_1
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08546__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07450__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07250_ _07250_/A _07250_/B vssd1 vssd1 vccd1 vccd1 _07272_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11205__B1 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07181_ _08733_/A _07174_/B _07180_/X vssd1 vssd1 vccd1 vccd1 _07181_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_60_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12953__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10035__B _11147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09822_ _09040_/B _09821_/X _11184_/A vssd1 vssd1 vccd1 vccd1 _09822_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09753_ _07308_/A _07308_/B _12760_/A vssd1 vssd1 vccd1 vccd1 _09754_/C sky130_fd_sc_hd__a21o_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08137__B1 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout282_A _06569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _08703_/B _08703_/C _08703_/A vssd1 vssd1 vccd1 vccd1 _08705_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__11147__A _11147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12250__B _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06965_ _12143_/A _11780_/A _06965_/C vssd1 vssd1 vccd1 vccd1 _06965_/X sky130_fd_sc_hd__and3_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09684_ reg1_val[3] curr_PC[3] vssd1 vssd1 vccd1 vccd1 _09684_/Y sky130_fd_sc_hd__nor2_1
X_06896_ instruction[12] _06897_/B vssd1 vssd1 vccd1 vccd1 dest_pred[1] sky130_fd_sc_hd__and2_4
X_08635_ _08635_/A _08635_/B vssd1 vssd1 vccd1 vccd1 _09070_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11692__B1 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _08568_/B _08567_/B _08567_/C vssd1 vssd1 vccd1 vccd1 _08568_/C sky130_fd_sc_hd__nor3_1
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07360__A _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout12 _07322_/X vssd1 vssd1 vccd1 vccd1 fanout12/X sky130_fd_sc_hd__buf_4
X_07517_ _09243_/B _07517_/B vssd1 vssd1 vccd1 vccd1 _07526_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout34 _06989_/X vssd1 vssd1 vccd1 vccd1 _09295_/A sky130_fd_sc_hd__buf_4
X_08497_ _08589_/A _08497_/B vssd1 vssd1 vccd1 vccd1 _08528_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout45 _07529_/Y vssd1 vssd1 vccd1 vccd1 _11147_/B sky130_fd_sc_hd__buf_6
Xfanout23 _12782_/A vssd1 vssd1 vccd1 vccd1 _12203_/A sky130_fd_sc_hd__clkbuf_8
Xfanout56 _07181_/Y vssd1 vssd1 vccd1 vccd1 fanout56/X sky130_fd_sc_hd__buf_8
XANTENNA__10798__A2 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07663__A2 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout67 _10280_/A vssd1 vssd1 vccd1 vccd1 _12255_/A sky130_fd_sc_hd__clkbuf_8
Xfanout89 _08836_/A vssd1 vssd1 vccd1 vccd1 _10180_/A sky130_fd_sc_hd__buf_6
Xfanout78 _07055_/Y vssd1 vssd1 vccd1 vccd1 _11794_/A sky130_fd_sc_hd__buf_8
X_07448_ _07448_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _07451_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_91_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07379_ _07379_/A _07379_/B vssd1 vssd1 vccd1 vccd1 _07385_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11747__A1 _11746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09118_ _09116_/X _09117_/X _12726_/A vssd1 vssd1 vccd1 vccd1 _09118_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10390_ reg1_val[8] curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10391_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09049_ _09049_/A _09049_/B _09049_/C vssd1 vssd1 vccd1 vccd1 _09050_/B sky130_fd_sc_hd__and3_1
XFILLER_0_102_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12060_ _12124_/B _12122_/B hold209/A vssd1 vssd1 vccd1 vccd1 _12060_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08376__B1 _08774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11011_ _12206_/A _11011_/B vssd1 vssd1 vccd1 vccd1 _11014_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06926__A1 _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06926__B2 _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10183__B1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12962_ _07148_/B _12742_/B hold84/X vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_99_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12893_ hold211/X _13168_/B1 fanout2/X _12955_/A2 vssd1 vssd1 vccd1 vccd1 _12894_/B
+ sky130_fd_sc_hd__a22o_1
X_11913_ _12361_/B _11913_/B vssd1 vssd1 vccd1 vccd1 _11913_/X sky130_fd_sc_hd__or2_1
XANTENNA__09340__A2 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10896__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11844_ _11184_/A _11819_/Y _11820_/X _11843_/X _11818_/X vssd1 vssd1 vccd1 vccd1
+ _11844_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_68_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__A1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11775_ _11864_/A _11775_/B vssd1 vssd1 vccd1 vccd1 _11777_/C sky130_fd_sc_hd__nand2_1
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10726_ _10728_/B _10728_/A vssd1 vssd1 vccd1 vccd1 _10726_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_125_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10657_ _11125_/A _10657_/B vssd1 vssd1 vccd1 vccd1 _10658_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12935__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11520__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_311 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06614__A _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07406__A2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10588_ _10588_/A _10588_/B vssd1 vssd1 vccd1 vccd1 _10589_/B sky130_fd_sc_hd__xor2_4
X_12327_ _12326_/A _12326_/B _12326_/Y _11184_/A vssd1 vssd1 vccd1 vccd1 _12327_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12258_ _12259_/B _12258_/B vssd1 vssd1 vccd1 vccd1 _12308_/A sky130_fd_sc_hd__and2b_1
X_11209_ _12373_/A1 _11208_/X _11196_/Y _09184_/X vssd1 vssd1 vccd1 vccd1 _11209_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_12189_ _12189_/A _12189_/B vssd1 vssd1 vccd1 vccd1 _12194_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07445__A _10180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06750_ _06750_/A _06750_/B vssd1 vssd1 vccd1 vccd1 _10108_/A sky130_fd_sc_hd__and2_1
XFILLER_0_116_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06681_ _06679_/Y _06680_/B1 _06569_/X reg2_val[17] vssd1 vssd1 vccd1 vccd1 _06684_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_78_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08420_ _08588_/A _08420_/B vssd1 vssd1 vccd1 vccd1 _08461_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07342__A1 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07342__B2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07893__A2 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08351_ _08365_/A _08351_/B vssd1 vssd1 vccd1 vccd1 _08351_/X sky130_fd_sc_hd__and2_1
XFILLER_0_74_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08282_ _08302_/A _08281_/B _08270_/X vssd1 vssd1 vccd1 vccd1 _08290_/B sky130_fd_sc_hd__a21oi_2
X_07302_ _07303_/B _07303_/C _07303_/A vssd1 vssd1 vccd1 vccd1 _08305_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_6_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07233_ _07233_/A _07233_/B vssd1 vssd1 vccd1 vccd1 _07234_/B sky130_fd_sc_hd__and2_1
XFILLER_0_116_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07164_ _07164_/A _07384_/A vssd1 vssd1 vccd1 vccd1 _07225_/B sky130_fd_sc_hd__or2_1
XFILLER_0_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07095_ reg1_val[28] _07095_/B vssd1 vssd1 vccd1 vccd1 _07097_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout213 _06785_/X vssd1 vssd1 vccd1 vccd1 _09362_/S sky130_fd_sc_hd__buf_6
Xfanout202 _09109_/Y vssd1 vssd1 vccd1 vccd1 _12223_/B1 sky130_fd_sc_hd__buf_4
Xfanout235 _09384_/X vssd1 vssd1 vccd1 vccd1 _09385_/C sky130_fd_sc_hd__clkbuf_4
Xfanout246 _09114_/Y vssd1 vssd1 vccd1 vccd1 _12373_/A1 sky130_fd_sc_hd__buf_4
XANTENNA__11901__A1 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout224 _06964_/A vssd1 vssd1 vccd1 vccd1 _11089_/A sky130_fd_sc_hd__buf_4
XFILLER_0_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout257 _06881_/Y vssd1 vssd1 vccd1 vccd1 _12487_/S sky130_fd_sc_hd__buf_6
Xfanout268 _13168_/A2 vssd1 vssd1 vccd1 vccd1 _12955_/A2 sky130_fd_sc_hd__buf_4
X_07997_ _07997_/A _07997_/B vssd1 vssd1 vccd1 vccd1 _07998_/B sky130_fd_sc_hd__xnor2_4
Xfanout279 _12658_/A vssd1 vssd1 vccd1 vccd1 _12708_/B sky130_fd_sc_hd__buf_4
X_09805_ _09650_/A _09650_/B _09648_/Y vssd1 vssd1 vccd1 vccd1 _09806_/B sky130_fd_sc_hd__a21boi_4
X_06948_ _06964_/A _10249_/S _09679_/S _08588_/A vssd1 vssd1 vccd1 vccd1 _06951_/C
+ sky130_fd_sc_hd__and4_1
X_09736_ _09736_/A _09736_/B _09736_/C _09736_/D vssd1 vssd1 vccd1 vccd1 _09737_/B
+ sky130_fd_sc_hd__or4_2
X_09667_ _10617_/A _09668_/B _09668_/C vssd1 vssd1 vccd1 vccd1 _09667_/Y sky130_fd_sc_hd__o21ai_1
X_08618_ _09009_/A _08616_/X _09007_/B _08431_/Y vssd1 vssd1 vccd1 vccd1 _09058_/A
+ sky130_fd_sc_hd__a31o_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06879_ _09200_/B _06879_/B vssd1 vssd1 vccd1 vccd1 dest_pred_val sky130_fd_sc_hd__xnor2_4
XANTENNA__07333__A1 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07333__B2 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09598_ _09597_/B _09597_/C _09597_/A vssd1 vssd1 vccd1 vccd1 _09599_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08549_ _08549_/A _08549_/B _08549_/C vssd1 vssd1 vccd1 vccd1 _08559_/A sky130_fd_sc_hd__or3_2
XANTENNA__11417__B1 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11560_ _06865_/B _11470_/B _06676_/A vssd1 vssd1 vccd1 vccd1 _11560_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_107_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10511_ hold198/A _12124_/B _10632_/B _10510_/Y _12290_/C1 vssd1 vssd1 vccd1 vccd1
+ _10511_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13031__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ _13241_/CLK _13230_/D vssd1 vssd1 vccd1 vccd1 hold215/A sky130_fd_sc_hd__dfxtp_1
X_11491_ _09205_/B _11479_/X _11490_/X _11473_/X vssd1 vssd1 vccd1 vccd1 _11491_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09389__A2 _09392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10442_ _10442_/A _10442_/B vssd1 vssd1 vccd1 vccd1 _10445_/A sky130_fd_sc_hd__xor2_2
X_13161_ _13166_/A hold245/X vssd1 vssd1 vccd1 vccd1 _13310_/D sky130_fd_sc_hd__and2_1
X_10373_ _10373_/A _10373_/B vssd1 vssd1 vccd1 vccd1 _10373_/Y sky130_fd_sc_hd__nand2_1
X_13092_ _13092_/A _13092_/B vssd1 vssd1 vccd1 vccd1 _13093_/B sky130_fd_sc_hd__nand2_1
X_12112_ _12053_/A _12050_/Y _12052_/B vssd1 vssd1 vccd1 vccd1 _12112_/X sky130_fd_sc_hd__o21a_1
XANTENNA__08349__A0 _08853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12043_ _06604_/X _11979_/Y _06602_/Y vssd1 vssd1 vccd1 vccd1 _12043_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10156__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12945_ hold209/X _12947_/A2 _12947_/B1 hold183/X vssd1 vssd1 vccd1 vccd1 hold210/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08096__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12876_ hold256/X hold19/X vssd1 vssd1 vccd1 vccd1 _12877_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11827_ reg1_val[22] curr_PC[22] vssd1 vssd1 vccd1 vccd1 _11828_/B sky130_fd_sc_hd__or2_1
XFILLER_0_68_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11408__B1 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11758_ _09115_/X _10629_/X _10642_/Y _09184_/X _11757_/X vssd1 vssd1 vccd1 vccd1
+ _11758_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10709_ _10710_/A _10710_/B vssd1 vssd1 vccd1 vccd1 _10711_/A sky130_fd_sc_hd__or2_1
XFILLER_0_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11689_ _11690_/A _11690_/B vssd1 vssd1 vccd1 vccd1 _11691_/A sky130_fd_sc_hd__or2_1
XFILLER_0_126_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07920_ _07918_/Y _08034_/B _07915_/Y vssd1 vssd1 vccd1 vccd1 _07924_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06998__B _07005_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ _08836_/A _07851_/B vssd1 vssd1 vccd1 vccd1 _07855_/A sky130_fd_sc_hd__xnor2_1
X_07782_ _07782_/A _07782_/B vssd1 vssd1 vccd1 vccd1 _07887_/A sky130_fd_sc_hd__xnor2_4
X_06802_ _06542_/Y _07015_/B _06801_/X vssd1 vssd1 vccd1 vccd1 _06802_/Y sky130_fd_sc_hd__o21ai_1
X_06733_ reg1_val[9] _07324_/A vssd1 vssd1 vccd1 vccd1 _06734_/B sky130_fd_sc_hd__nand2_1
X_09521_ _09128_/X _09133_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09521_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09304__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08512__B1 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11111__A2 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07866__A2 _11147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06664_ reg2_val[19] _06752_/A _06680_/B1 _06663_/Y vssd1 vssd1 vccd1 vccd1 _07077_/A
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__11425__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ _09452_/A _09452_/B vssd1 vssd1 vccd1 vccd1 _09454_/B sky130_fd_sc_hd__xnor2_1
X_08403_ _08403_/A _08403_/B vssd1 vssd1 vccd1 vccd1 _08620_/C sky130_fd_sc_hd__xnor2_1
X_06595_ reg2_val[25] _06752_/A _06688_/B1 _06594_/Y vssd1 vssd1 vccd1 vccd1 _07157_/A
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_93_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09383_ _09383_/A _09383_/B vssd1 vssd1 vccd1 vccd1 _09383_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08334_ _08334_/A _08334_/B vssd1 vssd1 vccd1 vccd1 _08344_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_74_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout245_A _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08265_ _08841_/B2 _08772_/B2 _08772_/A2 _09888_/B2 vssd1 vssd1 vccd1 vccd1 _08266_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07094__A3 _12697_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08196_ _08242_/A _08242_/B _08185_/X vssd1 vssd1 vccd1 vccd1 _08205_/B sky130_fd_sc_hd__a21boi_2
X_07216_ _12250_/A _06837_/B _07128_/X _07135_/B vssd1 vssd1 vccd1 vccd1 _07217_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07147_ _09621_/A _07148_/B vssd1 vssd1 vccd1 vccd1 _07149_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_70_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12375__A1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09565__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07251__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07078_ _07079_/A _07079_/B vssd1 vssd1 vccd1 vccd1 _07078_/X sky130_fd_sc_hd__and2_1
XFILLER_0_100_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06701__B _07192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09543__A2 _09392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10689__A1 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10689__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__A1 _07308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout60_A _07153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13026__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10991_ _10972_/A _09383_/B _10987_/Y _10988_/X _10990_/X vssd1 vssd1 vccd1 vccd1
+ _10991_/X sky130_fd_sc_hd__o221a_1
X_09719_ _09635_/A _09635_/B _09633_/Y vssd1 vssd1 vccd1 vccd1 _09733_/A sky130_fd_sc_hd__a21o_2
XANTENNA__07857__A2 _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_6_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13306_/CLK sky130_fd_sc_hd__clkbuf_8
X_12730_ _12730_/A _12744_/B vssd1 vssd1 vccd1 vccd1 _12730_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ _12661_/A _12661_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[20] sky130_fd_sc_hd__nor2_8
XFILLER_0_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12063__B1 _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11612_/A _11612_/B vssd1 vssd1 vccd1 vccd1 _11613_/B sky130_fd_sc_hd__or2_1
XFILLER_0_65_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11405__A3 _11404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12592_ reg1_val[7] _12593_/B vssd1 vssd1 vccd1 vccd1 _12592_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_80_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11543_ _11544_/A _11544_/B _11544_/C vssd1 vssd1 vccd1 vccd1 _11632_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11474_ reg1_val[18] curr_PC[18] vssd1 vssd1 vccd1 vccd1 _11476_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13213_ _13306_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10425_ _10551_/B _10425_/B vssd1 vssd1 vccd1 vccd1 _10429_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13144_ _13144_/A _13144_/B vssd1 vssd1 vccd1 vccd1 _13144_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__12118__A1 _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12613__B _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10356_ _10356_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10357_/B sky130_fd_sc_hd__xor2_1
X_13075_ hold291/X _12721_/B _13074_/X _12722_/A vssd1 vssd1 vccd1 vccd1 _13076_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ _10527_/A fanout20/X fanout18/X _10452_/B2 vssd1 vssd1 vccd1 vccd1 _10288_/B
+ sky130_fd_sc_hd__o22a_1
X_12026_ _12026_/A _12026_/B vssd1 vssd1 vccd1 vccd1 _12027_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07545__A1 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07545__B2 _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09298__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09298__B2 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12928_ _13166_/A hold208/X vssd1 vssd1 vccd1 vccd1 _13234_/D sky130_fd_sc_hd__and2_1
XFILLER_0_29_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12859_ hold58/X hold258/X vssd1 vssd1 vccd1 vccd1 _13097_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_29_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12054__B1 _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08273__A2 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_3_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08050_ _08050_/A _08050_/B vssd1 vssd1 vccd1 vccd1 _08105_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_43_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07001_ _09968_/A _12370_/B _07001_/C vssd1 vssd1 vccd1 vccd1 _07001_/X sky130_fd_sc_hd__and3_1
XFILLER_0_12_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08025__A2 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08952_ _08950_/A _08950_/B _08953_/B vssd1 vssd1 vccd1 vccd1 _08952_/X sky130_fd_sc_hd__o21ba_1
X_07903_ _08030_/A _08030_/B vssd1 vssd1 vccd1 vccd1 _07907_/A sky130_fd_sc_hd__or2_1
X_08883_ _08883_/A _08883_/B _08883_/C vssd1 vssd1 vccd1 vccd1 _08884_/B sky130_fd_sc_hd__and3_1
XANTENNA_fanout195_A _13151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ _07804_/B _08020_/B _07804_/A vssd1 vssd1 vccd1 vccd1 _07885_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13085__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07765_ _09621_/A _07765_/B vssd1 vssd1 vccd1 vccd1 _07767_/B sky130_fd_sc_hd__xnor2_4
X_06716_ reg2_val[11] _06729_/B vssd1 vssd1 vccd1 vccd1 _06716_/X sky130_fd_sc_hd__and2_1
X_07696_ _07696_/A _07696_/B vssd1 vssd1 vccd1 vccd1 _08966_/A sky130_fd_sc_hd__xnor2_4
X_09504_ _09506_/A _09506_/B vssd1 vssd1 vccd1 vccd1 _09504_/X sky130_fd_sc_hd__or2_1
X_06647_ _06647_/A _06647_/B vssd1 vssd1 vccd1 vccd1 _11824_/A sky130_fd_sc_hd__nor2_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09435_ _09436_/A _09436_/B vssd1 vssd1 vccd1 vccd1 _09435_/Y sky130_fd_sc_hd__nand2_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06578_ instruction[24] _12658_/A _06898_/B instruction[41] _06574_/X vssd1 vssd1
+ vccd1 vccd1 _06579_/B sky130_fd_sc_hd__a221o_1
X_09366_ _09147_/X _09173_/X _12726_/A vssd1 vssd1 vccd1 vccd1 _09366_/X sky130_fd_sc_hd__mux2_1
X_08317_ _08320_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _08317_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_40 reg2_val[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09297_ _09296_/B _09296_/C _10555_/A vssd1 vssd1 vccd1 vccd1 _09302_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08248_ _08297_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08298_/A sky130_fd_sc_hd__nand2_1
XANTENNA_51 reg2_val[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_62 reg2_val[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_84 reg1_val[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_73 reg1_val[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08179_ _08183_/A _08183_/B vssd1 vssd1 vccd1 vccd1 _08179_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_104_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12899__A2 _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10210_ _10077_/A _10076_/B _10074_/Y vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07808__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06578__A2 _12658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ reg1_val[15] curr_PC[15] vssd1 vssd1 vccd1 vccd1 _11191_/B sky130_fd_sc_hd__or2_1
XANTENNA__09295__A _09295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ _10003_/B _10273_/B _10617_/A vssd1 vssd1 vccd1 vccd1 _10141_/Y sky130_fd_sc_hd__a21oi_1
X_10072_ _10072_/A _10072_/B vssd1 vssd1 vccd1 vccd1 _10073_/B sky130_fd_sc_hd__xnor2_2
X_10974_ reg1_val[13] curr_PC[13] vssd1 vssd1 vccd1 vccd1 _10976_/A sky130_fd_sc_hd__nand2_1
Xmax_cap97 _11147_/A vssd1 vssd1 vccd1 vccd1 _07179_/A sky130_fd_sc_hd__buf_6
XFILLER_0_69_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12713_ _12713_/A _12713_/B vssd1 vssd1 vccd1 vccd1 _12714_/B sky130_fd_sc_hd__xnor2_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12644_ _12644_/A _12644_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[16] sky130_fd_sc_hd__xor2_4
XFILLER_0_127_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12575_ _12575_/A _12575_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[3] sky130_fd_sc_hd__xnor2_4
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06606__B _06633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10062__A2 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11526_ _11525_/B _11526_/B vssd1 vssd1 vccd1 vccd1 _11527_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_108_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13000__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08821__B _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11457_ _11457_/A _11457_/B _11457_/C vssd1 vssd1 vccd1 vccd1 _11458_/B sky130_fd_sc_hd__nand3_1
X_11388_ reg1_val[17] curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11389_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07718__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10408_ _10411_/A vssd1 vssd1 vccd1 vccd1 _10408_/Y sky130_fd_sc_hd__inv_2
X_13127_ hold252/X _13126_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13127_/X sky130_fd_sc_hd__mux2_1
X_10339_ _10340_/A _10340_/B vssd1 vssd1 vccd1 vccd1 _10339_/Y sky130_fd_sc_hd__nor2_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _13058_/A _13058_/B vssd1 vssd1 vccd1 vccd1 _13058_/Y sky130_fd_sc_hd__xnor2_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07518__A1 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07518__B2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ _12200_/A _12009_/B vssd1 vssd1 vccd1 vccd1 _12011_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08191__A1 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08191__B2 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06741__A2 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07550_ _10064_/B2 _08680_/B fanout30/X _09888_/B2 vssd1 vssd1 vccd1 vccd1 _07551_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09691__A1 _11194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08494__A2 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09220_ curr_PC[0] _12005_/A vssd1 vssd1 vccd1 vccd1 _09220_/X sky130_fd_sc_hd__or2_1
X_07481_ _07482_/B _07583_/A _07482_/A vssd1 vssd1 vccd1 vccd1 _09316_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_124_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09151_ reg1_val[27] reg1_val[4] _09158_/S vssd1 vssd1 vccd1 vccd1 _09151_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08102_ _08103_/A _08103_/B vssd1 vssd1 vccd1 vccd1 _08102_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_83_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09082_ _09098_/A _09082_/B vssd1 vssd1 vccd1 vccd1 _09082_/X sky130_fd_sc_hd__xor2_1
XANTENNA__10053__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08033_ _08033_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08106_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout208_A _07763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07206__B1 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07757__B2 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07757__A1 _10281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10054__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09984_ hold284/A _09385_/C _09982_/X _11400_/A vssd1 vssd1 vccd1 vccd1 _09984_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10761__B1 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08935_ _08935_/A _08935_/B vssd1 vssd1 vccd1 vccd1 _08935_/X sky130_fd_sc_hd__or2_1
XANTENNA__07509__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__A1 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08866_ _08866_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _08880_/A sky130_fd_sc_hd__xor2_2
XANTENNA__10513__B1 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07817_ _08857_/A _07817_/B vssd1 vssd1 vccd1 vccd1 _07842_/B sky130_fd_sc_hd__xnor2_4
X_08797_ _08798_/A _08798_/B vssd1 vssd1 vccd1 vccd1 _08883_/A sky130_fd_sc_hd__nand2_1
X_07748_ fanout70/X _08692_/A2 _08692_/B1 _12762_/A vssd1 vssd1 vccd1 vccd1 _07749_/B
+ sky130_fd_sc_hd__o22a_1
X_07679_ _08772_/B2 _12766_/A fanout69/X _07058_/A vssd1 vssd1 vccd1 vccd1 _07680_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout23_A _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09418_ _09418_/A _09418_/B _09418_/C vssd1 vssd1 vccd1 vccd1 _09419_/B sky130_fd_sc_hd__nand3_1
X_10690_ _12255_/B _10690_/B vssd1 vssd1 vccd1 vccd1 _10696_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09349_ _09135_/X _09138_/X _09359_/S vssd1 vssd1 vccd1 vccd1 _09349_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09434__A1 _09283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12360_ _12360_/A _12360_/B vssd1 vssd1 vccd1 vccd1 _12360_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10044__A2 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11311_ curr_PC[16] _11314_/C vssd1 vssd1 vccd1 vccd1 _11311_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12291_ reg1_val[29] _09202_/B wire201/A _06583_/X vssd1 vssd1 vccd1 vccd1 _12291_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_50_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11242_ _11119_/A _11119_/B _11115_/X vssd1 vssd1 vccd1 vccd1 _11244_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12741__A1 _10149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__B2 _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__A1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ _11173_/A _11462_/A vssd1 vssd1 vccd1 vccd1 _11374_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_30_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10124_ hold266/A _09385_/C _10256_/B _12339_/B1 vssd1 vssd1 vccd1 vccd1 _10124_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09472__B _09472_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10055_ _10058_/A vssd1 vssd1 vccd1 vccd1 _10147_/A sky130_fd_sc_hd__inv_2
X_10957_ _10958_/A _10958_/B vssd1 vssd1 vccd1 vccd1 _10957_/X sky130_fd_sc_hd__and2_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10888_ curr_PC[12] _10772_/B _10400_/S vssd1 vssd1 vccd1 vccd1 _10888_/Y sky130_fd_sc_hd__o21ai_2
X_12627_ _12635_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _12629_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07436__B1 _06622_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09425__A1 _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09425__B2 _09295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11232__A1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12558_ _12558_/A _12558_/B vssd1 vssd1 vccd1 vccd1 new_PC[27] sky130_fd_sc_hd__xnor2_4
XFILLER_0_81_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08832__A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11232__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12489_ _12490_/A _12490_/B _12490_/C vssd1 vssd1 vccd1 vccd1 _12500_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12980__A1 _10453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold107 hold107/A vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
X_11509_ _11509_/A _11509_/B vssd1 vssd1 vccd1 vccd1 _11510_/B sky130_fd_sc_hd__nor2_1
Xhold118 hold118/A vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _07974_/A _06987_/B vssd1 vssd1 vccd1 vccd1 _09294_/A sky130_fd_sc_hd__xnor2_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11299__B2 _06928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08720_ _08720_/A _08720_/B vssd1 vssd1 vccd1 vccd1 _08805_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09382__B _12726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06962__A2 _09392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _12762_/A _08772_/B2 _08772_/A2 _12760_/A vssd1 vssd1 vccd1 vccd1 _08652_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07911__A1 _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07911__B2 _07869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07602_ _07600_/X _07602_/B vssd1 vssd1 vccd1 vccd1 _07603_/B sky130_fd_sc_hd__and2b_1
X_08582_ _08596_/A _08596_/B vssd1 vssd1 vccd1 vccd1 _08585_/A sky130_fd_sc_hd__nor2_1
X_07533_ _09968_/A _07528_/C reg1_val[29] reg1_val[30] _12713_/A vssd1 vssd1 vccd1
+ vccd1 _12301_/C sky130_fd_sc_hd__a2111o_2
XFILLER_0_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11471__A1 _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout158_A _08681_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07464_ _07464_/A _07464_/B vssd1 vssd1 vccd1 vccd1 _07584_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_119_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09203_ _09180_/A _10377_/B _09198_/X hold211/A vssd1 vssd1 vccd1 vccd1 _09203_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07395_ _09898_/A _07395_/B vssd1 vssd1 vccd1 vccd1 _07396_/C sky130_fd_sc_hd__xor2_1
X_09134_ reg1_val[10] reg1_val[21] _09172_/S vssd1 vssd1 vccd1 vccd1 _09134_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_115_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08742__A _09600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11223__A1 _11222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09065_ _11379_/B _11379_/C _11468_/A vssd1 vssd1 vccd1 vccd1 _11559_/B sky130_fd_sc_hd__nand3_2
X_08016_ _08016_/A _08016_/B vssd1 vssd1 vccd1 vccd1 _08638_/B sky130_fd_sc_hd__xor2_4
XANTENNA__07358__A _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09967_ _06762_/Y _09824_/X _06764_/B vssd1 vssd1 vccd1 vccd1 _09968_/B sky130_fd_sc_hd__o21a_1
X_08918_ _08862_/A _08862_/B _08865_/A vssd1 vssd1 vccd1 vccd1 _08923_/A sky130_fd_sc_hd__a21o_2
XANTENNA__06953__A2 _07087_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08189__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07093__A _09392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09898_ _09898_/A _09898_/B vssd1 vssd1 vccd1 vccd1 _09900_/B sky130_fd_sc_hd__xnor2_1
X_08849_ _08850_/A _08850_/B vssd1 vssd1 vccd1 vccd1 _08849_/X sky130_fd_sc_hd__and2_1
XANTENNA__12239__B1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11860_ _11861_/A _11861_/B vssd1 vssd1 vccd1 vccd1 _11955_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12439__A _12603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07821__A _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11791_ _11791_/A _11791_/B _11791_/C vssd1 vssd1 vccd1 vccd1 _11792_/B sky130_fd_sc_hd__or3_1
X_10811_ _10811_/A _12255_/B _10812_/A vssd1 vssd1 vccd1 vccd1 _10811_/X sky130_fd_sc_hd__and3_1
X_10742_ _06806_/Y _10741_/Y _11738_/S vssd1 vssd1 vccd1 vccd1 _10743_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_67_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09407__A1 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09407__B2 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10673_ _10674_/A _10674_/B vssd1 vssd1 vccd1 vccd1 _10824_/B sky130_fd_sc_hd__and2_1
XFILLER_0_106_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08652__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12412_ _12583_/B _12412_/B vssd1 vssd1 vccd1 vccd1 _12413_/B sky130_fd_sc_hd__or2_1
XANTENNA__11214__A1 _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12962__A1 _07148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12174__A _12174_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12343_ _12319_/Y _12320_/X _12324_/X _12342_/Y vssd1 vssd1 vccd1 vccd1 _12343_/X
+ sky130_fd_sc_hd__o211a_1
X_12274_ _06591_/B _12226_/Y _06591_/A vssd1 vssd1 vccd1 vccd1 _12274_/X sky130_fd_sc_hd__a21bo_1
X_11225_ _11688_/A fanout27/X _12205_/A fanout70/X vssd1 vssd1 vccd1 vccd1 _11226_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11517__A2 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11156_ _11045_/A _11045_/B _11043_/X vssd1 vssd1 vccd1 vccd1 _11156_/Y sky130_fd_sc_hd__a21oi_1
X_11087_ _10978_/A _10978_/B _10976_/A vssd1 vssd1 vccd1 vccd1 _11088_/B sky130_fd_sc_hd__o21a_1
X_10107_ _06796_/X _10106_/Y _12322_/S vssd1 vssd1 vccd1 vccd1 _10108_/B sky130_fd_sc_hd__mux2_1
XANTENNA__11518__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10038_ _10206_/A _10038_/B vssd1 vssd1 vccd1 vccd1 _10040_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_105_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11989_ hold256/A hold293/A _11989_/C vssd1 vssd1 vccd1 vccd1 _12056_/B sky130_fd_sc_hd__or3_1
XFILLER_0_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12349__A _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07180_ _08733_/A _07180_/B vssd1 vssd1 vccd1 vccd1 _07180_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08082__B1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07178__A _07178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09821_ _12278_/A _09821_/B vssd1 vssd1 vccd1 vccd1 _09821_/X sky130_fd_sc_hd__and2_1
XFILLER_0_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09752_ _12762_/A _09752_/B vssd1 vssd1 vccd1 vccd1 _09754_/B sky130_fd_sc_hd__or2_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08137__B2 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08137__A1 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ _08703_/A _08703_/B _08703_/C vssd1 vssd1 vccd1 vccd1 _08705_/A sky130_fd_sc_hd__and3_1
X_06964_ _06964_/A _06964_/B vssd1 vssd1 vccd1 vccd1 _09600_/A sky130_fd_sc_hd__xnor2_4
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11147__B _11147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09683_ _09538_/A _09535_/Y _09537_/B vssd1 vssd1 vccd1 vccd1 _09683_/X sky130_fd_sc_hd__o21a_1
X_06895_ instruction[11] _06897_/B vssd1 vssd1 vccd1 vccd1 dest_pred[0] sky130_fd_sc_hd__and2_4
X_08634_ _08635_/A _08635_/B vssd1 vssd1 vccd1 vccd1 _08634_/X sky130_fd_sc_hd__and2b_1
XANTENNA__08737__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11692__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11692__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _08559_/A _08559_/B _08559_/C vssd1 vssd1 vccd1 vccd1 _08567_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout13 fanout14/X vssd1 vssd1 vccd1 vccd1 fanout13/X sky130_fd_sc_hd__buf_6
XFILLER_0_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07516_ _07516_/A _07516_/B vssd1 vssd1 vccd1 vccd1 _07517_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08496_ _07969_/A _08692_/A2 _09273_/A1 _09772_/A vssd1 vssd1 vccd1 vccd1 _08497_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout46 fanout47/X vssd1 vssd1 vccd1 vccd1 fanout46/X sky130_fd_sc_hd__buf_6
Xfanout24 _07132_/Y vssd1 vssd1 vccd1 vccd1 _12782_/A sky130_fd_sc_hd__buf_8
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout35 fanout36/X vssd1 vssd1 vccd1 vccd1 fanout35/X sky130_fd_sc_hd__buf_6
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout79 _06982_/Y vssd1 vssd1 vccd1 vccd1 _10553_/A sky130_fd_sc_hd__buf_8
Xfanout68 _07090_/X vssd1 vssd1 vccd1 vccd1 _10280_/A sky130_fd_sc_hd__buf_12
Xfanout57 _07179_/Y vssd1 vssd1 vccd1 vccd1 fanout57/X sky130_fd_sc_hd__buf_6
X_07447_ _07447_/A _07447_/B vssd1 vssd1 vccd1 vccd1 _07448_/B sky130_fd_sc_hd__or2_1
X_07378_ _07376_/A _07376_/B _07693_/A vssd1 vssd1 vccd1 vccd1 _07417_/A sky130_fd_sc_hd__a21oi_1
X_09117_ _09180_/A reg1_val[31] _09158_/S vssd1 vssd1 vccd1 vccd1 _09117_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09048_ _10370_/B _10370_/C vssd1 vssd1 vccd1 vccd1 _09048_/X sky130_fd_sc_hd__and2_1
XFILLER_0_102_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12722__A _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08376__B2 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08376__A1 _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ _11431_/A fanout27/X fanout26/X _11347_/A vssd1 vssd1 vccd1 vccd1 _11011_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10183__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11380__B1 _11379_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10183__B2 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ hold1/X _12723_/A _13170_/B hold83/X _13179_/A vssd1 vssd1 vccd1 vccd1 hold84/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA__11132__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12892_ _13167_/A _13167_/C _13167_/B vssd1 vssd1 vccd1 vccd1 hold243/A sky130_fd_sc_hd__o21bai_2
X_11912_ _11912_/A _11912_/B vssd1 vssd1 vccd1 vccd1 _11912_/Y sky130_fd_sc_hd__xnor2_1
X_11843_ _11824_/Y _11825_/X _11831_/X _09205_/B _11842_/X vssd1 vssd1 vccd1 vccd1
+ _11843_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09089__C1 _09079_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07551__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07103__A2 _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11774_ _11773_/B _11774_/B vssd1 vssd1 vccd1 vccd1 _11775_/B sky130_fd_sc_hd__nand2b_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10725_ _10725_/A _10725_/B vssd1 vssd1 vccd1 vccd1 _10728_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08382__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10656_ _12782_/A fanout54/X fanout20/X fanout95/X vssd1 vssd1 vccd1 vccd1 _10657_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06614__B _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10587_ _10587_/A _10587_/B vssd1 vssd1 vccd1 vccd1 _10588_/B sky130_fd_sc_hd__nor2_2
X_12326_ _12326_/A _12326_/B vssd1 vssd1 vccd1 vccd1 _12326_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_51_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12257_ _12257_/A _12257_/B vssd1 vssd1 vccd1 vccd1 _12259_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12188_ hold213/A _12332_/B _12237_/B _12290_/C1 vssd1 vssd1 vccd1 vccd1 _12189_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11208_ _10251_/S _09177_/X _09214_/A vssd1 vssd1 vccd1 vccd1 _11208_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09564__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11139_ _11139_/A _11139_/B vssd1 vssd1 vccd1 vccd1 _11140_/B sky130_fd_sc_hd__nor2_1
X_06680_ reg2_val[17] _06569_/X _06680_/B1 _06679_/Y vssd1 vssd1 vccd1 vccd1 _07049_/C
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__11674__A1 _12345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07342__A2 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07461__A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08350_ _08365_/B vssd1 vssd1 vccd1 vccd1 _08351_/B sky130_fd_sc_hd__inv_2
XFILLER_0_74_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07301_ _11429_/A _11429_/B vssd1 vssd1 vccd1 vccd1 _07301_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_19_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08281_ _08270_/X _08281_/B vssd1 vssd1 vccd1 vccd1 _08302_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10634__C1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07232_ _07233_/A _07233_/B vssd1 vssd1 vccd1 vccd1 _07234_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_116_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07163_ _07383_/A _07383_/B _07383_/C vssd1 vssd1 vccd1 vccd1 _07384_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07094_ _07087_/B _07087_/C _12697_/B _07165_/A vssd1 vssd1 vccd1 vccd1 _07095_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_42_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07636__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout203 _08311_/A vssd1 vssd1 vccd1 vccd1 _08589_/A sky130_fd_sc_hd__buf_8
Xfanout214 _08821_/A vssd1 vssd1 vccd1 vccd1 _08588_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__06540__A _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout236 _10377_/B vssd1 vssd1 vccd1 vccd1 _11099_/B sky130_fd_sc_hd__buf_4
Xfanout225 _06761_/Y vssd1 vssd1 vccd1 vccd1 _10752_/S sky130_fd_sc_hd__clkbuf_8
Xfanout247 _07869_/B vssd1 vssd1 vccd1 vccd1 _08758_/A2 sky130_fd_sc_hd__buf_6
XFILLER_0_5_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09804_ _09804_/A _09804_/B vssd1 vssd1 vccd1 vccd1 _09806_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_10_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout269 _13168_/A2 vssd1 vssd1 vccd1 vccd1 _13146_/B2 sky130_fd_sc_hd__buf_4
X_07996_ _07997_/A _07997_/B vssd1 vssd1 vccd1 vccd1 _07996_/X sky130_fd_sc_hd__and2b_1
Xfanout258 _12345_/A vssd1 vssd1 vccd1 vccd1 _10400_/S sky130_fd_sc_hd__clkbuf_16
X_06947_ _11823_/S _12370_/B vssd1 vssd1 vccd1 vccd1 _07075_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09851__A _12284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09858__A1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ _09736_/A _09736_/B _09736_/C _09736_/D vssd1 vssd1 vccd1 vccd1 _09735_/X
+ sky130_fd_sc_hd__o22a_1
X_09666_ _09666_/A _10273_/C vssd1 vssd1 vccd1 vccd1 _09666_/Y sky130_fd_sc_hd__nand2_1
X_08617_ _09008_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _09007_/B sky130_fd_sc_hd__nand2_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06878_ instruction[3] _06860_/X _06872_/X _09200_/C _06874_/X vssd1 vssd1 vccd1
+ vccd1 _06879_/B sky130_fd_sc_hd__a221o_2
XANTENNA__07333__A2 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ _09597_/A _09597_/B _09597_/C vssd1 vssd1 vccd1 vccd1 _09599_/A sky130_fd_sc_hd__and3_1
XFILLER_0_77_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08548_ _08589_/A _08548_/B vssd1 vssd1 vccd1 vccd1 _08549_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__11417__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11417__A1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08479_ _08506_/A _08506_/B vssd1 vssd1 vccd1 vccd1 _08489_/A sky130_fd_sc_hd__and2b_1
X_11490_ _11490_/A _11490_/B _11490_/C vssd1 vssd1 vccd1 vccd1 _11490_/X sky130_fd_sc_hd__and3_1
XFILLER_0_92_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10640__A2 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10510_ _12124_/B _10632_/B hold198/A vssd1 vssd1 vccd1 vccd1 _10510_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ _10442_/A _10442_/B vssd1 vssd1 vccd1 vccd1 _10441_/X sky130_fd_sc_hd__and2_1
XFILLER_0_17_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09389__A3 wire201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13160_ hold244/X _13165_/A2 _13159_/X _13168_/A2 vssd1 vssd1 vccd1 vccd1 hold245/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10372_ _06801_/B _10371_/Y _11738_/S vssd1 vssd1 vccd1 vccd1 _10373_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_33_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13091_ _13166_/A hold283/X vssd1 vssd1 vccd1 vccd1 _13295_/D sky130_fd_sc_hd__and2_1
X_12111_ _06620_/B _12109_/X _12110_/Y vssd1 vssd1 vccd1 vccd1 _12111_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09546__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ _12007_/X _12072_/B _12041_/Y vssd1 vssd1 vccd1 vccd1 _12042_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07546__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 hold290/A vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10156__A1 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10156__B2 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11656__A1 _11746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ _12946_/A hold174/X vssd1 vssd1 vccd1 vccd1 hold175/A sky130_fd_sc_hd__and2_1
XFILLER_0_99_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08377__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07281__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ _13130_/A _13131_/A _13130_/B vssd1 vssd1 vccd1 vccd1 _13135_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__10864__C1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ reg1_val[22] curr_PC[22] vssd1 vssd1 vccd1 vccd1 _11828_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11408__A1 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11408__B2 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ reg1_val[21] _11099_/B _11755_/X _06660_/B _11756_/Y vssd1 vssd1 vccd1 vccd1
+ _11757_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_448 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10708_ _10708_/A _10708_/B vssd1 vssd1 vccd1 vccd1 _10710_/B sky130_fd_sc_hd__xnor2_1
X_11688_ _11688_/A _12304_/B _11610_/A vssd1 vssd1 vccd1 vccd1 _11690_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_113_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10639_ _07318_/A _11923_/A2 _11099_/B reg1_val[10] _10638_/Y vssd1 vssd1 vccd1 vccd1
+ _10639_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_51_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11250__B _11250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09785__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12309_ _12308_/A _12308_/B _12308_/C vssd1 vssd1 vccd1 vccd1 _12309_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11592__B1 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13289_ _13289_/CLK _13289_/D vssd1 vssd1 vccd1 vccd1 hold268/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07456__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07850_ _12734_/A _08134_/B fanout51/X _09478_/B2 vssd1 vssd1 vccd1 vccd1 _07851_/B
+ sky130_fd_sc_hd__o22a_1
X_07781_ _07781_/A _07781_/B vssd1 vssd1 vccd1 vccd1 _07782_/B sky130_fd_sc_hd__xnor2_4
X_06801_ _10373_/A _06801_/B vssd1 vssd1 vccd1 vccd1 _06801_/X sky130_fd_sc_hd__or2_1
X_06732_ reg1_val[9] _07324_/A vssd1 vssd1 vccd1 vccd1 _06732_/Y sky130_fd_sc_hd__nor2_1
X_09520_ _09121_/X _09125_/X _09676_/S vssd1 vssd1 vccd1 vccd1 _09520_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07191__A _07192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08512__A1 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08512__B2 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06663_ _06687_/A _12578_/B vssd1 vssd1 vccd1 vccd1 _06663_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09451_ _10156_/B2 _10677_/A fanout58/X _10156_/A1 vssd1 vssd1 vccd1 vccd1 _09452_/B
+ sky130_fd_sc_hd__o22a_1
X_08402_ _08430_/A _08430_/B vssd1 vssd1 vccd1 vccd1 _08620_/B sky130_fd_sc_hd__and2_1
X_06594_ _06687_/A _12607_/B vssd1 vssd1 vccd1 vccd1 _06594_/Y sky130_fd_sc_hd__nor2_1
X_09382_ _11823_/S _12726_/A _09382_/C vssd1 vssd1 vccd1 vccd1 _09382_/X sky130_fd_sc_hd__or3_1
XFILLER_0_47_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08333_ _08360_/A _08330_/B _08372_/A vssd1 vssd1 vccd1 vccd1 _08344_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__08276__B1 _08672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08264_ _08264_/A _08264_/B vssd1 vssd1 vccd1 vccd1 _08290_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__13132__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout238_A _09201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout140_A _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08195_ _08244_/A _08195_/B vssd1 vssd1 vccd1 vccd1 _08242_/B sky130_fd_sc_hd__xor2_1
X_07215_ _09467_/A _07215_/B vssd1 vssd1 vccd1 vccd1 _07221_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07146_ _08695_/A _07148_/B vssd1 vssd1 vccd1 vccd1 _07150_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07077_ _07077_/A _07077_/B _07077_/C vssd1 vssd1 vccd1 vccd1 _07079_/B sky130_fd_sc_hd__or3_2
XANTENNA__07251__A1 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07251__B2 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12127__A2 wire201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10689__A2 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__A2 _07308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07979_ _08658_/A _07978_/C _07978_/A vssd1 vssd1 vccd1 vccd1 _07980_/C sky130_fd_sc_hd__a21oi_1
X_09718_ _09651_/A _09651_/B _09652_/Y vssd1 vssd1 vccd1 vccd1 _09811_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_97_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10990_ _06710_/B _09188_/X _09191_/X _06708_/Y _10989_/X vssd1 vssd1 vccd1 vccd1
+ _10990_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_93_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout53_A _07260_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09649_ _09649_/A _09649_/B vssd1 vssd1 vccd1 vccd1 _09650_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _12678_/A _12660_/B _12660_/C vssd1 vssd1 vccd1 vccd1 _12661_/B sky130_fd_sc_hd__and3_2
XANTENNA__08267__B1 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12063__A1 _07157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11611_ _11612_/A _11612_/B vssd1 vssd1 vccd1 vccd1 _11613_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12447__A _12607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12591_ _12590_/A _12589_/A _12589_/B vssd1 vssd1 vccd1 vccd1 _12595_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_53_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11542_ _11542_/A _11542_/B vssd1 vssd1 vccd1 vccd1 _11544_/C sky130_fd_sc_hd__xor2_1
X_11473_ _06865_/B _11471_/Y _11472_/Y vssd1 vssd1 vccd1 vccd1 _11473_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13212_ _13306_/CLK _13212_/D vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08660__A _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10424_ _07278_/B fanout81/X _09295_/B fanout7/X vssd1 vssd1 vccd1 vccd1 _10425_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13143_ _13147_/A _13143_/B vssd1 vssd1 vccd1 vccd1 _13306_/D sky130_fd_sc_hd__and2_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10355_ _10356_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10355_/X sky130_fd_sc_hd__or2_1
X_13074_ hold276/X _13073_/Y hold243/X vssd1 vssd1 vccd1 vccd1 _13074_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10286_ _10158_/A _10158_/B _10154_/X vssd1 vssd1 vccd1 vccd1 _10295_/A sky130_fd_sc_hd__o21ba_1
X_12025_ _12025_/A _12025_/B _12025_/C vssd1 vssd1 vccd1 vccd1 _12026_/B sky130_fd_sc_hd__and3_1
XANTENNA__07545__A2 _09295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06753__B1 _12284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09298__A2 _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12927_ hold207/X _13146_/B2 _13165_/A2 hold178/X vssd1 vssd1 vccd1 vccd1 hold208/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12858_ _13092_/A _13093_/A _13092_/B vssd1 vssd1 vccd1 vccd1 _13098_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_87_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11809_ _11809_/A _11809_/B _11809_/C vssd1 vssd1 vccd1 vccd1 _11810_/B sky130_fd_sc_hd__and3_1
X_12789_ _07435_/Y _13020_/B2 hold76/X _13086_/A vssd1 vssd1 vccd1 vccd1 _13216_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09470__A2 _07435_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07000_ _07000_/A _11933_/A vssd1 vssd1 vccd1 vccd1 _07000_/X sky130_fd_sc_hd__or2_4
XFILLER_0_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08951_ _08910_/A _08910_/C _08910_/B vssd1 vssd1 vccd1 vccd1 _08953_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_11_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07902_ _09452_/A _07902_/B vssd1 vssd1 vccd1 vccd1 _08030_/B sky130_fd_sc_hd__xnor2_2
X_08882_ _08883_/A _08883_/B _08883_/C vssd1 vssd1 vccd1 vccd1 _08884_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__07914__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07833_ _07833_/A _07833_/B vssd1 vssd1 vccd1 vccd1 _08020_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09930__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13127__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _07134_/A fanout77/X _12768_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07765_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_79_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06715_ _06713_/Y _06715_/B vssd1 vssd1 vccd1 vccd1 _10863_/A sky130_fd_sc_hd__nand2b_2
X_07695_ _07697_/A _07697_/B vssd1 vssd1 vccd1 vccd1 _07695_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12293__A1 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09503_ _09503_/A _09503_/B vssd1 vssd1 vccd1 vccd1 _09506_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06646_ reg1_val[22] _07112_/B vssd1 vssd1 vccd1 vccd1 _06647_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_66_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09434_ _09283_/A _09775_/A _09289_/B _09287_/X vssd1 vssd1 vccd1 vccd1 _09436_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06577_ instruction[41] _06898_/B _06574_/X vssd1 vssd1 vccd1 vccd1 _06577_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10056__B1 _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09365_ _09170_/X _09172_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09365_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08316_ _10453_/A _08316_/B vssd1 vssd1 vccd1 vccd1 _08320_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_41 reg2_val[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 reg1_val[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ _10555_/A _09296_/B _09296_/C vssd1 vssd1 vccd1 vccd1 _09302_/A sky130_fd_sc_hd__and3_1
X_08247_ _08247_/A _08247_/B vssd1 vssd1 vccd1 vccd1 _08297_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_52 reg2_val[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 reg2_val[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_74 reg1_val[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_85 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08178_ _08394_/A _08178_/B vssd1 vssd1 vccd1 vccd1 _08183_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11556__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07129_ _07153_/A _07129_/B _07129_/C _07129_/D vssd1 vssd1 vccd1 vccd1 _07434_/C
+ sky130_fd_sc_hd__or4_1
XANTENNA__09295__B _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07096__A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10140_ _10397_/C _10139_/Y _10137_/X vssd1 vssd1 vccd1 vccd1 dest_val[6] sky130_fd_sc_hd__o21ai_4
XFILLER_0_30_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07965__A2_N _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ _10071_/A _10071_/B vssd1 vssd1 vccd1 vccd1 _10072_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__12730__A _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07824__A _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap10 _07435_/Y vssd1 vssd1 vccd1 vccd1 _12349_/A sky130_fd_sc_hd__buf_6
XANTENNA__11346__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07035__S _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10973_ _10972_/A _10972_/B _10972_/Y _12277_/B1 vssd1 vssd1 vccd1 vccd1 _10973_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11492__C1 _11466_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12712_ _12709_/B _12711_/B _12707_/X vssd1 vssd1 vccd1 vccd1 _12713_/B sky130_fd_sc_hd__a21oi_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12643_ _12644_/A _12644_/B vssd1 vssd1 vccd1 vccd1 _12657_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_92_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12574_ _12572_/Y _12574_/B vssd1 vssd1 vccd1 vccd1 _12575_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_25_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11525_ _11526_/B _11525_/B vssd1 vssd1 vccd1 vccd1 _11616_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11456_ _11457_/A _11457_/B _11457_/C vssd1 vssd1 vccd1 vccd1 _11456_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11387_ reg1_val[17] curr_PC[17] vssd1 vssd1 vccd1 vccd1 _11387_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_68_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10407_ _11499_/A _10407_/B vssd1 vssd1 vccd1 vccd1 _10411_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10425__A _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13126_ _13126_/A _13126_/B vssd1 vssd1 vccd1 vccd1 _13126_/Y sky130_fd_sc_hd__xnor2_1
X_10338_ _10150_/A _10150_/B _10148_/A vssd1 vssd1 vccd1 vccd1 _10340_/B sky130_fd_sc_hd__o21a_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13057_/A _13057_/B vssd1 vssd1 vccd1 vccd1 _13058_/B sky130_fd_sc_hd__nand2_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _10269_/A _10269_/B _10269_/C _10269_/D vssd1 vssd1 vccd1 vccd1 _10269_/X
+ sky130_fd_sc_hd__or4_2
XANTENNA__07518__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ _12150_/A fanout15/X fanout6/X _12150_/B vssd1 vssd1 vccd1 vccd1 _12009_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10522__A1 _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08191__A2 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06741__A3 _12598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07480_ _07582_/A _07582_/B vssd1 vssd1 vccd1 vccd1 _07583_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09160__S _09392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12087__A _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09150_ reg1_val[26] reg1_val[5] _09158_/S vssd1 vssd1 vccd1 vccd1 _09150_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08101_ _08099_/A _08099_/B _08155_/A vssd1 vssd1 vccd1 vccd1 _08123_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__08651__B1 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09081_ _09098_/A _09082_/B vssd1 vssd1 vccd1 vccd1 _12133_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_44_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08032_ _08033_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08032_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_32_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07206__A1 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07206__B2 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07757__A2 _07182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09983_ _09842_/B _09982_/X hold284/A vssd1 vssd1 vccd1 vccd1 _09983_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08934_ _08932_/A _08932_/B _08884_/A vssd1 vssd1 vccd1 vccd1 _08935_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09903__B1 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07509__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ _08865_/A _08865_/B vssd1 vssd1 vccd1 vccd1 _08866_/B sky130_fd_sc_hd__nor2_1
X_07816_ _08837_/B2 _08217_/B fanout55/X _07969_/A vssd1 vssd1 vccd1 vccd1 _07817_/B
+ sky130_fd_sc_hd__o22a_2
X_08796_ _08796_/A _08796_/B vssd1 vssd1 vccd1 vccd1 _08798_/B sky130_fd_sc_hd__xnor2_2
X_07747_ _07747_/A _07747_/B _07747_/C vssd1 vssd1 vccd1 vccd1 _07751_/A sky130_fd_sc_hd__and3_1
XANTENNA__07390__B1 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10277__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07678_ _07678_/A _07678_/B _07678_/C vssd1 vssd1 vccd1 vccd1 _07686_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_66_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06629_ reg1_val[30] _07434_/B vssd1 vssd1 vccd1 vccd1 _06631_/A sky130_fd_sc_hd__and2_1
X_09417_ _09418_/A _09418_/B _09418_/C vssd1 vssd1 vccd1 vccd1 _09645_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_118_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09348_ _09132_/X _09134_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09348_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_124_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout16_A _07277_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09434__A2 _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11310_ curr_PC[16] _11314_/C vssd1 vssd1 vccd1 vccd1 _11310_/Y sky130_fd_sc_hd__nand2_1
X_09279_ _09620_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _09280_/B sky130_fd_sc_hd__xnor2_4
X_12290_ _13246_/Q _12332_/B _12330_/B _12289_/Y _12290_/C1 vssd1 vssd1 vccd1 vccd1
+ _12295_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11241_ _11328_/A _11328_/B vssd1 vssd1 vccd1 vccd1 _11244_/A sky130_fd_sc_hd__xor2_1
XANTENNA__12741__A2 _12980_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07748__A2 _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11172_ _11170_/Y _11172_/B vssd1 vssd1 vccd1 vccd1 _11462_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10123_ _09385_/C _10256_/B hold266/A vssd1 vssd1 vccd1 vccd1 _10123_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12460__A _12620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ _10458_/A _10054_/B vssd1 vssd1 vccd1 vccd1 _10058_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12619__B _12620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10956_ _10958_/A _10958_/B vssd1 vssd1 vccd1 vccd1 _10956_/X sky130_fd_sc_hd__or2_1
XFILLER_0_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10887_ curr_PC[11] curr_PC[12] _10887_/C vssd1 vssd1 vccd1 vccd1 _11107_/C sky130_fd_sc_hd__and3_2
XFILLER_0_85_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12626_ reg1_val[13] _12626_/B vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__or2_1
XFILLER_0_66_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07436__A1 _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09425__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12557_ _12557_/A _12557_/B vssd1 vssd1 vccd1 vccd1 _12558_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11232__A2 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12980__A2 _12980_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12488_ _12551_/A _12488_/B vssd1 vssd1 vccd1 vccd1 _12490_/C sky130_fd_sc_hd__xnor2_1
Xhold108 hold108/A vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11508_ _11509_/A _11509_/B vssd1 vssd1 vccd1 vccd1 _11618_/C sky130_fd_sc_hd__and2_1
XFILLER_0_22_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09189__A1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11439_ _11439_/A _11439_/B vssd1 vssd1 vccd1 vccd1 _11453_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10155__A _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13109_ hold260/X _13108_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13109_/X sky130_fd_sc_hd__mux2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11940__B1 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06980_ reg1_val[22] _06980_/B vssd1 vssd1 vccd1 vccd1 _06987_/B sky130_fd_sc_hd__xor2_4
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06962__A3 _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08650_ _08650_/A _08650_/B vssd1 vssd1 vccd1 vccd1 _08654_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07911__A2 _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07601_ _07601_/A _07601_/B _07601_/C vssd1 vssd1 vccd1 vccd1 _07602_/B sky130_fd_sc_hd__or3_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08581_ _08589_/A _08581_/B vssd1 vssd1 vccd1 vccd1 _08596_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07532_ _07441_/A _07441_/B _07439_/Y vssd1 vssd1 vccd1 vccd1 _07538_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_48_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07463_ _07463_/A vssd1 vssd1 vccd1 vccd1 _07584_/A sky130_fd_sc_hd__inv_2
XFILLER_0_64_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09202_ _09202_/A _09202_/B vssd1 vssd1 vccd1 vccd1 _09202_/X sky130_fd_sc_hd__or2_1
XFILLER_0_29_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07394_ fanout77/X _09618_/A1 fanout62/X _09618_/B2 vssd1 vssd1 vccd1 vccd1 _07395_/B
+ sky130_fd_sc_hd__o22a_1
X_09133_ _09131_/X _09132_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09133_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08742__B _09294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11223__A2 _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09064_ _09070_/A _09064_/B vssd1 vssd1 vccd1 vccd1 _11468_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_71_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07639__A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08015_ _08016_/A _08016_/B vssd1 vssd1 vccd1 vccd1 _08806_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10065__A _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07060__C1 _07052_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _10617_/A _09966_/B _09966_/C vssd1 vssd1 vccd1 vccd1 _09966_/X sky130_fd_sc_hd__or3_1
X_08917_ _08866_/A _08866_/B _08849_/X vssd1 vssd1 vccd1 vccd1 _08927_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07374__A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09897_ _09898_/B vssd1 vssd1 vccd1 vccd1 _09897_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_99_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08848_ _08848_/A _08848_/B vssd1 vssd1 vccd1 vccd1 _08850_/B sky130_fd_sc_hd__xnor2_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07363__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ _08779_/A _08779_/B vssd1 vssd1 vccd1 vccd1 _08780_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11790_ _11791_/A _11791_/B _11791_/C vssd1 vssd1 vccd1 vccd1 _11878_/A sky130_fd_sc_hd__o21ai_1
X_10810_ _10811_/A _12255_/B vssd1 vssd1 vccd1 vccd1 _10812_/B sky130_fd_sc_hd__nand2_1
X_10741_ _10621_/A _10619_/X _06728_/B vssd1 vssd1 vccd1 vccd1 _10741_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12411_ _12583_/B _12412_/B vssd1 vssd1 vccd1 vccd1 _12422_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08933__A _09077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09407__A2 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10672_ _11780_/A _10672_/B vssd1 vssd1 vccd1 vccd1 _10674_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12962__A2 _12742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12342_ _09851_/B _12329_/X _12341_/X vssd1 vssd1 vccd1 vccd1 _12342_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10422__B1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12273_ _12317_/B _12272_/B _09110_/X vssd1 vssd1 vccd1 vccd1 _12273_/X sky130_fd_sc_hd__a21o_1
X_11224_ _11224_/A _11224_/B vssd1 vssd1 vccd1 vccd1 _11257_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_120_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11155_ _11007_/A _11007_/B _11006_/A vssd1 vssd1 vccd1 vccd1 _11160_/A sky130_fd_sc_hd__a21o_1
X_11086_ _11086_/A _11086_/B vssd1 vssd1 vccd1 vccd1 _11088_/A sky130_fd_sc_hd__nand2_1
X_10106_ _06755_/Y _09968_/B _06758_/B vssd1 vssd1 vccd1 vccd1 _10106_/Y sky130_fd_sc_hd__o21ai_1
X_10037_ _10037_/A _10037_/B _10037_/C vssd1 vssd1 vccd1 vccd1 _10038_/B sky130_fd_sc_hd__and3_1
XFILLER_0_98_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11988_ _10245_/X _11987_/Y _12361_/B vssd1 vssd1 vccd1 vccd1 _11988_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08854__B1 _07179_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12349__B _12349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10939_ _10827_/A _10827_/B _10816_/A vssd1 vssd1 vccd1 vccd1 _10949_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11205__A2 _09188_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12609_ _12605_/A _12609_/B vssd1 vssd1 vccd1 vccd1 _12611_/C sky130_fd_sc_hd__nand2b_1
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08082__B2 _08774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08082__A1 _08774_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12953__A2 _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09820_ _09716_/X _10002_/B _09819_/Y vssd1 vssd1 vccd1 vccd1 _09820_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07194__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06963_ _11194_/S _06964_/B vssd1 vssd1 vccd1 vccd1 _06963_/Y sky130_fd_sc_hd__xnor2_2
X_09751_ _11125_/A _09751_/B vssd1 vssd1 vccd1 vccd1 _09757_/A sky130_fd_sc_hd__xnor2_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08137__A2 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08702_ _08701_/A _08701_/B _08701_/C vssd1 vssd1 vccd1 vccd1 _08703_/C sky130_fd_sc_hd__o21ai_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06894_ instruction[2] instruction[1] pred_val instruction[0] vssd1 vssd1 vccd1 vccd1
+ _06897_/B sky130_fd_sc_hd__and4b_4
X_09682_ _09675_/X _09681_/X _10251_/S vssd1 vssd1 vccd1 vccd1 _09682_/X sky130_fd_sc_hd__mux2_2
XANTENNA__07345__B1 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ _08633_/A _08633_/B vssd1 vssd1 vccd1 vccd1 _08633_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07922__A _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout170_A _07047_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11692__A2 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08564_ _08570_/A _08570_/B vssd1 vssd1 vccd1 vccd1 _08567_/B sky130_fd_sc_hd__or2_1
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07515_ _07516_/A _07516_/B vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__or2_1
XFILLER_0_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout14 _07308_/X vssd1 vssd1 vccd1 vccd1 fanout14/X sky130_fd_sc_hd__buf_6
X_08495_ _09621_/A _08495_/B vssd1 vssd1 vccd1 vccd1 _08528_/A sky130_fd_sc_hd__xnor2_1
Xfanout47 _07852_/B vssd1 vssd1 vccd1 vccd1 fanout47/X sky130_fd_sc_hd__buf_8
Xfanout25 fanout26/X vssd1 vssd1 vccd1 vccd1 _12205_/A sky130_fd_sc_hd__buf_6
Xfanout36 _06966_/Y vssd1 vssd1 vccd1 vccd1 fanout36/X sky130_fd_sc_hd__buf_6
XFILLER_0_91_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout69 fanout70/X vssd1 vssd1 vccd1 vccd1 fanout69/X sky130_fd_sc_hd__buf_8
XFILLER_0_76_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout58 _07157_/Y vssd1 vssd1 vccd1 vccd1 fanout58/X sky130_fd_sc_hd__buf_6
XFILLER_0_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07446_ _07447_/A _07447_/B vssd1 vssd1 vccd1 vccd1 _07448_/A sky130_fd_sc_hd__nand2_1
X_07377_ _07692_/B _07377_/B vssd1 vssd1 vccd1 vccd1 _07693_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_45_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07369__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09116_ _12563_/A reg1_val[30] _09158_/S vssd1 vssd1 vccd1 vccd1 _09116_/X sky130_fd_sc_hd__mux2_1
XANTENNA__06623__A2 _06898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09047_ _09047_/A _09047_/B vssd1 vssd1 vccd1 vccd1 _10370_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08376__A2 _08774_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11380__A1 _11379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout83_A _07305_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ _09804_/A _09804_/B _09802_/Y vssd1 vssd1 vccd1 vccd1 _09950_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__10183__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12960_ hold1/X _13170_/B _08394_/A _12980_/A2 _12959_/Y vssd1 vssd1 vccd1 vccd1
+ hold2/A sky130_fd_sc_hd__o221a_1
XANTENNA__07336__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11132__A1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11132__B2 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12891_ hold75/X _12891_/B _12891_/C vssd1 vssd1 vccd1 vccd1 _13167_/C sky130_fd_sc_hd__and3_1
X_11911_ _11830_/A _11830_/B _11828_/A vssd1 vssd1 vccd1 vccd1 _11912_/B sky130_fd_sc_hd__o21a_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _11836_/Y _11837_/X _11841_/X _11834_/X vssd1 vssd1 vccd1 vccd1 _11842_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__09089__B1 _09079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10891__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11773_ _11774_/B _11773_/B vssd1 vssd1 vccd1 vccd1 _11864_/A sky130_fd_sc_hd__nand2b_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10724_ _10724_/A _10724_/B vssd1 vssd1 vccd1 vccd1 _10725_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10655_ _10894_/A _10655_/B vssd1 vssd1 vccd1 vccd1 _10660_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07279__A _07279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12325_ _12278_/B _12279_/A _12278_/A vssd1 vssd1 vccd1 vccd1 _12326_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_51_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10586_ _10586_/A _10586_/B _10586_/C vssd1 vssd1 vccd1 vccd1 _10587_/B sky130_fd_sc_hd__and3_1
XFILLER_0_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12256_ fanout19/X _12255_/Y _12254_/Y vssd1 vssd1 vccd1 vccd1 _12257_/B sky130_fd_sc_hd__o21a_1
XANTENNA__12632__B _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11207_ _11400_/A _11199_/X _11200_/Y _11206_/X vssd1 vssd1 vccd1 vccd1 _11207_/X
+ sky130_fd_sc_hd__o31a_1
X_12187_ _12187_/A1 _12237_/B hold213/A vssd1 vssd1 vccd1 vccd1 _12189_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__09564__B2 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09564__A1 _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10433__A _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11138_ _11139_/A _11139_/B vssd1 vssd1 vccd1 vccd1 _11262_/C sky130_fd_sc_hd__and2_1
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08838__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12320__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11069_ _10959_/B _10956_/X _10957_/X vssd1 vssd1 vccd1 vccd1 _11069_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07300_ reg1_val[18] _07300_/B vssd1 vssd1 vccd1 vccd1 _11429_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08280_ _10819_/A _08329_/A vssd1 vssd1 vccd1 vccd1 _08281_/B sky130_fd_sc_hd__or2_1
XFILLER_0_41_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07231_ _10658_/A _07231_/B vssd1 vssd1 vccd1 vccd1 _07233_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07162_ _07162_/A _07162_/B vssd1 vssd1 vccd1 vccd1 _07383_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07093_ _09392_/S _07093_/B vssd1 vssd1 vccd1 vccd1 _07093_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07917__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout204 _08311_/A vssd1 vssd1 vccd1 vccd1 _09622_/A sky130_fd_sc_hd__buf_8
Xfanout226 _07001_/C vssd1 vssd1 vccd1 vccd1 _10251_/S sky130_fd_sc_hd__clkbuf_8
Xfanout237 _09202_/X vssd1 vssd1 vccd1 vccd1 _10377_/B sky130_fd_sc_hd__buf_4
Xfanout215 _12726_/A vssd1 vssd1 vccd1 vccd1 _08821_/A sky130_fd_sc_hd__buf_8
XFILLER_0_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09803_ _09803_/A _09803_/B vssd1 vssd1 vccd1 vccd1 _09804_/B sky130_fd_sc_hd__xor2_4
X_07995_ _07995_/A _07995_/B vssd1 vssd1 vccd1 vccd1 _07997_/B sky130_fd_sc_hd__xnor2_4
Xfanout259 _06898_/C vssd1 vssd1 vccd1 vccd1 _12345_/A sky130_fd_sc_hd__buf_8
XFILLER_0_66_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout248 _09621_/A vssd1 vssd1 vccd1 vccd1 _08595_/A sky130_fd_sc_hd__buf_12
XANTENNA__09307__A1 _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06946_ _11823_/S _12370_/B vssd1 vssd1 vccd1 vccd1 _06946_/X sky130_fd_sc_hd__and2_1
XANTENNA__09851__B _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09734_ _09632_/A _09632_/B _09629_/A vssd1 vssd1 vccd1 vccd1 _09738_/A sky130_fd_sc_hd__o21ai_4
X_06877_ instruction[4] _09198_/B vssd1 vssd1 vccd1 vccd1 _09188_/C sky130_fd_sc_hd__or2_2
X_09665_ _09666_/A _10273_/C vssd1 vssd1 vccd1 vccd1 _09665_/X sky130_fd_sc_hd__or2_1
X_08616_ _08611_/X _08613_/X _09055_/A _08486_/Y vssd1 vssd1 vccd1 vccd1 _08616_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09596_ _09596_/A _09596_/B _09596_/C _09596_/D vssd1 vssd1 vccd1 vccd1 _09597_/C
+ sky130_fd_sc_hd__or4_2
X_08547_ _09478_/B2 _08588_/B _09273_/A1 _09476_/A vssd1 vssd1 vccd1 vccd1 _08548_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11417__A2 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08478_ _08777_/A _08478_/B vssd1 vssd1 vccd1 vccd1 _08506_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07429_ _12782_/A _09273_/A1 fanout20/X _08588_/B vssd1 vssd1 vccd1 vccd1 _07430_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12378__A0 _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11430__A1_N _07308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10440_ _11604_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10442_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10371_ _06742_/Y _10240_/Y _06744_/B vssd1 vssd1 vccd1 vccd1 _10371_/Y sky130_fd_sc_hd__o21ai_1
X_13090_ hold282/X _13165_/A2 _13089_/X _13168_/A2 vssd1 vssd1 vccd1 vccd1 hold283/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07827__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12110_ _06620_/B _12109_/X _12277_/B1 vssd1 vssd1 vccd1 vccd1 _12110_/Y sky130_fd_sc_hd__a21oi_1
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12041_ _12007_/X _12072_/B _12223_/B1 vssd1 vssd1 vccd1 vccd1 _12041_/Y sky130_fd_sc_hd__o21ai_1
Xhold291 hold291/A vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10156__A2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11105__B2 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12943_ hold173/X _12947_/A2 _12947_/B1 hold209/A vssd1 vssd1 vccd1 vccd1 hold174/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12302__B1 _12349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12874_ hold15/X hold293/A vssd1 vssd1 vccd1 vccd1 _13130_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ _11824_/A _11824_/B _09193_/X vssd1 vssd1 vccd1 vccd1 _11825_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_68_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11408__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11756_ _11756_/A wire201/X vssd1 vssd1 vccd1 vccd1 _11756_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_126_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ _10707_/A _10707_/B vssd1 vssd1 vccd1 vccd1 _10708_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06625__B _06633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12369__B1 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11687_ _11777_/B _11687_/B vssd1 vssd1 vccd1 vccd1 _11690_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10638_ _10638_/A _10638_/B vssd1 vssd1 vccd1 vccd1 _10638_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10147__B _10147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10862__S _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12643__A _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09785__B2 _07179_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09785__A1 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10569_ _10570_/A _10570_/B vssd1 vssd1 vccd1 vccd1 _10569_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_121_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13288_ _13289_/CLK _13288_/D vssd1 vssd1 vccd1 vccd1 hold292/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12308_ _12308_/A _12308_/B _12308_/C vssd1 vssd1 vccd1 vccd1 _12311_/A sky130_fd_sc_hd__or3_1
XFILLER_0_11_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11592__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11592__A1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12239_ hold165/A _12332_/B _12288_/B _12290_/C1 vssd1 vssd1 vccd1 vccd1 _12239_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10163__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07780_ _07780_/A _07780_/B vssd1 vssd1 vccd1 vccd1 _07781_/B sky130_fd_sc_hd__xnor2_4
X_06800_ _06866_/D _06798_/Y _06799_/X vssd1 vssd1 vccd1 vccd1 _06801_/B sky130_fd_sc_hd__a21oi_1
X_06731_ _07324_/A vssd1 vssd1 vccd1 vccd1 _07325_/A sky130_fd_sc_hd__inv_2
XANTENNA__08512__A2 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09450_ _09450_/A _09450_/B vssd1 vssd1 vccd1 vccd1 _09453_/B sky130_fd_sc_hd__xor2_1
X_06662_ instruction[29] _06678_/B vssd1 vssd1 vccd1 vccd1 _12578_/B sky130_fd_sc_hd__and2_4
X_08401_ _08401_/A _08401_/B vssd1 vssd1 vccd1 vccd1 _08430_/B sky130_fd_sc_hd__or2_1
X_06593_ instruction[35] _06633_/B vssd1 vssd1 vccd1 vccd1 _12607_/B sky130_fd_sc_hd__and2_4
X_09381_ _11823_/S _12726_/A _09382_/C vssd1 vssd1 vccd1 vccd1 _09381_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_59_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08276__B2 _08692_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08332_ _08371_/A _08371_/B vssd1 vssd1 vccd1 vccd1 _08372_/A sky130_fd_sc_hd__or2_1
XANTENNA__08276__A1 _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08263_ _08263_/A _08263_/B vssd1 vssd1 vccd1 vccd1 _08296_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07214_ _12774_/A _09618_/A1 fanout58/X _09618_/B2 vssd1 vssd1 vccd1 vccd1 _07215_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08194_ _08190_/A _08190_/B _08193_/Y vssd1 vssd1 vccd1 vccd1 _08242_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_6_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07145_ _09621_/A _07148_/B vssd1 vssd1 vccd1 vccd1 _07149_/A sky130_fd_sc_hd__and2_1
XFILLER_0_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07076_ _07077_/B _07077_/C _07077_/A vssd1 vssd1 vccd1 vccd1 _07079_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__07647__A _08853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07251__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07978_ _07978_/A _08658_/A _07978_/C vssd1 vssd1 vccd1 vccd1 _07980_/B sky130_fd_sc_hd__and3_1
XANTENNA__08478__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06929_ _09200_/A _09200_/B _12322_/S _09202_/A vssd1 vssd1 vccd1 vccd1 _06929_/X
+ sky130_fd_sc_hd__or4_2
X_09717_ _09656_/A _09656_/B _09654_/X vssd1 vssd1 vccd1 vccd1 _09814_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_96_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07711__B1 _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout46_A fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ _09649_/A _09649_/B vssd1 vssd1 vccd1 vccd1 _09648_/Y sky130_fd_sc_hd__nand2_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ _12760_/A _09752_/B fanout14/X _11134_/B2 vssd1 vssd1 vccd1 vccd1 _09580_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08267__B2 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08267__A1 _07004_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12063__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12590_/A _12590_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[6] sky130_fd_sc_hd__xor2_4
X_11610_ _11610_/A _11610_/B vssd1 vssd1 vccd1 vccd1 _11612_/B sky130_fd_sc_hd__xor2_1
X_11541_ _11542_/A _11542_/B vssd1 vssd1 vccd1 vccd1 _11632_/A sky130_fd_sc_hd__or2_1
XFILLER_0_107_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13012__A1 _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11472_ _06865_/B _11471_/Y _12228_/B1 vssd1 vssd1 vccd1 vccd1 _11472_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13211_ _13306_/CLK _13211_/D vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
X_10423_ _12255_/A _10423_/B vssd1 vssd1 vccd1 vccd1 _10432_/A sky130_fd_sc_hd__xnor2_1
X_13142_ hold286/X _13165_/A2 _13141_/X _13146_/B2 vssd1 vssd1 vccd1 vccd1 _13143_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10354_ _10356_/A _10356_/B vssd1 vssd1 vccd1 vccd1 _10354_/X sky130_fd_sc_hd__and2_1
XANTENNA__07557__A _09294_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13073_ _13073_/A _13073_/B vssd1 vssd1 vccd1 vccd1 _13073_/Y sky130_fd_sc_hd__xnor2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10285_ _10185_/A _10185_/B _10181_/Y vssd1 vssd1 vccd1 vccd1 _10297_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__09772__A _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12024_ _12025_/A _12025_/B _12025_/C vssd1 vssd1 vccd1 vccd1 _12026_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07950__B1 _10551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12926_ _13169_/A _12926_/B vssd1 vssd1 vccd1 vccd1 _13233_/D sky130_fd_sc_hd__and2_1
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12857_ hold65/X hold282/X vssd1 vssd1 vccd1 vccd1 _13092_/B sky130_fd_sc_hd__nand2b_1
X_11808_ _11808_/A vssd1 vssd1 vccd1 vccd1 _11810_/A sky130_fd_sc_hd__inv_2
XFILLER_0_29_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12788_ hold75/X _12788_/B vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__or2_1
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11739_ _11739_/A _11739_/B vssd1 vssd1 vccd1 vccd1 _11739_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07467__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08950_ _08950_/A _08950_/B vssd1 vssd1 vccd1 vccd1 _08953_/A sky130_fd_sc_hd__or2_1
XFILLER_0_20_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07901_ _08477_/B _08672_/B _10433_/A _08776_/B1 vssd1 vssd1 vccd1 vccd1 _07902_/B
+ sky130_fd_sc_hd__o22a_1
X_08881_ _08881_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _08883_/C sky130_fd_sc_hd__xnor2_2
X_07832_ _07833_/A _07833_/B vssd1 vssd1 vccd1 vccd1 _07832_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09930__A1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09930__B2 _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07763_ _07763_/A _07763_/B vssd1 vssd1 vccd1 vccd1 _07767_/A sky130_fd_sc_hd__xnor2_4
X_09502_ _09502_/A _09502_/B vssd1 vssd1 vccd1 vccd1 _09503_/B sky130_fd_sc_hd__xor2_4
X_06714_ reg1_val[12] _07303_/A vssd1 vssd1 vccd1 vccd1 _06715_/B sky130_fd_sc_hd__nand2_1
X_07694_ _07694_/A _07694_/B vssd1 vssd1 vccd1 vccd1 _07697_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06645_ _06645_/A vssd1 vssd1 vccd1 vccd1 _06647_/A sky130_fd_sc_hd__inv_2
X_09433_ _09596_/B _09433_/B vssd1 vssd1 vccd1 vccd1 _09436_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_93_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09364_ _09362_/X _09363_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09364_/X sky130_fd_sc_hd__mux2_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06576_ instruction[41] _06898_/B _06574_/X vssd1 vssd1 vccd1 vccd1 _06923_/A sky130_fd_sc_hd__a21o_1
X_08315_ _09478_/B2 _08420_/B _08854_/B2 _12730_/A vssd1 vssd1 vccd1 vccd1 _08316_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06546__A _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_20 reg1_val[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_31 reg1_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09295_ _09295_/A _09295_/B vssd1 vssd1 vccd1 vccd1 _09296_/C sky130_fd_sc_hd__or2_1
X_08246_ _08246_/A _08246_/B vssd1 vssd1 vccd1 vccd1 _08297_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_53 reg2_val[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_42 reg2_val[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_64 reg2_val[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_75 reg1_val[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08177_ _09180_/A _07179_/A _11012_/A _08544_/C vssd1 vssd1 vccd1 vccd1 _08178_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06680__B1 _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_86 _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07128_ _07153_/A _07128_/B _07128_/C _07128_/D vssd1 vssd1 vccd1 vccd1 _07128_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_113_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07059_ _07068_/A _07135_/B vssd1 vssd1 vccd1 vccd1 _07059_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07096__B _07097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11308__B2 _12228_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10070_ _10071_/A _10071_/B vssd1 vssd1 vccd1 vccd1 _10187_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_11_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10972_ _10972_/A _10972_/B vssd1 vssd1 vccd1 vccd1 _10972_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_69_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12711_ _12711_/A _12711_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[30] sky130_fd_sc_hd__xnor2_4
XFILLER_0_97_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap99 _07168_/Y vssd1 vssd1 vccd1 vccd1 _11222_/A sky130_fd_sc_hd__buf_6
X_12642_ reg1_val[15] _12637_/B _12640_/A vssd1 vssd1 vccd1 vccd1 _12644_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_38_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12573_ reg1_val[3] _12573_/B vssd1 vssd1 vccd1 vccd1 _12574_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08671__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11524_ _12022_/A _11524_/B vssd1 vssd1 vccd1 vccd1 _11525_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06671__B1 _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11455_ _11455_/A _11455_/B vssd1 vssd1 vccd1 vccd1 _11457_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07287__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ _12772_/A _10557_/B fanout13/X _11794_/A vssd1 vssd1 vccd1 vccd1 _10407_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11386_ _11294_/A _11291_/Y _11293_/B vssd1 vssd1 vccd1 vccd1 _11390_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13125_ _13147_/A hold253/X vssd1 vssd1 vccd1 vccd1 _13302_/D sky130_fd_sc_hd__and2_1
X_10337_ _10337_/A _10337_/B vssd1 vssd1 vccd1 vccd1 _10340_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _13066_/A _13056_/B vssd1 vssd1 vccd1 vccd1 _13288_/D sky130_fd_sc_hd__and2_1
X_10268_ _12373_/A1 _10245_/X _10251_/X _09837_/A _10267_/Y vssd1 vssd1 vccd1 vccd1
+ _10269_/D sky130_fd_sc_hd__a221o_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12007_ _12072_/A _11973_/B _11973_/A vssd1 vssd1 vccd1 vccd1 _12007_/X sky130_fd_sc_hd__a21o_1
X_10199_ _10200_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10201_/A sky130_fd_sc_hd__and2_1
XFILLER_0_17_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12909_ _13224_/Q _12947_/A2 _12947_/B1 hold187/X vssd1 vssd1 vccd1 vccd1 hold188/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12087__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08100_ _08154_/A _08154_/B vssd1 vssd1 vccd1 vccd1 _08155_/A sky130_fd_sc_hd__or2_1
XANTENNA__08651__A1 _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09080_ _09077_/A _08933_/B _08937_/Y vssd1 vssd1 vccd1 vccd1 _09082_/B sky130_fd_sc_hd__o21a_2
XANTENNA__08581__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08031_ _08033_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08031_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08651__B2 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06651__A2_N _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07197__A _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07206__A2 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09982_ hold288/A _10122_/C vssd1 vssd1 vccd1 vccd1 _09982_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08933_ _09077_/A _08933_/B _09098_/A _09103_/A vssd1 vssd1 vccd1 vccd1 _09090_/A
+ sky130_fd_sc_hd__or4_2
XFILLER_0_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12550__B _12551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout298_A _11647_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08864_ _08864_/A _08864_/B _08864_/C vssd1 vssd1 vccd1 vccd1 _08865_/B sky130_fd_sc_hd__and3_1
XANTENNA__10513__A2 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ _08733_/A _07815_/B vssd1 vssd1 vccd1 vccd1 _07842_/A sky130_fd_sc_hd__xor2_4
X_08795_ _08796_/B _08796_/A vssd1 vssd1 vccd1 vccd1 _08795_/Y sky130_fd_sc_hd__nand2b_1
X_07746_ _08775_/A _07746_/B vssd1 vssd1 vccd1 vccd1 _07747_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10277__A1 _07277_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__B2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10497__S _11647_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07677_ _08831_/A _07675_/Y _07672_/Y vssd1 vssd1 vccd1 vccd1 _07678_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12278__A _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09416_ _09416_/A _09416_/B vssd1 vssd1 vccd1 vccd1 _09418_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06628_ _06626_/Y _06680_/B1 _06778_/B reg2_val[30] vssd1 vssd1 vccd1 vccd1 _07434_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_06559_ instruction[18] _06915_/B vssd1 vssd1 vccd1 vccd1 _06559_/X sky130_fd_sc_hd__or2_1
X_09347_ _09343_/X _09346_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09347_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_118_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ _09621_/A _09279_/B vssd1 vssd1 vccd1 vccd1 _09278_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08229_ _08227_/Y _08284_/B _08224_/Y vssd1 vssd1 vccd1 vccd1 _08240_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11240_ _11604_/A _11240_/B vssd1 vssd1 vccd1 vccd1 _11328_/B sky130_fd_sc_hd__xnor2_2
X_11171_ _11171_/A _11171_/B _11171_/C vssd1 vssd1 vccd1 vccd1 _11172_/B sky130_fd_sc_hd__nand3_1
X_10122_ hold284/A hold288/A _10122_/C vssd1 vssd1 vccd1 vccd1 _10256_/B sky130_fd_sc_hd__or3_1
XFILLER_0_101_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10053_ _10156_/A1 fanout20/X fanout18/X _10156_/B2 vssd1 vssd1 vccd1 vccd1 _10054_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_89_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08666__A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10268__A1 _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11465__B1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10955_ _10843_/A _10841_/X _10840_/X vssd1 vssd1 vccd1 vccd1 _10958_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_128_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10886_ _10857_/Y _10860_/Y _10864_/X _10885_/X _12345_/A vssd1 vssd1 vccd1 vccd1
+ _10886_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12625_ reg1_val[13] _12626_/B vssd1 vssd1 vccd1 vccd1 _12635_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_503 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12556_ reg1_val[27] curr_PC[27] _12556_/S vssd1 vssd1 vccd1 vccd1 _12557_/B sky130_fd_sc_hd__mux2_2
XANTENNA_max_cap10_A _07435_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11507_ _12200_/A _11507_/B vssd1 vssd1 vccd1 vccd1 _11509_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06633__B _06633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12487_ reg1_val[16] curr_PC[16] _12487_/S vssd1 vssd1 vccd1 vccd1 _12488_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10991__A2 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09189__A2 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11438_ _11438_/A _11438_/B vssd1 vssd1 vccd1 vccd1 _11439_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_111_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12193__A1 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11369_ _11369_/A _11369_/B _11369_/C vssd1 vssd1 vccd1 vccd1 _11370_/B sky130_fd_sc_hd__nand3_1
X_13108_ _13108_/A _13108_/B vssd1 vssd1 vccd1 vccd1 _13108_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11940__B2 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11940__A1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12370__B _12370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13039_ _13039_/A _13039_/B vssd1 vssd1 vccd1 vccd1 _13039_/Y sky130_fd_sc_hd__xnor2_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08580_ _08825_/A2 _08588_/B _09273_/A1 _08588_/A vssd1 vssd1 vccd1 vccd1 _08581_/B
+ sky130_fd_sc_hd__o22a_1
X_07600_ _07601_/A _07601_/B _07601_/C vssd1 vssd1 vccd1 vccd1 _07600_/X sky130_fd_sc_hd__o21a_1
X_07531_ _09362_/S _10551_/B vssd1 vssd1 vccd1 vccd1 _07539_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07462_ _07462_/A _07462_/B vssd1 vssd1 vccd1 vccd1 _07463_/A sky130_fd_sc_hd__xnor2_1
X_09201_ instruction[5] _09201_/B _09200_/A vssd1 vssd1 vccd1 vccd1 _09201_/X sky130_fd_sc_hd__or3b_4
X_07393_ _08595_/A _07393_/B _07393_/C vssd1 vssd1 vccd1 vccd1 _07396_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_17_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09132_ reg1_val[9] reg1_val[22] _09172_/S vssd1 vssd1 vccd1 vccd1 _09132_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12545__B _12545_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09063_ _09063_/A _09063_/B vssd1 vssd1 vccd1 vccd1 _11379_/C sky130_fd_sc_hd__xnor2_4
XANTENNA__06635__B1 _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08014_ _08014_/A _08014_/B vssd1 vssd1 vccd1 vccd1 _08016_/B sky130_fd_sc_hd__or2_2
XFILLER_0_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08388__B1 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11931__A1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10195__B1 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09965_ _10617_/A _09966_/B _09966_/C vssd1 vssd1 vccd1 vccd1 _09965_/Y sky130_fd_sc_hd__o21ai_1
X_08916_ _08916_/A _08916_/B vssd1 vssd1 vccd1 vccd1 _08929_/A sky130_fd_sc_hd__nor2_2
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09896_ _10458_/A _09896_/B vssd1 vssd1 vccd1 vccd1 _09898_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09888__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08847_ _08847_/A _08847_/B vssd1 vssd1 vccd1 vccd1 _08848_/B sky130_fd_sc_hd__xnor2_2
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07363__B2 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07363__A1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08560__B1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08778_ _08779_/A _08779_/B vssd1 vssd1 vccd1 vccd1 _08778_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07729_ _07173_/Y _10551_/A _07325_/Y _07182_/X vssd1 vssd1 vccd1 vccd1 _07730_/B
+ sky130_fd_sc_hd__a22o_1
X_10740_ _12131_/A _10740_/B _10740_/C vssd1 vssd1 vccd1 vccd1 _10740_/X sky130_fd_sc_hd__or3_1
XFILLER_0_48_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10671_ fanout29/X _11431_/A fanout70/X fanout32/X vssd1 vssd1 vccd1 vccd1 _10672_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12736__A _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12410_ reg1_val[5] curr_PC[5] _12524_/S vssd1 vssd1 vccd1 vccd1 _12412_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_106_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12341_ _09198_/X _12331_/X _12332_/Y _12336_/X _12340_/Y vssd1 vssd1 vccd1 vccd1
+ _12341_/X sky130_fd_sc_hd__a311o_1
XANTENNA__10422__B2 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10422__A1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12272_ _12317_/B _12272_/B vssd1 vssd1 vccd1 vccd1 _12272_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_120_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11223_ _11222_/A _12200_/A _11222_/C vssd1 vssd1 vccd1 vccd1 _11224_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09764__B fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07565__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11154_ _11052_/A _11052_/B _11055_/A vssd1 vssd1 vccd1 vccd1 _11162_/A sky130_fd_sc_hd__a21bo_1
X_11085_ reg1_val[14] curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11086_/B sky130_fd_sc_hd__or2_1
X_10105_ _11184_/A _10105_/B _10104_/X vssd1 vssd1 vccd1 vccd1 _10105_/X sky130_fd_sc_hd__or3b_1
X_10036_ _10037_/A _10037_/B _10037_/C vssd1 vssd1 vccd1 vccd1 _10206_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11987_ _11987_/A _11987_/B vssd1 vssd1 vccd1 vccd1 _11987_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08854__A1 _07031_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10938_ _10938_/A _10938_/B vssd1 vssd1 vccd1 vccd1 _10951_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08854__B2 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10869_ reg1_val[12] curr_PC[12] vssd1 vssd1 vccd1 vccd1 _10869_/X sky130_fd_sc_hd__or2_1
XFILLER_0_73_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12608_ _12617_/A _12608_/B vssd1 vssd1 vccd1 vccd1 _12611_/B sky130_fd_sc_hd__nand2_1
X_12539_ _12539_/A _12539_/B _12539_/C _12539_/D vssd1 vssd1 vccd1 vccd1 _12541_/C
+ sky130_fd_sc_hd__or4_1
XANTENNA__08082__A2 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10177__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07194__B _10819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06962_ _07279_/A _09392_/S _09362_/S _12370_/B _09968_/A vssd1 vssd1 vccd1 vccd1
+ _06964_/B sky130_fd_sc_hd__o311a_2
X_09750_ fanout77/X fanout95/X fanout54/X fanout75/X vssd1 vssd1 vccd1 vccd1 _09751_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08701_ _08701_/A _08701_/B _08701_/C vssd1 vssd1 vccd1 vccd1 _08703_/B sky130_fd_sc_hd__or3_1
X_09681_ _09677_/X _09680_/X _11089_/A vssd1 vssd1 vccd1 vccd1 _09681_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11677__B1 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06893_ hold163/A _12721_/B vssd1 vssd1 vccd1 vccd1 busy sky130_fd_sc_hd__nor2_8
X_08632_ _08633_/A _08633_/B vssd1 vssd1 vccd1 vccd1 _09072_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07345__B2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07345__A1 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08563_ _09620_/A _08563_/B vssd1 vssd1 vccd1 vccd1 _08570_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08494_ _06864_/A _08841_/B2 _08837_/B2 _08758_/A2 vssd1 vssd1 vccd1 vccd1 _08495_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10101__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07514_ _10184_/A _07514_/B vssd1 vssd1 vccd1 vccd1 _07516_/B sky130_fd_sc_hd__xnor2_1
Xfanout15 _07278_/B vssd1 vssd1 vccd1 vccd1 fanout15/X sky130_fd_sc_hd__clkbuf_8
Xfanout26 _07099_/X vssd1 vssd1 vccd1 vccd1 fanout26/X sky130_fd_sc_hd__buf_8
Xfanout37 _08821_/B vssd1 vssd1 vccd1 vccd1 fanout37/X sky130_fd_sc_hd__buf_6
X_07445_ _10180_/A _07445_/B vssd1 vssd1 vccd1 vccd1 _07447_/B sky130_fd_sc_hd__xnor2_1
Xfanout59 _07157_/Y vssd1 vssd1 vccd1 vccd1 _12776_/A sky130_fd_sc_hd__buf_6
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout48 _09752_/B vssd1 vssd1 vccd1 vccd1 _10557_/B sky130_fd_sc_hd__buf_6
XFILLER_0_91_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07376_ _07376_/A _07376_/B vssd1 vssd1 vccd1 vccd1 _07692_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09115_ _11738_/S _09184_/B vssd1 vssd1 vccd1 vccd1 _09115_/X sky130_fd_sc_hd__or2_4
XANTENNA__06608__B1 _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11601__B1 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09046_ _09046_/A _09046_/B vssd1 vssd1 vccd1 vccd1 _10370_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_4_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09865__A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10804__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10168__B1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09948_ _09948_/A _09948_/B vssd1 vssd1 vccd1 vccd1 _09950_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08533__B1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07336__B2 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07336__A1 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _09879_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _09879_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11132__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12890_ _12891_/B _12891_/C hold75/X vssd1 vssd1 vccd1 vccd1 _13167_/B sky130_fd_sc_hd__a21oi_1
X_11910_ _11910_/A _11910_/B vssd1 vssd1 vccd1 vccd1 _11912_/A sky130_fd_sc_hd__nor2_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _09115_/X _10507_/Y _10518_/Y _09184_/X _11840_/X vssd1 vssd1 vccd1 vccd1
+ _11841_/X sky130_fd_sc_hd__o221a_1
XANTENNA__10891__A1 _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10891__B2 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ _12022_/A _11772_/B vssd1 vssd1 vccd1 vccd1 _11773_/B sky130_fd_sc_hd__xnor2_1
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10723_ _10724_/A _10724_/B vssd1 vssd1 vccd1 vccd1 _10723_/X sky130_fd_sc_hd__and2_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_125_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10654_ fanout56/X fanout18/X fanout9/X fanout98/X vssd1 vssd1 vccd1 vccd1 _10655_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10585_ _10586_/A _10586_/B _10586_/C vssd1 vssd1 vccd1 vccd1 _10587_/A sky130_fd_sc_hd__a21oi_1
X_12324_ _06856_/A _12322_/X _12323_/Y vssd1 vssd1 vccd1 vccd1 _12324_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09775__A _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06911__B _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12255_ _12255_/A _12255_/B vssd1 vssd1 vccd1 vccd1 _12255_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_121_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11206_ _11187_/A _09383_/B _11202_/Y _11203_/X _11205_/X vssd1 vssd1 vccd1 vccd1
+ _11206_/X sky130_fd_sc_hd__o221a_1
X_12186_ hold183/A _12186_/B vssd1 vssd1 vccd1 vccd1 _12237_/B sky130_fd_sc_hd__or2_1
XANTENNA__09564__A2 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08772__B1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11137_ _12022_/A _11137_/B vssd1 vssd1 vccd1 vccd1 _11139_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10433__B _12349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11068_ _11068_/A _11068_/B vssd1 vssd1 vccd1 vccd1 _11462_/A sky130_fd_sc_hd__or2_2
XANTENNA__09660__D _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10019_ _10019_/A _10019_/B vssd1 vssd1 vccd1 vccd1 _10020_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_59_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07230_ _10452_/B2 _10553_/B fanout69/X _10527_/A vssd1 vssd1 vccd1 vccd1 _07231_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07161_ _07411_/A _07411_/B vssd1 vssd1 vccd1 vccd1 _07383_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07263__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07092_ _09679_/S _07093_/B vssd1 vssd1 vccd1 vccd1 _09283_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_41_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09004__A1 _08018_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 _08311_/A vssd1 vssd1 vccd1 vccd1 _08443_/A sky130_fd_sc_hd__buf_12
XFILLER_0_10_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout238 _09201_/X vssd1 vssd1 vccd1 vccd1 _11400_/A sky130_fd_sc_hd__buf_4
Xfanout227 _07001_/C vssd1 vssd1 vccd1 vccd1 _11195_/A sky130_fd_sc_hd__clkbuf_4
Xfanout216 _06784_/Y vssd1 vssd1 vccd1 vccd1 _12726_/A sky130_fd_sc_hd__buf_4
X_09802_ _09803_/A _09803_/B vssd1 vssd1 vccd1 vccd1 _09802_/Y sky130_fd_sc_hd__nor2_1
X_07994_ _07994_/A _07994_/B vssd1 vssd1 vccd1 vccd1 _07995_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_66_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout249 _08695_/A vssd1 vssd1 vccd1 vccd1 _09621_/A sky130_fd_sc_hd__buf_12
XANTENNA__09307__A2 _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout280_A _06569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06945_ reg1_val[27] _06945_/B vssd1 vssd1 vccd1 vccd1 _12143_/A sky130_fd_sc_hd__xnor2_4
X_09733_ _09733_/A _09733_/B vssd1 vssd1 vccd1 vccd1 _09797_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_69_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06876_ _09201_/B vssd1 vssd1 vccd1 vccd1 _09200_/C sky130_fd_sc_hd__inv_2
X_09664_ _10229_/A _09664_/B vssd1 vssd1 vccd1 vccd1 _10273_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_96_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08615_ _08611_/X _08613_/X _08486_/Y vssd1 vssd1 vccd1 vccd1 _09055_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_49_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09595_ _09596_/A _09596_/B _09596_/C _09596_/D vssd1 vssd1 vccd1 vccd1 _09597_/B
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_77_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08546_ _08595_/A _08546_/B _08546_/C vssd1 vssd1 vccd1 vccd1 _08549_/B sky130_fd_sc_hd__and3_1
XFILLER_0_65_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08477_ _08588_/A _08477_/B vssd1 vssd1 vccd1 vccd1 _08478_/B sky130_fd_sc_hd__nor2_1
X_07428_ _07426_/A _07426_/B _07427_/Y vssd1 vssd1 vccd1 vccd1 _07620_/A sky130_fd_sc_hd__o21ai_4
X_07359_ fanout36/X _08825_/A2 _09476_/A _08821_/B vssd1 vssd1 vccd1 vccd1 _07360_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10370_ _11973_/A _10370_/B _10370_/C vssd1 vssd1 vccd1 vccd1 _10370_/X sky130_fd_sc_hd__or3_1
XFILLER_0_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09029_ _08806_/X _09029_/B _09076_/A vssd1 vssd1 vccd1 vccd1 _09029_/Y sky130_fd_sc_hd__nand3b_1
Xhold270 hold270/A vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__dlygate4sd3_1
X_12040_ _12163_/A _12040_/B vssd1 vssd1 vccd1 vccd1 _12072_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold281 hold281/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 hold292/A vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08004__A _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_12_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12302__A1 _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12942_ _13169_/A hold227/X vssd1 vssd1 vccd1 vccd1 _13241_/D sky130_fd_sc_hd__and2_1
XANTENNA__06780__A2 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12873_ _13126_/A _12872_/B _12802_/X vssd1 vssd1 vccd1 vccd1 _13131_/A sky130_fd_sc_hd__a21o_1
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08674__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11824_ _11824_/A _11824_/B vssd1 vssd1 vccd1 vccd1 _11824_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_68_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11755_ _11756_/A _09383_/B _09191_/X vssd1 vssd1 vccd1 vccd1 _11755_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10706_ _10706_/A _10706_/B vssd1 vssd1 vccd1 vccd1 _10707_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_126_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11686_ _11686_/A _11686_/B vssd1 vssd1 vccd1 vccd1 _11687_/B sky130_fd_sc_hd__or2_1
X_10637_ hold301/A _09842_/B _10758_/B _10636_/Y _12339_/B1 vssd1 vssd1 vccd1 vccd1
+ _10641_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_11_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10568_ _10705_/C _10568_/B vssd1 vssd1 vccd1 vccd1 _10570_/B sky130_fd_sc_hd__nor2_2
XANTENNA__09785__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13287_ _13310_/CLK _13287_/D vssd1 vssd1 vccd1 vccd1 hold266/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10499_ _10498_/A _10498_/B _10498_/Y _12277_/B1 vssd1 vssd1 vccd1 vccd1 _10499_/X
+ sky130_fd_sc_hd__a211o_1
X_12307_ _12307_/A _12307_/B vssd1 vssd1 vccd1 vccd1 _12308_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10444__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11592__A2 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12238_ _12332_/B _12288_/B hold165/A vssd1 vssd1 vccd1 vccd1 _12238_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06641__B _12593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08745__B1 _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12169_ _06620_/B _12108_/X _06619_/A vssd1 vssd1 vccd1 vccd1 _12169_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06730_ _06783_/A _06641_/A _12607_/B _06729_/X vssd1 vssd1 vccd1 vccd1 _07324_/A
+ sky130_fd_sc_hd__a31o_4
X_06661_ _11906_/A _11824_/A _06661_/C _11739_/A vssd1 vssd1 vccd1 vccd1 _06872_/B
+ sky130_fd_sc_hd__nor4_1
X_08400_ _08407_/A _08407_/B vssd1 vssd1 vccd1 vccd1 _08401_/B sky130_fd_sc_hd__and2b_1
X_09380_ _09383_/A _09380_/B vssd1 vssd1 vccd1 vccd1 _09382_/C sky130_fd_sc_hd__xnor2_1
X_06592_ _06605_/B vssd1 vssd1 vccd1 vccd1 _06592_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_47_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08276__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08331_ _08331_/A _08331_/B vssd1 vssd1 vccd1 vccd1 _08371_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08262_ _08263_/A _08263_/B vssd1 vssd1 vccd1 vccd1 _08295_/A sky130_fd_sc_hd__or2_1
XFILLER_0_116_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07213_ _07222_/A vssd1 vssd1 vccd1 vccd1 _07213_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08193_ _08247_/B _08247_/A vssd1 vssd1 vccd1 vccd1 _08193_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout126_A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07144_ reg1_val[2] _07144_/B vssd1 vssd1 vccd1 vccd1 _07148_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_15_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07075_ _07075_/A _07075_/B vssd1 vssd1 vccd1 vccd1 _07077_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08736__B1 _08672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08759__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ _07977_/A _07977_/B _07977_/C vssd1 vssd1 vccd1 vccd1 _07978_/C sky130_fd_sc_hd__nand3_1
X_06928_ _09198_/C instruction[5] _09968_/A _06928_/D vssd1 vssd1 vccd1 vccd1 _06928_/X
+ sky130_fd_sc_hd__and4b_4
X_09716_ _10617_/A _10002_/A vssd1 vssd1 vccd1 vccd1 _09716_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06859_ _12713_/A _12370_/B _06858_/X vssd1 vssd1 vccd1 vccd1 _06859_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09647_ _09485_/A _09485_/B _09483_/X vssd1 vssd1 vccd1 vccd1 _09649_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12048__B1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11913__A _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09578_ _09416_/A _09416_/B _09413_/A vssd1 vssd1 vccd1 vccd1 _09593_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__08267__A2 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08529_ _08529_/A _08529_/B vssd1 vssd1 vccd1 vccd1 _08531_/B sky130_fd_sc_hd__nor2_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout39_A _12349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ _11540_/A _11540_/B vssd1 vssd1 vccd1 vccd1 _11542_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13012__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11471_ _11738_/S _06820_/Y _11470_/Y vssd1 vssd1 vccd1 vccd1 _11471_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13210_ _13305_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_751 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10422_ fanout27/X _10927_/A fanout83/X _12205_/A vssd1 vssd1 vccd1 vccd1 _10423_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12771__A1 _11793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13141_ hold262/X _13140_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13141_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07557__B _10551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10353_ _10353_/A _10353_/B vssd1 vssd1 vccd1 vccd1 _10356_/B sky130_fd_sc_hd__xnor2_1
X_13072_ _13072_/A _13072_/B vssd1 vssd1 vccd1 vccd1 _13073_/B sky130_fd_sc_hd__nand2_1
X_10284_ _10284_/A _10284_/B vssd1 vssd1 vccd1 vccd1 _10312_/A sky130_fd_sc_hd__xnor2_1
X_12023_ _12023_/A _12023_/B vssd1 vssd1 vccd1 vccd1 _12025_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__08669__A _08853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09772__B _12349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10534__B1 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07950__A1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07950__B2 _07182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06753__A2 _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12925_ hold203/X _12955_/A2 _13168_/B1 hold207/X vssd1 vssd1 vccd1 vccd1 _12926_/B
+ sky130_fd_sc_hd__a22o_1
X_12856_ _13087_/A _13088_/A _13087_/B vssd1 vssd1 vccd1 vccd1 _13093_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11934__A2_N fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _11809_/A _11809_/B _11809_/C vssd1 vssd1 vccd1 vccd1 _11808_/A sky130_fd_sc_hd__a21o_1
X_12787_ hold3/X _12786_/B _12786_/Y _13166_/A vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__o211a_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07466__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11738_ _11736_/X _11737_/X _11738_/S vssd1 vssd1 vccd1 vccd1 _11739_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11669_ _11644_/Y _11645_/X _11668_/X _11643_/X vssd1 vssd1 vccd1 vccd1 _11669_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07218__B1 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07900_ _08773_/A _07900_/B vssd1 vssd1 vccd1 vccd1 _08030_/A sky130_fd_sc_hd__xnor2_2
X_08880_ _08880_/A _08880_/B vssd1 vssd1 vccd1 vccd1 _08881_/B sky130_fd_sc_hd__xor2_2
XANTENNA__08579__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10902__A _11780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07831_ _07831_/A _07831_/B vssd1 vssd1 vccd1 vccd1 _07833_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_47_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09930__A2 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07762_ _07023_/Y _08774_/A2 _08774_/B1 _12760_/A vssd1 vssd1 vccd1 vccd1 _07763_/B
+ sky130_fd_sc_hd__o22a_2
X_09501_ _09502_/A _09502_/B vssd1 vssd1 vccd1 vccd1 _09501_/X sky130_fd_sc_hd__and2_1
X_06713_ reg1_val[12] _07303_/A vssd1 vssd1 vccd1 vccd1 _06713_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07693_ _07693_/A _07693_/B vssd1 vssd1 vccd1 vccd1 _07697_/A sky130_fd_sc_hd__or2_1
XFILLER_0_2_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06644_ reg1_val[22] _07112_/B vssd1 vssd1 vccd1 vccd1 _06645_/A sky130_fd_sc_hd__nand2_1
X_09432_ _09432_/A _09432_/B vssd1 vssd1 vccd1 vccd1 _09433_/B sky130_fd_sc_hd__nor2_1
X_06575_ instruction[1] instruction[2] instruction[25] pred_val vssd1 vssd1 vccd1
+ vccd1 _06575_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_93_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09363_ _09166_/X _09169_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09363_/X sky130_fd_sc_hd__mux2_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08314_ _08362_/A _08313_/B _08309_/X vssd1 vssd1 vccd1 vccd1 _08320_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_74_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10056__A2 _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_21 reg1_val[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09294_ _09294_/A _10694_/A vssd1 vssd1 vccd1 vccd1 _09296_/B sky130_fd_sc_hd__nand2_1
XANTENNA_32 reg1_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 reg1_val[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08245_ _08245_/A _08245_/B vssd1 vssd1 vccd1 vccd1 _08246_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_43 reg2_val[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_65 reg2_val[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_54 reg2_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08176_ _08775_/A _08176_/B vssd1 vssd1 vccd1 vccd1 _08183_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_76 reg1_val[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07127_ _07128_/B _07128_/C _07128_/D vssd1 vssd1 vccd1 vccd1 _07127_/X sky130_fd_sc_hd__and3_1
XFILLER_0_15_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07058_ _07058_/A vssd1 vssd1 vccd1 vccd1 _09253_/A sky130_fd_sc_hd__inv_2
XFILLER_0_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06983__A2 _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07393__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10971_ _06810_/X _10970_/X _11738_/S vssd1 vssd1 vccd1 vccd1 _10972_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_97_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11492__A1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12710_ _12704_/A _12706_/B _12704_/B vssd1 vssd1 vccd1 vccd1 _12711_/B sky130_fd_sc_hd__a21bo_2
XFILLER_0_84_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ _12641_/A _12658_/A vssd1 vssd1 vccd1 vccd1 _12644_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12572_ reg1_val[3] _12573_/B vssd1 vssd1 vccd1 vccd1 _12572_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_108_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12474__A _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12992__A1 _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11523_ fanout35/X _11935_/A _12776_/A fanout37/X vssd1 vssd1 vccd1 vccd1 _11524_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_18_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11454_ _11455_/A _11455_/B vssd1 vssd1 vccd1 vccd1 _11547_/B sky130_fd_sc_hd__and2_1
XFILLER_0_123_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _10351_/A _10351_/B _10352_/Y vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__o21ai_4
X_11385_ _06865_/C _11383_/X _11384_/Y vssd1 vssd1 vccd1 vccd1 _11404_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13124_ hold252/X _13165_/A2 _13123_/X _13146_/B2 vssd1 vssd1 vccd1 vccd1 hold253/A
+ sky130_fd_sc_hd__a22o_1
X_10336_ _11499_/A _10336_/B vssd1 vssd1 vccd1 vccd1 _10337_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ hold292/X _12721_/B _13054_/X _12722_/A vssd1 vssd1 vccd1 vccd1 _13056_/B
+ sky130_fd_sc_hd__a22o_1
X_10267_ _11197_/S _09205_/B _10266_/Y _10261_/X vssd1 vssd1 vccd1 vccd1 _10267_/Y
+ sky130_fd_sc_hd__o31ai_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12006_ _12005_/A _12002_/X _12003_/X _12005_/Y vssd1 vssd1 vccd1 vccd1 dest_val[24]
+ sky130_fd_sc_hd__a22o_4
X_10198_ _10559_/A _10198_/B vssd1 vssd1 vccd1 vccd1 _10200_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11180__B1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12908_ _12946_/A hold229/X vssd1 vssd1 vccd1 vccd1 hold230/A sky130_fd_sc_hd__and2_1
XFILLER_0_69_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12839_ hold77/X hold284/X vssd1 vssd1 vccd1 vccd1 _13047_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_33_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10169__A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08651__A2 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12384__A _12563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08030_ _08030_/A _08030_/B vssd1 vssd1 vccd1 vccd1 _08033_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_114_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_4_5_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13303_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09981_ hold189/A _09980_/B _09198_/X vssd1 vssd1 vccd1 vccd1 _09981_/X sky130_fd_sc_hd__o21a_1
X_08932_ _08932_/A _08932_/B vssd1 vssd1 vccd1 vccd1 _09103_/A sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout193_A _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08863_ _08864_/A _08864_/B _08864_/C vssd1 vssd1 vccd1 vccd1 _08865_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07814_ _10281_/A _07173_/Y _07182_/X _10149_/A vssd1 vssd1 vccd1 vccd1 _07815_/B
+ sky130_fd_sc_hd__a22o_2
X_08794_ _08794_/A _08794_/B vssd1 vssd1 vccd1 vccd1 _08796_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09116__A0 _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07745_ _12760_/A _08774_/A2 _08774_/B1 _09925_/A1 vssd1 vssd1 vccd1 vccd1 _07746_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13154__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__A2 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ _07676_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _08831_/B sky130_fd_sc_hd__xnor2_1
X_09415_ _10301_/A _09415_/B vssd1 vssd1 vccd1 vccd1 _09416_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06627_ reg2_val[30] _06778_/B _06680_/B1 _06626_/Y vssd1 vssd1 vccd1 vccd1 _06834_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_06558_ instruction[14] _06552_/X _06557_/X _06678_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[3]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09346_ _09344_/X _09345_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09346_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12974__A1 _07080_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09277_ _09467_/A _09277_/B vssd1 vssd1 vccd1 vccd1 _09279_/B sky130_fd_sc_hd__xnor2_4
X_08228_ _08228_/A _08228_/B vssd1 vssd1 vccd1 vccd1 _08284_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10985__B1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07850__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08159_ _08167_/B _08167_/A vssd1 vssd1 vccd1 vccd1 _08160_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_43_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10737__B1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11170_ _11171_/A _11171_/B _11171_/C vssd1 vssd1 vccd1 vccd1 _11170_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ hold228/A _12124_/B _10252_/B _12290_/C1 vssd1 vssd1 vccd1 vccd1 _10121_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09108__A _09559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10542__A _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10052_ _10052_/A _10052_/B vssd1 vssd1 vccd1 vccd1 _10061_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07851__A _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13064__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10954_ _11067_/B _10954_/B vssd1 vssd1 vccd1 vccd1 _10958_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10885_ _09184_/X _10867_/Y _10873_/X _09205_/B _10884_/X vssd1 vssd1 vccd1 vccd1
+ _10885_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_66_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12624_ _12629_/B _12624_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[12] sky130_fd_sc_hd__and2_4
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12555_ _12552_/B _12554_/B _12552_/A vssd1 vssd1 vccd1 vccd1 _12558_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_108_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11506_ _11704_/A fanout15/X fanout6/X _11688_/A vssd1 vssd1 vccd1 vccd1 _11507_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_110_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12486_ _12490_/B _12486_/B vssd1 vssd1 vccd1 vccd1 new_PC[15] sky130_fd_sc_hd__and2_4
XFILLER_0_110_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11437_ _11437_/A _11437_/B vssd1 vssd1 vccd1 vccd1 _11438_/B sky130_fd_sc_hd__or2_1
XFILLER_0_22_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11368_ _11369_/A _11369_/B _11369_/C vssd1 vssd1 vccd1 vccd1 _11368_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13107_ _12806_/X _13107_/B vssd1 vssd1 vccd1 vccd1 _13108_/B sky130_fd_sc_hd__nand2b_1
X_10319_ _10320_/A _10320_/B _10320_/C vssd1 vssd1 vccd1 vccd1 _10473_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11940__A2 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13142__B2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11299_ reg1_val[16] _11099_/B _07168_/A _06928_/X vssd1 vssd1 vccd1 vccd1 _11299_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13086_/A hold247/X vssd1 vssd1 vccd1 vccd1 _13284_/D sky130_fd_sc_hd__and2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08857__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10259__A2 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12379__A _12560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07530_ _09968_/A _07528_/X _12713_/A vssd1 vssd1 vccd1 vccd1 _07530_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07461_ _09452_/A _07461_/B vssd1 vssd1 vccd1 vccd1 _07462_/B sky130_fd_sc_hd__xnor2_1
X_09200_ _09200_/A _09200_/B _09200_/C vssd1 vssd1 vccd1 vccd1 _09200_/X sky130_fd_sc_hd__and3_2
X_07392_ _07393_/B _07393_/C _08595_/A vssd1 vssd1 vccd1 vccd1 _07396_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09131_ reg1_val[8] reg1_val[23] _09172_/S vssd1 vssd1 vccd1 vccd1 _09131_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09062_ _11183_/B _11183_/C _11285_/A vssd1 vssd1 vccd1 vccd1 _11379_/B sky130_fd_sc_hd__and3_1
XFILLER_0_72_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08013_ _08013_/A _08013_/B vssd1 vssd1 vccd1 vccd1 _08016_/A sky130_fd_sc_hd__xor2_4
XANTENNA_fanout206_A _07763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07001__A _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08388__B2 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08388__A1 _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09585__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07060__A1 _06653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10195__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10195__A1 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09964_ _09859_/X _10002_/C _09963_/Y vssd1 vssd1 vccd1 vccd1 _09964_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_0_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13133__B2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08915_ _08914_/B _08914_/C _08914_/A vssd1 vssd1 vccd1 vccd1 _08916_/B sky130_fd_sc_hd__a21oi_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09895_ _10156_/A1 _12782_/A fanout20/X _10156_/B2 vssd1 vssd1 vccd1 vccd1 _09896_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09888__A1 _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09888__B2 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08846_ _08847_/A _08847_/B vssd1 vssd1 vccd1 vccd1 _08846_/X sky130_fd_sc_hd__and2b_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07671__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09362__S _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07363__A2 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08560__A1 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08560__B2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08777_ _08777_/A _08777_/B vssd1 vssd1 vccd1 vccd1 _08779_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07728_ _07727_/A _07727_/B _07727_/C vssd1 vssd1 vccd1 vccd1 _07738_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11998__A2 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07659_ _10015_/A _07659_/B vssd1 vssd1 vccd1 vccd1 _07661_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout21_A _07138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10670_ _10670_/A _10670_/B vssd1 vssd1 vccd1 vccd1 _10674_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_125_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12736__B _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09329_ _09331_/A _09331_/B vssd1 vssd1 vccd1 vccd1 _09329_/X sky130_fd_sc_hd__or2_1
XFILLER_0_48_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10537__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07823__B1 _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12340_ _12338_/Y _12339_/X _12327_/X vssd1 vssd1 vccd1 vccd1 _12340_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__09110__B _09199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10422__A2 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12752__A _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10971__S _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12271_ _11973_/B _12317_/A _12221_/X _11973_/A vssd1 vssd1 vccd1 vccd1 _12272_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11907__C1 _12228_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11222_ _11222_/A _12200_/A _11222_/C vssd1 vssd1 vccd1 vccd1 _11224_/A sky130_fd_sc_hd__and3_1
XFILLER_0_120_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13059__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10989__A2_N _06928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ _11046_/A _11046_/B _11047_/X vssd1 vssd1 vccd1 vccd1 _11164_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__13124__B2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11084_ reg1_val[14] curr_PC[14] vssd1 vssd1 vccd1 vccd1 _11086_/A sky130_fd_sc_hd__nand2_1
X_10104_ _10617_/A _10104_/B _10104_/C vssd1 vssd1 vccd1 vccd1 _10104_/X sky130_fd_sc_hd__or3_1
X_10035_ _10035_/A _11147_/B vssd1 vssd1 vccd1 vccd1 _10037_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06909__B _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08303__A1 _10281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ _11984_/Y _11986_/B vssd1 vssd1 vccd1 vccd1 _11987_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08303__B2 _10149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08854__A2 _09925_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10937_ _10937_/A _10937_/B vssd1 vssd1 vccd1 vccd1 _10938_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06925__A _12487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10868_ reg1_val[12] curr_PC[12] vssd1 vssd1 vccd1 vccd1 _10868_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12607_ reg1_val[10] _12607_/B vssd1 vssd1 vccd1 vccd1 _12608_/B sky130_fd_sc_hd__or2_1
XFILLER_0_14_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10799_ _11853_/A _10799_/B vssd1 vssd1 vccd1 vccd1 _10801_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12538_ _12557_/A _12538_/B vssd1 vssd1 vccd1 vccd1 _12542_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07814__B1 _07182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12469_ _12478_/A _12469_/B vssd1 vssd1 vccd1 vccd1 _12471_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10177__B2 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10177__A1 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13115__B2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06961_ _09392_/S _09362_/S _11823_/S _12370_/B vssd1 vssd1 vccd1 vccd1 _07279_/B
+ sky130_fd_sc_hd__o211a_1
X_08700_ _08700_/A _08700_/B vssd1 vssd1 vccd1 vccd1 _08701_/C sky130_fd_sc_hd__xnor2_1
X_09680_ _09678_/X _09679_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09680_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11677__A1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08631_ _09070_/A _09064_/B _09070_/C _08629_/Y vssd1 vssd1 vccd1 vccd1 _09068_/A
+ sky130_fd_sc_hd__a31o_4
X_06892_ _12723_/A _12722_/B vssd1 vssd1 vccd1 vccd1 _06892_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_55_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07345__A2 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08587__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11677__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08562_ reg1_val[0] _08544_/A _08544_/B _09600_/A _08544_/C vssd1 vssd1 vccd1 vccd1
+ _08563_/B sky130_fd_sc_hd__a32o_1
X_08493_ _10458_/A _08499_/B vssd1 vssd1 vccd1 vccd1 _08493_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_49_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07513_ _12762_/A fanout95/X fanout54/X _11347_/A vssd1 vssd1 vccd1 vccd1 _07514_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout156_A _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout16 _07277_/Y vssd1 vssd1 vccd1 vccd1 _07278_/B sky130_fd_sc_hd__buf_8
Xfanout27 _07389_/B vssd1 vssd1 vccd1 vccd1 fanout27/X sky130_fd_sc_hd__buf_6
Xfanout38 _06960_/X vssd1 vssd1 vccd1 vccd1 _08821_/B sky130_fd_sc_hd__buf_6
X_07444_ fanout57/X fanout52/X _10677_/B _07553_/A vssd1 vssd1 vccd1 vccd1 _07445_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout49 _07301_/Y vssd1 vssd1 vccd1 vccd1 _09752_/B sky130_fd_sc_hd__buf_8
X_07375_ _07655_/A _07655_/B _07372_/A vssd1 vssd1 vccd1 vccd1 _07377_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_127_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07805__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09114_ _11738_/S _09184_/B vssd1 vssd1 vccd1 vccd1 _09114_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11601__B2 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11601__A1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09045_ _09045_/A _09045_/B vssd1 vssd1 vccd1 vccd1 _09046_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10168__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10168__A1 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11117__B1 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09947_ _09947_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09948_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout69_A fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08497__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__A1 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__B2 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07336__A2 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09878_ _09879_/A _09879_/B vssd1 vssd1 vccd1 vccd1 _10018_/A sky130_fd_sc_hd__nor2_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ _08891_/B _08829_/B vssd1 vssd1 vccd1 vccd1 _08848_/A sky130_fd_sc_hd__or2_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _06645_/A _12243_/B1 _11838_/Y _06647_/B _11839_/X vssd1 vssd1 vccd1 vccd1
+ _11840_/X sky130_fd_sc_hd__o221a_1
XANTENNA__09105__B _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10891__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11771_ fanout37/X _12203_/A _12150_/A fanout35/X vssd1 vssd1 vccd1 vccd1 _11772_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10722_ _10722_/A _10722_/B vssd1 vssd1 vccd1 vccd1 _10724_/B sky130_fd_sc_hd__xnor2_2
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08049__A0 _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10653_ _10551_/A _10551_/B _10552_/A _10549_/X vssd1 vssd1 vccd1 vccd1 _10664_/A
+ sky130_fd_sc_hd__a31o_1
X_10584_ _10584_/A _10584_/B vssd1 vssd1 vccd1 vccd1 _10586_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12323_ _06856_/A _12322_/X _09192_/Y vssd1 vssd1 vccd1 vccd1 _12323_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12482__A _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12254_ fanout19/X _12304_/B _12255_/A vssd1 vssd1 vccd1 vccd1 _12254_/Y sky130_fd_sc_hd__o21bai_1
X_12185_ hold254/A _11398_/B _12240_/B _12184_/Y _11400_/A vssd1 vssd1 vccd1 vccd1
+ _12185_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_102_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11205_ _06698_/B _09188_/X _09191_/X _06696_/Y _11204_/X vssd1 vssd1 vccd1 vccd1
+ _11205_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08772__A1 _07023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08772__B2 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ fanout37/X _11704_/A _11688_/A fanout35/X vssd1 vssd1 vccd1 vccd1 _11137_/B
+ sky130_fd_sc_hd__o22a_1
X_11067_ _11067_/A _11067_/B _11067_/C vssd1 vssd1 vccd1 vccd1 _11068_/B sky130_fd_sc_hd__and3_1
XANTENNA__07742__C _08544_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _10018_/A _10018_/B _10018_/C vssd1 vssd1 vccd1 vccd1 _10019_/B sky130_fd_sc_hd__or3_1
XANTENNA__10882__A2 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11969_ _11969_/A _11969_/B vssd1 vssd1 vccd1 vccd1 _12216_/B sky130_fd_sc_hd__or2_1
XFILLER_0_86_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07160_ _07160_/A _07160_/B vssd1 vssd1 vccd1 vccd1 _07411_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07091_ _09968_/A _12370_/B _09362_/S vssd1 vssd1 vccd1 vccd1 _07093_/B sky130_fd_sc_hd__and3_2
XANTENNA__07263__A1 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07263__B2 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout206 _07763_/A vssd1 vssd1 vccd1 vccd1 _09898_/A sky130_fd_sc_hd__buf_8
Xfanout228 _06760_/X vssd1 vssd1 vccd1 vccd1 _07001_/C sky130_fd_sc_hd__clkbuf_4
Xfanout217 _09392_/S vssd1 vssd1 vccd1 vccd1 _09678_/S sky130_fd_sc_hd__clkbuf_8
X_09801_ _09638_/A _09638_/B _09636_/Y vssd1 vssd1 vccd1 vccd1 _09803_/B sky130_fd_sc_hd__o21a_2
Xfanout239 _09201_/X vssd1 vssd1 vccd1 vccd1 _12339_/B1 sky130_fd_sc_hd__clkbuf_4
X_07993_ _07994_/A _07994_/B vssd1 vssd1 vccd1 vccd1 _07993_/Y sky130_fd_sc_hd__nor2_1
X_09732_ _09733_/B _09733_/A vssd1 vssd1 vccd1 vccd1 _09732_/Y sky130_fd_sc_hd__nand2b_1
X_06944_ reg1_val[27] _06945_/B vssd1 vssd1 vccd1 vccd1 _06944_/X sky130_fd_sc_hd__xor2_2
XANTENNA__09206__A _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06875_ instruction[4] instruction[3] vssd1 vssd1 vccd1 vccd1 _09201_/B sky130_fd_sc_hd__nand2_2
X_09663_ _10230_/A _10230_/B _09661_/X _09662_/X vssd1 vssd1 vccd1 vccd1 _09664_/B
+ sky130_fd_sc_hd__o211a_2
X_08614_ _08614_/A _09009_/B vssd1 vssd1 vccd1 vccd1 _09054_/A sky130_fd_sc_hd__and2_1
X_09594_ _09465_/A _09465_/B _09462_/A vssd1 vssd1 vccd1 vccd1 _09597_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_82_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _08546_/B _08546_/C _08595_/A vssd1 vssd1 vccd1 vccd1 _08549_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08476_ _10155_/A _08476_/B vssd1 vssd1 vccd1 vccd1 _08506_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07427_ _07622_/B _07622_/A vssd1 vssd1 vccd1 vccd1 _07427_/Y sky130_fd_sc_hd__nand2b_1
X_07358_ _10015_/A _07358_/B vssd1 vssd1 vccd1 vccd1 _07362_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_33_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07289_ _07213_/Y _07222_/B _07220_/Y vssd1 vssd1 vccd1 vccd1 _07291_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09028_ _09028_/A _09028_/B vssd1 vssd1 vccd1 vccd1 _09076_/B sky130_fd_sc_hd__nand2_2
XANTENNA__11338__B1 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 hold260/A vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__buf_1
Xhold271 hold271/A vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07006__A1 _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold282 hold282/A vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 hold293/A vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
X_12941_ hold192/X _12955_/A2 _13168_/B1 hold173/X vssd1 vssd1 vccd1 vccd1 hold227/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06780__A3 _12568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12302__A2 _07277_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12872_ _12802_/X _12872_/B vssd1 vssd1 vccd1 vccd1 _13126_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11823_ _11821_/X _11822_/X _11823_/S vssd1 vssd1 vccd1 vccd1 _11824_/B sky130_fd_sc_hd__mux2_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11381__A _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _11754_/A _11754_/B vssd1 vssd1 vccd1 vccd1 _11754_/X sky130_fd_sc_hd__or2_1
XFILLER_0_68_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13015__B1 _13151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11685_ _11686_/A _11686_/B vssd1 vssd1 vccd1 vccd1 _11777_/B sky130_fd_sc_hd__nand2_1
X_10705_ _10705_/A _10705_/B _10705_/C vssd1 vssd1 vccd1 vccd1 _10706_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_126_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10636_ _09385_/C _10758_/B hold301/A vssd1 vssd1 vccd1 vccd1 _10636_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12369__A2 _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09786__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10567_ _10567_/A _10567_/B vssd1 vssd1 vccd1 vccd1 _10568_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13286_ _13310_/CLK _13286_/D vssd1 vssd1 vccd1 vccd1 hold284/A sky130_fd_sc_hd__dfxtp_1
X_10498_ _10498_/A _10498_/B vssd1 vssd1 vccd1 vccd1 _10498_/Y sky130_fd_sc_hd__nor2_1
X_12306_ _12348_/A _12305_/B _12301_/X vssd1 vssd1 vccd1 vccd1 _12307_/B sky130_fd_sc_hd__o21a_1
X_12237_ hold213/A _12237_/B vssd1 vssd1 vccd1 vccd1 _12288_/B sky130_fd_sc_hd__or2_1
X_12168_ _12221_/C _12166_/X _12167_/Y vssd1 vssd1 vccd1 vccd1 _12168_/X sky130_fd_sc_hd__o21a_1
X_12099_ _12099_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12215_/A sky130_fd_sc_hd__nor2_2
X_11119_ _11119_/A _11119_/B vssd1 vssd1 vccd1 vccd1 _11121_/B sky130_fd_sc_hd__xor2_1
X_06660_ _11756_/A _06660_/B vssd1 vssd1 vccd1 vccd1 _11739_/A sky130_fd_sc_hd__nor2_2
XANTENNA__11501__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06591_ _06591_/A _06591_/B vssd1 vssd1 vccd1 vccd1 _06605_/B sky130_fd_sc_hd__and2_1
X_08330_ _08360_/A _08330_/B vssd1 vssd1 vccd1 vccd1 _08371_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_604 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08261_ _08261_/A _08261_/B vssd1 vssd1 vccd1 vccd1 _08263_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_74_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07212_ _08589_/A _07212_/B vssd1 vssd1 vccd1 vccd1 _07222_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12765__C1 _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08192_ _09452_/A _08192_/B vssd1 vssd1 vccd1 vccd1 _08247_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07143_ _09180_/A reg1_val[1] _07105_/A vssd1 vssd1 vccd1 vccd1 _07144_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_14_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07074_ _08477_/B vssd1 vssd1 vccd1 vccd1 _07074_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08736__B2 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08736__A1 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11740__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07976_ _08658_/A vssd1 vssd1 vccd1 vccd1 _07976_/Y sky130_fd_sc_hd__inv_2
X_06927_ _12487_/S _06927_/B vssd1 vssd1 vccd1 vccd1 dest_mask[1] sky130_fd_sc_hd__nand2_8
XANTENNA__07155__S _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12296__A1 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09715_ _10273_/D _10273_/C vssd1 vssd1 vccd1 vccd1 _10002_/A sky130_fd_sc_hd__and2_1
XFILLER_0_97_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09646_ _09437_/A _09437_/B _09435_/Y vssd1 vssd1 vccd1 vccd1 _09649_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__08775__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06858_ _06858_/A _12357_/A _06834_/Y vssd1 vssd1 vccd1 vccd1 _06858_/X sky130_fd_sc_hd__or3b_1
X_06789_ reg1_val[2] _10249_/S vssd1 vssd1 vccd1 vccd1 _06789_/X sky130_fd_sc_hd__and2_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _09577_/A _09577_/B vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__xor2_4
X_08528_ _08528_/A _08528_/B vssd1 vssd1 vccd1 vccd1 _08529_/B sky130_fd_sc_hd__and2_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08459_ _08457_/X _09009_/A vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_65_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11470_ _11738_/S _11470_/B vssd1 vssd1 vccd1 vccd1 _11470_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09216__A2 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10421_ _10421_/A _10421_/B vssd1 vssd1 vccd1 vccd1 _10466_/A sky130_fd_sc_hd__and2_1
XANTENNA__12771__A2 _12781_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13140_ _13140_/A _13140_/B vssd1 vssd1 vccd1 vccd1 _13140_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10352_ _10353_/B _10353_/A vssd1 vssd1 vccd1 vccd1 _10352_/Y sky130_fd_sc_hd__nand2b_1
X_13071_ _13086_/A _13071_/B vssd1 vssd1 vccd1 vccd1 _13291_/D sky130_fd_sc_hd__and2_1
XFILLER_0_14_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12760__A _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10283_ _10283_/A _10283_/B vssd1 vssd1 vccd1 vccd1 _10284_/B sky130_fd_sc_hd__nor2_1
X_12022_ _12022_/A _12022_/B vssd1 vssd1 vccd1 vccd1 _12023_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10534__B2 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10534__A1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10280__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07950__A2 _10694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ _13169_/A hold204/X vssd1 vssd1 vccd1 vccd1 _13232_/D sky130_fd_sc_hd__and2_1
XANTENNA__10298__B1 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12855_ hold70/X hold295/A vssd1 vssd1 vccd1 vccd1 _13087_/B sky130_fd_sc_hd__nand2b_1
X_12786_ _12786_/A _12786_/B vssd1 vssd1 vccd1 vccd1 _12786_/Y sky130_fd_sc_hd__nand2_1
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11806_ _11888_/B _11806_/B vssd1 vssd1 vccd1 vccd1 _11809_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_126_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11737_ _06661_/C _11646_/X _06654_/A vssd1 vssd1 vccd1 vccd1 _11737_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07466__A1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07466__B2 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11668_ _11668_/A _11668_/B _11668_/C _11668_/D vssd1 vssd1 vccd1 vccd1 _11668_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06652__B _06653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10619_ _06732_/Y _10496_/Y _06734_/B vssd1 vssd1 vccd1 vccd1 _10619_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07218__A1 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07218__B2 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11599_ _11598_/B _11599_/B vssd1 vssd1 vccd1 vccd1 _11600_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_24_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10773__A1 _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13269_ _13277_/CLK _13269_/D vssd1 vssd1 vccd1 vccd1 hold128/A sky130_fd_sc_hd__dfxtp_1
X_07830_ _07829_/B _07829_/C _07829_/A vssd1 vssd1 vccd1 vccd1 _07831_/B sky130_fd_sc_hd__a21boi_4
X_07761_ _07783_/A _07783_/B vssd1 vssd1 vccd1 vccd1 _07781_/A sky130_fd_sc_hd__or2_2
XFILLER_0_37_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06712_ _06898_/A _06641_/A _12626_/B _06711_/X vssd1 vssd1 vccd1 vccd1 _07303_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__10289__B1 _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09500_ _09500_/A _09500_/B vssd1 vssd1 vccd1 vccd1 _09502_/B sky130_fd_sc_hd__xnor2_2
X_07692_ _07377_/B _07692_/B vssd1 vssd1 vccd1 vccd1 _07693_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08595__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06643_ _06641_/Y _06680_/B1 _06729_/B reg2_val[22] vssd1 vssd1 vccd1 vccd1 _07112_/B
+ sky130_fd_sc_hd__a2bb2o_2
X_09431_ _09432_/A _09432_/B vssd1 vssd1 vccd1 vccd1 _09596_/B sky130_fd_sc_hd__and2_1
X_06574_ instruction[1] instruction[2] instruction[25] pred_val vssd1 vssd1 vccd1
+ vccd1 _06574_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_87_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06827__B _07068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09362_ _09163_/X _09165_/X _09362_/S vssd1 vssd1 vccd1 vccd1 _09362_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08313_ _08309_/X _08313_/B vssd1 vssd1 vccd1 vccd1 _08362_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout236_A _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_11 reg1_val[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_22 reg1_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09293_ _07475_/A _07475_/B _07472_/A vssd1 vssd1 vccd1 vccd1 _09310_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_117_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08244_ _08244_/A _08244_/B vssd1 vssd1 vccd1 vccd1 _08246_/A sky130_fd_sc_hd__nand2_1
XANTENNA_55 reg2_val[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_44 reg2_val[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_66 reg2_val[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_33 reg2_val[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08175_ _08774_/A2 fanout82/X _08672_/B _08774_/B1 vssd1 vssd1 vccd1 vccd1 _08176_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_77 reg1_val[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12753__A2 _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07126_ _07157_/A _07126_/B vssd1 vssd1 vccd1 vccd1 _07129_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07057_ _10155_/A _07045_/Y _07056_/Y vssd1 vssd1 vccd1 vccd1 _07057_/X sky130_fd_sc_hd__o21a_2
XFILLER_0_30_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07674__A _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07959_ _08420_/B _12752_/A fanout84/X _08854_/B2 vssd1 vssd1 vccd1 vccd1 _07960_/B
+ sky130_fd_sc_hd__o22a_1
X_10970_ _10863_/A _10861_/Y _06715_/B vssd1 vssd1 vccd1 vccd1 _10970_/X sky130_fd_sc_hd__o21a_1
X_09629_ _09629_/A _09629_/B vssd1 vssd1 vccd1 vccd1 _09632_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_78_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ _12640_/A _12640_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[15] sky130_fd_sc_hd__nor2_8
XANTENNA__08645__B1 _08774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12571_ _12570_/A _12567_/Y _12569_/B vssd1 vssd1 vccd1 vccd1 _12575_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_108_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12992__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire201 wire201/A vssd1 vssd1 vccd1 vccd1 wire201/X sky130_fd_sc_hd__clkbuf_4
X_11522_ _11522_/A _11522_/B vssd1 vssd1 vccd1 vccd1 _11526_/B sky130_fd_sc_hd__xor2_1
XANTENNA__10452__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11453_ _11453_/A _11453_/B vssd1 vssd1 vccd1 vccd1 _11455_/B sky130_fd_sc_hd__xor2_1
X_10404_ _10357_/A _10355_/X _10354_/X vssd1 vssd1 vccd1 vccd1 _10485_/A sky130_fd_sc_hd__a21oi_4
X_13123_ hold277/A _13122_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13123_/X sky130_fd_sc_hd__mux2_1
X_11384_ _06865_/C _11383_/X _12277_/B1 vssd1 vssd1 vccd1 vccd1 _11384_/Y sky130_fd_sc_hd__a21oi_1
X_10335_ fanout77/X _10557_/B fanout13/X _11704_/A vssd1 vssd1 vccd1 vccd1 _10336_/B
+ sky130_fd_sc_hd__o22a_1
X_13054_ hold266/X _13053_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13054_/X sky130_fd_sc_hd__mux2_1
X_10266_ _10266_/A _10266_/B vssd1 vssd1 vccd1 vccd1 _10266_/Y sky130_fd_sc_hd__xnor2_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12005_ _12005_/A _12069_/B vssd1 vssd1 vccd1 vccd1 _12005_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_108_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10197_ _11704_/A _10557_/B fanout13/X _11688_/A vssd1 vssd1 vccd1 vccd1 _10198_/B
+ sky130_fd_sc_hd__o22a_1
X_12907_ hold228/X _12947_/A2 _12947_/B1 _13224_/Q vssd1 vssd1 vccd1 vccd1 hold229/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ _12822_/B _13043_/B _12820_/X vssd1 vssd1 vccd1 vccd1 _13048_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_69_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10691__B1 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12769_ hold5/X _12778_/B _12768_/Y _13147_/A vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__o211a_1
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06663__A _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10443__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10994__B2 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12735__A2 _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09980_ hold189/A _09980_/B vssd1 vssd1 vccd1 vccd1 _09980_/Y sky130_fd_sc_hd__nand2_1
X_08931_ _08932_/A _08932_/B vssd1 vssd1 vccd1 vccd1 _08935_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_58_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13160__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08862_ _08862_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _08864_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07813_ _07809_/A _07809_/B _07847_/A vssd1 vssd1 vccd1 vccd1 _07833_/A sky130_fd_sc_hd__o21bai_4
XANTENNA__06717__A3 _12620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08793_ _08713_/A _08713_/B _08711_/Y vssd1 vssd1 vccd1 vccd1 _08794_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_74_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout186_A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07744_ _08394_/A _07744_/B _07744_/C vssd1 vssd1 vccd1 vccd1 _07747_/B sky130_fd_sc_hd__or3_1
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12120__B1 _09200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ _07676_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _07675_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12559__B _12560_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06557__B _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06626_ _06649_/A _12637_/B vssd1 vssd1 vccd1 vccd1 _06626_/Y sky130_fd_sc_hd__nor2_1
X_09414_ _08821_/B _10144_/B2 _10064_/B2 fanout36/X vssd1 vssd1 vccd1 vccd1 _09415_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06557_ instruction[21] _06915_/B vssd1 vssd1 vccd1 vccd1 _06557_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09345_ _09127_/X _09131_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09345_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09276_ _09618_/A1 _12782_/A fanout20/X _09618_/B2 vssd1 vssd1 vccd1 vccd1 _09277_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_35_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10434__B1 _07325_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07850__A1 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08227_ _08284_/A vssd1 vssd1 vccd1 vccd1 _08227_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07850__B2 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09884__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08158_ _08158_/A _08158_/B vssd1 vssd1 vccd1 vccd1 _08167_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_120_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08089_ _08089_/A _08089_/B vssd1 vssd1 vccd1 vccd1 _08150_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07109_ _09764_/A _07110_/B vssd1 vssd1 vccd1 vccd1 _08572_/B sky130_fd_sc_hd__and2_2
X_10120_ _12124_/B _10252_/B hold228/A vssd1 vssd1 vccd1 vccd1 _10120_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13151__A2 _13151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10051_ _10052_/B _10052_/A vssd1 vssd1 vccd1 vccd1 _10194_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07366__B1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10953_ _10953_/A _10953_/B _10953_/C vssd1 vssd1 vccd1 vccd1 _10954_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_97_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10884_ _10875_/Y _10876_/X _10883_/Y _09115_/X _10882_/X vssd1 vssd1 vccd1 vccd1
+ _10884_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12623_ _12623_/A _12623_/B _12623_/C vssd1 vssd1 vccd1 vccd1 _12624_/B sky130_fd_sc_hd__nand3_1
X_12554_ _12554_/A _12554_/B vssd1 vssd1 vccd1 vccd1 new_PC[26] sky130_fd_sc_hd__xnor2_4
XANTENNA__11820__C _11820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11505_ _11618_/B _11505_/B vssd1 vssd1 vccd1 vccd1 _11516_/A sky130_fd_sc_hd__or2_1
XFILLER_0_124_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12485_ _12485_/A _12485_/B _12485_/C vssd1 vssd1 vccd1 vccd1 _12486_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11436_ _11437_/A _11437_/B vssd1 vssd1 vccd1 vccd1 _11438_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12424__S _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ _11367_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _11369_/C sky130_fd_sc_hd__xor2_1
X_13106_ _13116_/A hold261/X vssd1 vssd1 vccd1 vccd1 _13298_/D sky130_fd_sc_hd__and2_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10318_ _10433_/C _10433_/D vssd1 vssd1 vccd1 vccd1 _10320_/C sky130_fd_sc_hd__xnor2_1
X_11298_ hold294/A _11398_/B _11397_/B _11400_/A vssd1 vssd1 vccd1 vccd1 _11298_/Y
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__13142__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13037_ hold246/X _12721_/B _13036_/X _12722_/A vssd1 vssd1 vccd1 vccd1 hold247/A
+ sky130_fd_sc_hd__a22o_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10249_ _09676_/X _09679_/X _10249_/S vssd1 vssd1 vccd1 vccd1 _10249_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07357__B1 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07460_ fanout77/X _10156_/A1 fanout62/X _10156_/B2 vssd1 vssd1 vccd1 vccd1 _07461_/B
+ sky130_fd_sc_hd__o22a_1
X_07391_ _08544_/C _12087_/A vssd1 vssd1 vccd1 vccd1 _07393_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09130_ _09122_/X _09129_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09130_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09061_ _09061_/A _09061_/B vssd1 vssd1 vccd1 vccd1 _11285_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_71_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08012_ _08013_/A _08013_/B vssd1 vssd1 vccd1 vccd1 _08806_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11916__B1 _09200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07001__B _12370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08388__A2 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09585__B2 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09585__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11392__A1 _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_95 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06840__B _07126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09963_ _09859_/X _10002_/C _09110_/X vssd1 vssd1 vccd1 vccd1 _09963_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10195__A2 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13133__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08914_ _08914_/A _08914_/B _08914_/C vssd1 vssd1 vccd1 vccd1 _08916_/A sky130_fd_sc_hd__and3_1
XFILLER_0_110_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09894_ _10155_/A _09894_/B vssd1 vssd1 vccd1 vccd1 _09900_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09888__A2 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__A1 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07899__B2 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08845_ _08899_/B _08845_/B vssd1 vssd1 vccd1 vccd1 _08847_/B sky130_fd_sc_hd__and2_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08776_ _12760_/A _08477_/B _08776_/B1 _09925_/A1 vssd1 vssd1 vccd1 vccd1 _08777_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08560__A2 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07727_ _07727_/A _07727_/B _07727_/C vssd1 vssd1 vccd1 vccd1 _07738_/A sky130_fd_sc_hd__and3_1
XFILLER_0_79_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07658_ _09772_/A _09295_/A _07969_/A _08681_/A vssd1 vssd1 vccd1 vccd1 _07659_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07520__B1 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06609_ _06607_/Y _06680_/B1 _06778_/B reg2_val[27] vssd1 vssd1 vccd1 vccd1 _07434_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_07589_ _07589_/A _07589_/B vssd1 vssd1 vccd1 vccd1 _07590_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_48_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09328_ _09328_/A _09328_/B vssd1 vssd1 vccd1 vccd1 _09331_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09273__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09259_ _10156_/A1 _10557_/A fanout58/X _10156_/B2 vssd1 vssd1 vccd1 vccd1 _09260_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12270_ _12312_/B _12270_/B vssd1 vssd1 vccd1 vccd1 _12317_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_31_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12752__B _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ _11221_/A _11221_/B vssd1 vssd1 vccd1 vccd1 _11222_/C sky130_fd_sc_hd__xor2_1
XANTENNA__10553__A _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11152_ _11152_/A _11152_/B vssd1 vssd1 vccd1 vccd1 _11166_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13124__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10103_ _10617_/A _10104_/B _10104_/C vssd1 vssd1 vccd1 vccd1 _10105_/B sky130_fd_sc_hd__o21a_1
X_11083_ _06705_/A _11081_/X _11082_/Y vssd1 vssd1 vccd1 vccd1 _11083_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07862__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _09898_/A _09897_/Y _09899_/Y vssd1 vssd1 vccd1 vccd1 _10040_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__08303__A2 _08572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11985_ reg1_val[24] curr_PC[24] vssd1 vssd1 vccd1 vccd1 _11986_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_105_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08693__A _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10936_ _10937_/B _10937_/A vssd1 vssd1 vccd1 vccd1 _11054_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_14_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10867_ _10251_/S _09691_/X _10866_/X vssd1 vssd1 vccd1 vccd1 _10867_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_73_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12606_ reg1_val[10] _12607_/B vssd1 vssd1 vccd1 vccd1 _12617_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13060__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10798_ _10553_/A _11794_/A _11704_/A fanout33/X vssd1 vssd1 vccd1 vccd1 _10799_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09264__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07814__A1 _10281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07814__B2 _10149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12537_ reg1_val[24] curr_PC[24] _12556_/S vssd1 vssd1 vccd1 vccd1 _12538_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_30_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12468_ _12626_/B _12468_/B vssd1 vssd1 vccd1 vccd1 _12469_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11419_ _12301_/A fanout47/X _11603_/A fanout19/X vssd1 vssd1 vccd1 vccd1 _11420_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_111_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12399_ _12408_/A _12399_/B vssd1 vssd1 vccd1 vccd1 _12401_/C sky130_fd_sc_hd__nand2_1
XANTENNA__10177__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13115__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06960_ _06960_/A _12078_/A vssd1 vssd1 vccd1 vccd1 _06960_/X sky130_fd_sc_hd__or2_1
X_06891_ _12722_/A _12723_/B vssd1 vssd1 vccd1 vccd1 _06891_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07772__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11677__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08630_ _08630_/A _08630_/B vssd1 vssd1 vccd1 vccd1 _09070_/C sky130_fd_sc_hd__xor2_4
XFILLER_0_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08561_ _08589_/A _08561_/B vssd1 vssd1 vccd1 vccd1 _08570_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11834__C1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08492_ _08492_/A _08492_/B vssd1 vssd1 vccd1 vccd1 _08499_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07512_ _07512_/A _07512_/B vssd1 vssd1 vccd1 vccd1 _07516_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_119_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout17 _12786_/A vssd1 vssd1 vccd1 vccd1 _12301_/A sky130_fd_sc_hd__clkbuf_8
Xfanout28 _07098_/Y vssd1 vssd1 vccd1 vccd1 _07389_/B sky130_fd_sc_hd__buf_8
X_07443_ _10894_/A _07443_/B vssd1 vssd1 vccd1 vccd1 _07447_/A sky130_fd_sc_hd__xor2_1
XANTENNA__12929__A2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12329__S _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06835__B _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout149_A _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout39 _12349_/B vssd1 vssd1 vccd1 vccd1 _12304_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_9_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07374_ _09580_/A _07374_/B vssd1 vssd1 vccd1 vccd1 _07655_/B sky130_fd_sc_hd__xnor2_1
X_09113_ _09201_/B instruction[5] _06849_/X vssd1 vssd1 vccd1 vccd1 _09218_/C sky130_fd_sc_hd__or3b_1
XANTENNA__07805__B2 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07805__A1 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11601__A2 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09044_ _10104_/B _10104_/C vssd1 vssd1 vccd1 vccd1 _09046_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12572__B _12573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10168__A2 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11117__A1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09946_ _09946_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _09946_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07682__A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11117__B2 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10876__B1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08533__A2 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09877_ _09758_/B _09761_/B _09758_/A vssd1 vssd1 vccd1 vccd1 _09879_/B sky130_fd_sc_hd__o21ba_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07741__B1 _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08828_ _08827_/B _08828_/B vssd1 vssd1 vccd1 vccd1 _08829_/B sky130_fd_sc_hd__and2b_1
X_08759_ _09621_/A _08759_/B vssd1 vssd1 vccd1 vccd1 _08761_/B sky130_fd_sc_hd__xnor2_2
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ _12206_/A _11770_/B vssd1 vssd1 vccd1 vccd1 _11774_/B sky130_fd_sc_hd__xnor2_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ _10722_/B _10722_/A vssd1 vssd1 vccd1 vccd1 _10721_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11840__A2 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06745__B _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10548__A _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10652_ _10600_/A _10600_/B _10598_/Y vssd1 vssd1 vccd1 vccd1 _10725_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10982__S _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10583_ _11125_/A _10583_/B vssd1 vssd1 vccd1 vccd1 _10584_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12322_ _06856_/B _12321_/X _12322_/S vssd1 vssd1 vccd1 vccd1 _12322_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_36_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11379__A _11379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12253_ _12255_/B _12253_/B vssd1 vssd1 vccd1 vccd1 _12257_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11204_ _07178_/A _06928_/X _11099_/B reg1_val[15] vssd1 vssd1 vccd1 vccd1 _11204_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_12184_ _11398_/B _12240_/B hold254/A vssd1 vssd1 vccd1 vccd1 _12184_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08772__A2 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ _12255_/B _11135_/B vssd1 vssd1 vccd1 vccd1 _11139_/A sky130_fd_sc_hd__xnor2_1
X_11066_ _11068_/A vssd1 vssd1 vccd1 vccd1 _11066_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09182__C1 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10017_ _10018_/A _10018_/B _10018_/C vssd1 vssd1 vccd1 vccd1 _10019_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11968_ _11811_/X _11969_/B _11966_/Y vssd1 vssd1 vccd1 vccd1 _11968_/Y sky130_fd_sc_hd__o21bai_1
X_11899_ _11848_/X _11972_/D _12223_/B1 vssd1 vssd1 vccd1 vccd1 _11899_/Y sky130_fd_sc_hd__o21ai_1
X_10919_ _11604_/A _10919_/B vssd1 vssd1 vccd1 vccd1 _10920_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10458__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11988__S _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07799__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07090_ _07090_/A _07090_/B vssd1 vssd1 vccd1 vccd1 _07090_/X sky130_fd_sc_hd__or2_2
XFILLER_0_42_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07263__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07992_ _08775_/A _07992_/B vssd1 vssd1 vccd1 vccd1 _07994_/B sky130_fd_sc_hd__xnor2_4
Xfanout229 _11746_/A vssd1 vssd1 vccd1 vccd1 _11197_/S sky130_fd_sc_hd__clkbuf_8
Xfanout207 _07763_/A vssd1 vssd1 vccd1 vccd1 _09467_/A sky130_fd_sc_hd__buf_8
Xfanout218 _09392_/S vssd1 vssd1 vccd1 vccd1 _09676_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09800_ _09593_/A _09593_/B _09591_/Y vssd1 vssd1 vccd1 vccd1 _09803_/A sky130_fd_sc_hd__a21boi_4
X_06943_ reg1_val[26] _07087_/B _07087_/C _07086_/C _07165_/A vssd1 vssd1 vccd1 vccd1
+ _06945_/B sky130_fd_sc_hd__o41a_4
X_09731_ _09731_/A _09731_/B vssd1 vssd1 vccd1 vccd1 _09733_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_66_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07723__B1 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10858__B1 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06874_ _09200_/A _06872_/X _06873_/Y _06928_/D vssd1 vssd1 vccd1 vccd1 _06874_/X
+ sky130_fd_sc_hd__o211a_1
X_09662_ _07705_/X _08994_/Y _09660_/C _09816_/A _07706_/X vssd1 vssd1 vccd1 vccd1
+ _09662_/X sky130_fd_sc_hd__a2111o_1
X_08613_ _09010_/A _09009_/B vssd1 vssd1 vccd1 vccd1 _08613_/X sky130_fd_sc_hd__and2_1
X_09593_ _09593_/A _09593_/B vssd1 vssd1 vccd1 vccd1 _09640_/A sky130_fd_sc_hd__xor2_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08544_ _08544_/A _08544_/B _08544_/C vssd1 vssd1 vccd1 vccd1 _08546_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12567__B _12568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08475_ _07058_/A _08825_/A2 _09476_/A _08532_/B vssd1 vssd1 vccd1 vccd1 _08476_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07426_ _07426_/A _07426_/B vssd1 vssd1 vccd1 vccd1 _07622_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09228__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07357_ _08681_/A _08837_/B2 _12736_/A _09295_/A vssd1 vssd1 vccd1 vccd1 _07358_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09027_ _08633_/Y _08641_/Y _09025_/X _09026_/Y _08639_/Y vssd1 vssd1 vccd1 vccd1
+ _09028_/B sky130_fd_sc_hd__o32a_2
XANTENNA__06581__A _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07288_ _07355_/A _07355_/B vssd1 vssd1 vccd1 vccd1 _07356_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11338__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11338__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold261 hold261/A vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold250 hold250/A vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__buf_1
Xhold283 hold283/A vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold294 hold294/A vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06664__A2_N _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout81_A _07312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09929_ _09929_/A _09929_/B vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12940_ _12946_/A hold193/X vssd1 vssd1 vccd1 vccd1 hold194/A sky130_fd_sc_hd__and2_1
XANTENNA__12302__A3 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12871_ hold252/X hold86/X vssd1 vssd1 vccd1 vccd1 _12872_/B sky130_fd_sc_hd__nand2b_1
X_11822_ _11739_/A _11736_/X _06826_/Y vssd1 vssd1 vccd1 vccd1 _11822_/X sky130_fd_sc_hd__o21a_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08674__C _08674_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ hold221/A _12187_/A1 _11835_/B _11920_/C1 vssd1 vssd1 vccd1 vccd1 _11754_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10278__A _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11684_ _11684_/A vssd1 vssd1 vccd1 vccd1 _11686_/B sky130_fd_sc_hd__inv_2
X_10704_ _10705_/B _10705_/C _10705_/A vssd1 vssd1 vccd1 vccd1 _10706_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_125_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10635_ hold272/A _10635_/B vssd1 vssd1 vccd1 vccd1 _10758_/B sky130_fd_sc_hd__or2_1
XFILLER_0_71_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11026__B1 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08442__B2 _10035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08442__A1 _10149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ _12348_/A _12305_/B vssd1 vssd1 vccd1 vccd1 _12305_/Y sky130_fd_sc_hd__nor2_1
X_10566_ _10567_/A _10567_/B vssd1 vssd1 vccd1 vccd1 _10705_/C sky130_fd_sc_hd__and2_1
XFILLER_0_23_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13285_ _13310_/CLK _13285_/D vssd1 vssd1 vccd1 vccd1 hold288/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10497_ _06802_/Y _10496_/Y _11647_/S vssd1 vssd1 vccd1 vccd1 _10498_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_11_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12236_ _12361_/B _12234_/Y _12235_/Y _09205_/B vssd1 vssd1 vccd1 vccd1 _12236_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_32_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12167_ _12221_/C _12166_/X _09110_/X vssd1 vssd1 vccd1 vccd1 _12167_/Y sky130_fd_sc_hd__a21oi_1
X_11118_ _11853_/A _11118_/B vssd1 vssd1 vccd1 vccd1 _11119_/B sky130_fd_sc_hd__xnor2_1
X_12098_ _12098_/A _12098_/B _12098_/C vssd1 vssd1 vccd1 vccd1 _12099_/B sky130_fd_sc_hd__and3_1
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11501__A1 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11049_ _10931_/B _10938_/B _10929_/Y vssd1 vssd1 vccd1 vccd1 _11060_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__11501__B2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07181__A1 _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06590_ reg1_val[28] _12250_/A vssd1 vssd1 vccd1 vccd1 _06591_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09458__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08130__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ _08260_/A _08260_/B vssd1 vssd1 vccd1 vccd1 _08263_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__13006__A1 _07005_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08191_ _08841_/B2 _08477_/B _08776_/B1 _08837_/B2 vssd1 vssd1 vccd1 vccd1 _08192_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_62_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07211_ fanout22/X _08588_/B _10677_/A _09273_/A1 vssd1 vssd1 vccd1 vccd1 _07212_/B
+ sky130_fd_sc_hd__o22a_1
X_07142_ _07160_/A _07160_/B vssd1 vssd1 vccd1 vccd1 _07383_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09630__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07073_ _07073_/A _07073_/B vssd1 vssd1 vccd1 vccd1 _07073_/X sky130_fd_sc_hd__or2_2
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08736__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07975_ _07977_/A _07977_/B _07977_/C vssd1 vssd1 vccd1 vccd1 _08658_/A sky130_fd_sc_hd__a21o_1
X_06926_ _06687_/A _06923_/B _06923_/C is_load _11823_/S vssd1 vssd1 vccd1 vccd1 _06927_/B
+ sky130_fd_sc_hd__a32o_2
X_09714_ _12005_/A _09710_/X _09711_/X _09713_/Y vssd1 vssd1 vccd1 vccd1 dest_val[3]
+ sky130_fd_sc_hd__a22o_4
XANTENNA__07960__A _08232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06857_ _06856_/A _06856_/B _06834_/Y vssd1 vssd1 vccd1 vccd1 _06857_/X sky130_fd_sc_hd__o21a_1
X_09645_ _09645_/A _09645_/B vssd1 vssd1 vccd1 vccd1 _09650_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12048__A2 _09079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06788_ _09383_/A _09380_/B _06787_/X vssd1 vssd1 vccd1 vccd1 _06788_/X sky130_fd_sc_hd__a21o_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ _09576_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09577_/B sky130_fd_sc_hd__nor2_2
X_08527_ _08527_/A _08527_/B vssd1 vssd1 vccd1 vccd1 _08609_/A sky130_fd_sc_hd__xnor2_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08458_ _08457_/A _08457_/B _08457_/C vssd1 vssd1 vccd1 vccd1 _09009_/A sky130_fd_sc_hd__a21o_1
X_07409_ _07409_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07412_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11008__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08389_ _10453_/A _08389_/B vssd1 vssd1 vccd1 vccd1 _08390_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10420_ _10420_/A _10420_/B _10420_/C vssd1 vssd1 vccd1 vccd1 _10421_/B sky130_fd_sc_hd__or3_1
XANTENNA__08424__A1 _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10351_ _10351_/A _10351_/B vssd1 vssd1 vccd1 vccd1 _10353_/B sky130_fd_sc_hd__xnor2_1
X_13070_ hold276/X _12721_/B _13069_/X _12722_/A vssd1 vssd1 vccd1 vccd1 _13071_/B
+ sky130_fd_sc_hd__a22o_1
X_10282_ _10281_/A _10551_/B _10281_/C vssd1 vssd1 vccd1 vccd1 _10283_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08188__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12021_ fanout35/X _12301_/A fanout8/X fanout37/X vssd1 vssd1 vccd1 vccd1 _12022_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10534__A2 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ hold180/X _12955_/A2 _13151_/A2 hold203/X vssd1 vssd1 vccd1 vccd1 hold204/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10298__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__A1 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12854_ _13082_/A _13083_/A _13082_/B vssd1 vssd1 vccd1 vccd1 _13088_/A sky130_fd_sc_hd__a21bo_1
X_12785_ hold21/X _12786_/B _12784_/Y _13166_/A vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__o211a_1
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11247__B1 _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11805_ _11805_/A _11805_/B vssd1 vssd1 vccd1 vccd1 _11806_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_96_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11736_ _06661_/C _06824_/X _06827_/Y vssd1 vssd1 vccd1 vccd1 _11736_/X sky130_fd_sc_hd__o21a_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07466__A2 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_216 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11667_ _11658_/Y _11659_/X _11663_/X vssd1 vssd1 vccd1 vccd1 _11668_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_64_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10618_ _10618_/A _10618_/B vssd1 vssd1 vccd1 vccd1 _10618_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07218__A2 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11598_ _11599_/B _11598_/B vssd1 vssd1 vccd1 vccd1 _11706_/B sky130_fd_sc_hd__and2b_1
X_10549_ _10550_/A _10550_/B vssd1 vssd1 vccd1 vccd1 _10549_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_12_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10773__A2 _10769_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13268_ _13277_/CLK hold112/X vssd1 vssd1 vccd1 vccd1 hold110/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09376__C1 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13199_ _13310_/CLK hold72/X vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfxtp_1
X_12219_ _12313_/A _12218_/Y _12217_/X _12216_/X vssd1 vssd1 vccd1 vccd1 _12220_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07760_ _08857_/A _07760_/B vssd1 vssd1 vccd1 vccd1 _07783_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_47_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11486__B1 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06711_ reg2_val[12] _06729_/B vssd1 vssd1 vccd1 vccd1 _06711_/X sky130_fd_sc_hd__and2_1
XFILLER_0_2_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12398__A _12573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07691_ _08969_/A _08969_/B _07654_/Y vssd1 vssd1 vccd1 vccd1 _07700_/B sky130_fd_sc_hd__a21oi_2
X_09430_ _10565_/A _09430_/B vssd1 vssd1 vccd1 vccd1 _09432_/B sky130_fd_sc_hd__xnor2_1
X_06642_ reg2_val[22] _06729_/B _06680_/B1 _06641_/Y vssd1 vssd1 vccd1 vccd1 _07111_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_78_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06573_ instruction[25] _06633_/B vssd1 vssd1 vccd1 vccd1 _12560_/B sky130_fd_sc_hd__and2_4
X_09361_ _09358_/X _09360_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09361_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08312_ _08309_/B _08309_/C _08309_/A vssd1 vssd1 vccd1 vccd1 _08313_/B sky130_fd_sc_hd__a21o_1
X_09292_ _09292_/A _09292_/B vssd1 vssd1 vccd1 vccd1 _09312_/A sky130_fd_sc_hd__xnor2_1
X_08243_ _08243_/A _08243_/B vssd1 vssd1 vccd1 vccd1 _08244_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_12 reg1_val[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 reg1_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout131_A _09742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout229_A _11746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_45 reg2_val[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_34 reg2_val[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 reg2_val[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08174_ _08243_/A _08243_/B vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__or2_1
XFILLER_0_43_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_67 _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_78 reg1_val[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07125_ _07157_/A _07126_/B vssd1 vssd1 vccd1 vccd1 _07128_/D sky130_fd_sc_hd__and2_1
XANTENNA__11410__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10764__A2 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07056_ _10155_/A _07056_/B vssd1 vssd1 vccd1 vccd1 _07056_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_30_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07958_ _07958_/A _07958_/B vssd1 vssd1 vccd1 vccd1 _07980_/A sky130_fd_sc_hd__xnor2_1
X_06909_ instruction[27] _06915_/B vssd1 vssd1 vccd1 vccd1 _06909_/X sky130_fd_sc_hd__or2_1
X_07889_ _08841_/A1 _08854_/B2 _08835_/B1 _08420_/B vssd1 vssd1 vccd1 vccd1 _07891_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout44_A _11147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09628_ _09628_/A _09628_/B vssd1 vssd1 vccd1 vccd1 _09629_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_84_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09559_ _09559_/A wire3/X _09559_/C _09559_/D vssd1 vssd1 vccd1 vccd1 _10273_/D sky130_fd_sc_hd__and4_1
XFILLER_0_38_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _12570_/A _12570_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[2] sky130_fd_sc_hd__xnor2_4
XANTENNA__08645__A1 _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08645__B2 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09410__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10452__A1 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11521_ _11522_/A _11522_/B vssd1 vssd1 vccd1 vccd1 _11616_/A sky130_fd_sc_hd__and2b_1
XANTENNA__10452__B2 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08026__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11452_ _11453_/A _11453_/B vssd1 vssd1 vccd1 vccd1 _11547_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_104_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11383_ _06818_/X _11382_/X _11738_/S vssd1 vssd1 vccd1 vccd1 _11383_/X sky130_fd_sc_hd__mux2_1
X_10403_ _10617_/A _10524_/A vssd1 vssd1 vccd1 vccd1 _10403_/X sky130_fd_sc_hd__or2_1
XFILLER_0_33_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13122_ _13122_/A _13122_/B vssd1 vssd1 vccd1 vccd1 _13122_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10334_ _10334_/A _10334_/B vssd1 vssd1 vccd1 vccd1 _10337_/A sky130_fd_sc_hd__nor2_1
X_13053_ _13053_/A _13053_/B vssd1 vssd1 vccd1 vccd1 _13053_/Y sky130_fd_sc_hd__xnor2_1
X_10265_ _10263_/Y _10265_/B vssd1 vssd1 vccd1 vccd1 _10266_/B sky130_fd_sc_hd__nand2b_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12901__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12004_ curr_PC[24] _12070_/C vssd1 vssd1 vccd1 vccd1 _12069_/B sky130_fd_sc_hd__and2_1
X_10196_ _10555_/A _10196_/B vssd1 vssd1 vccd1 vccd1 _10200_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07136__A1 _07153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12906_ _12946_/A hold190/X vssd1 vssd1 vccd1 vccd1 hold191/A sky130_fd_sc_hd__and2_1
XANTENNA__10140__B1 _10137_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ _12825_/B _13039_/B _12823_/X vssd1 vssd1 vccd1 vccd1 _13043_/B sky130_fd_sc_hd__a21o_1
XANTENNA__10691__A1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10691__B2 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _12768_/A _12778_/B vssd1 vssd1 vccd1 vccd1 _12768_/Y sky130_fd_sc_hd__nand2_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06663__B _12578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12699_ _12700_/B _12700_/C _12700_/A vssd1 vssd1 vccd1 vccd1 _12705_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__10443__B2 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10443__A1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11719_ _11719_/A _11719_/B vssd1 vssd1 vccd1 vccd1 _11722_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12196__B2 _12382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08930_ _08930_/A _08930_/B vssd1 vssd1 vccd1 vccd1 _08932_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_58_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08861_ _08861_/A _08861_/B vssd1 vssd1 vccd1 vccd1 _08862_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07812_ _07846_/B _07812_/B vssd1 vssd1 vccd1 vccd1 _07847_/A sky130_fd_sc_hd__and2b_1
X_08792_ _08792_/A _08792_/B vssd1 vssd1 vccd1 vccd1 _08794_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07180__A_N _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07743_ _07744_/B _07744_/C _08394_/A vssd1 vssd1 vccd1 vccd1 _07747_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout179_A _12742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07674_ _09622_/A _07674_/B vssd1 vssd1 vccd1 vccd1 _08831_/A sky130_fd_sc_hd__xor2_2
XANTENNA__06838__B _07153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06625_ instruction[40] _06633_/B vssd1 vssd1 vccd1 vccd1 _12637_/B sky130_fd_sc_hd__and2_4
XFILLER_0_66_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09413_ _09413_/A _09413_/B vssd1 vssd1 vccd1 vccd1 _09416_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06556_ instruction[13] _06552_/X _06555_/X _06678_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[2]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09344_ _09124_/X _09126_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09344_/X sky130_fd_sc_hd__mux2_1
XANTENNA__06573__B _06633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09275_ _09280_/A vssd1 vssd1 vccd1 vccd1 _09275_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_35_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10434__B2 _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08226_ _08311_/A _08226_/B vssd1 vssd1 vccd1 vccd1 _08284_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08157_ _08157_/A _08212_/A vssd1 vssd1 vccd1 vccd1 _08167_/A sky130_fd_sc_hd__nand2_2
XANTENNA__07850__A2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07108_ _08589_/A _07115_/B vssd1 vssd1 vccd1 vccd1 _07110_/B sky130_fd_sc_hd__or2_1
XANTENNA__11934__B2 _11780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08088_ _08773_/A _08088_/B vssd1 vssd1 vccd1 vccd1 _08150_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07063__B1 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07039_ reg1_val[7] _07039_/B vssd1 vssd1 vccd1 vccd1 _08415_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_101_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10050_ _10050_/A _10050_/B vssd1 vssd1 vccd1 vccd1 _10052_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07366__A1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07366__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11935__A _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08315__B1 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10952_ _10953_/A _10953_/B _10953_/C vssd1 vssd1 vccd1 vccd1 _11067_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12766__A _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10883_ _10251_/S _09681_/X _09214_/A vssd1 vssd1 vccd1 vccd1 _10883_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_66_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12622_ _12623_/A _12623_/B _12623_/C vssd1 vssd1 vccd1 vccd1 _12629_/B sky130_fd_sc_hd__a21o_1
X_12553_ _12546_/B _12548_/B _12546_/A vssd1 vssd1 vccd1 vccd1 _12554_/B sky130_fd_sc_hd__o21ba_2
XFILLER_0_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11504_ _11503_/B _11504_/B vssd1 vssd1 vccd1 vccd1 _11505_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_19_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12484_ _12485_/A _12485_/B _12485_/C vssd1 vssd1 vccd1 vccd1 _12490_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11925__A1 _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11435_ _11435_/A _11435_/B vssd1 vssd1 vccd1 vccd1 _11437_/B sky130_fd_sc_hd__and2_1
XFILLER_0_123_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11925__B2 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11366_ _11367_/A _11367_/B vssd1 vssd1 vccd1 vccd1 _11457_/B sky130_fd_sc_hd__nand2b_1
X_13105_ hold260/X _13165_/A2 _13104_/X _13146_/B2 vssd1 vssd1 vccd1 vccd1 hold261/A
+ sky130_fd_sc_hd__a22o_1
X_11297_ _11398_/B _11397_/B hold294/A vssd1 vssd1 vccd1 vccd1 _11297_/X sky130_fd_sc_hd__a21o_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10317_ _11125_/A _10317_/B vssd1 vssd1 vccd1 vccd1 _10433_/D sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13036_ hold250/A _13035_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13036_/X sky130_fd_sc_hd__mux2_1
X_10248_ _10246_/X _10247_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _10248_/X sky130_fd_sc_hd__mux2_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07357__A1 _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07357__B2 _09295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10179_ fanout62/X fanout52/X _10677_/B fanout77/X vssd1 vssd1 vccd1 vccd1 _10180_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08306__B1 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07390_ _07139_/A _07139_/B _06864_/A vssd1 vssd1 vccd1 vccd1 _07393_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_57_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10196__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09060_ _09060_/A _09060_/B vssd1 vssd1 vccd1 vccd1 _11183_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_84_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08011_ _08011_/A _08011_/B vssd1 vssd1 vccd1 vccd1 _08013_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07001__C _07001_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09585__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09962_ _10229_/C _09962_/B vssd1 vssd1 vccd1 vccd1 _10002_/C sky130_fd_sc_hd__xnor2_2
X_08913_ _08912_/B _08912_/C _08912_/A vssd1 vssd1 vccd1 vccd1 _08914_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__09337__A2 _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12341__A1 _09198_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08545__B1 _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09893_ _07058_/A fanout18/X fanout9/X _08532_/B vssd1 vssd1 vccd1 vccd1 _09894_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07899__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08844_ _08844_/A _08844_/B vssd1 vssd1 vccd1 vccd1 _08845_/B sky130_fd_sc_hd__or2_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08775_ _08775_/A _08775_/B vssd1 vssd1 vccd1 vccd1 _08779_/A sky130_fd_sc_hd__xnor2_2
X_07726_ _07726_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07727_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07657_ _10169_/A _07657_/B vssd1 vssd1 vccd1 vccd1 _07661_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07520__B2 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07520__A1 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06608_ reg2_val[27] _06778_/B _06680_/B1 _06607_/Y vssd1 vssd1 vccd1 vccd1 _06837_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_48_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07588_ _07588_/A _07588_/B vssd1 vssd1 vccd1 vccd1 _07604_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06539_ instruction[5] vssd1 vssd1 vccd1 vccd1 _09200_/B sky130_fd_sc_hd__inv_6
XFILLER_0_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09273__A1 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09327_ _09327_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09328_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_63_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07284__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09273__B2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09258_ _09258_/A _09258_/B vssd1 vssd1 vccd1 vccd1 _09261_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_7_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08209_ _08209_/A _08209_/B vssd1 vssd1 vccd1 vccd1 _08630_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09189_ _11184_/A _12243_/B1 _08594_/B vssd1 vssd1 vccd1 vccd1 _09197_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08304__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07036__B1 _07034_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11220_ _12200_/A _11220_/B vssd1 vssd1 vccd1 vccd1 _11221_/B sky130_fd_sc_hd__xnor2_1
X_11151_ _11151_/A _11151_/B vssd1 vssd1 vccd1 vccd1 _11152_/B sky130_fd_sc_hd__nor2_1
XANTENNA__10553__B _10553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10102_ _10003_/X _10273_/B _10101_/Y vssd1 vssd1 vccd1 vccd1 _10102_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11082_ _06705_/A _11081_/X _12228_/B1 vssd1 vssd1 vccd1 vccd1 _11082_/Y sky130_fd_sc_hd__o21ai_1
X_10033_ _10033_/A _10033_/B vssd1 vssd1 vccd1 vccd1 _10075_/A sky130_fd_sc_hd__xnor2_1
X_11984_ reg1_val[24] curr_PC[24] vssd1 vssd1 vccd1 vccd1 _11984_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10935_ _11054_/A _10935_/B vssd1 vssd1 vccd1 vccd1 _10937_/B sky130_fd_sc_hd__or2_1
XFILLER_0_128_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10866_ _10750_/S _09831_/X _10865_/X _10752_/S vssd1 vssd1 vccd1 vccd1 _10866_/X
+ sky130_fd_sc_hd__o211a_1
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12605_ _12605_/A _12605_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[9] sky130_fd_sc_hd__xor2_4
XANTENNA__09264__A1 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13060__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10797_ _12022_/A _10797_/B vssd1 vssd1 vccd1 vccd1 _10801_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09264__B2 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12536_ _12539_/D _12536_/B vssd1 vssd1 vccd1 vccd1 new_PC[23] sky130_fd_sc_hd__xnor2_4
XANTENNA__07814__A2 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12467_ _12626_/B _12468_/B vssd1 vssd1 vccd1 vccd1 _12478_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11418_ _12019_/A _11418_/B vssd1 vssd1 vccd1 vccd1 _11422_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12398_ _12573_/B _12398_/B vssd1 vssd1 vccd1 vccd1 _12399_/B sky130_fd_sc_hd__or2_1
XFILLER_0_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11349_ _11349_/A _11349_/B vssd1 vssd1 vccd1 vccd1 _11350_/B sky130_fd_sc_hd__and2_1
XANTENNA__10582__B1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06890_ _06752_/A _06572_/X _09199_/B instruction[4] _06888_/Y vssd1 vssd1 vccd1
+ vccd1 _12722_/B sky130_fd_sc_hd__a221o_1
X_13019_ _06533_/Y _06537_/A rst vssd1 vssd1 vccd1 vccd1 _13019_/Y sky130_fd_sc_hd__a21oi_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10885__B2 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08560_ _08825_/A2 _09273_/A1 _09476_/A _08588_/B vssd1 vssd1 vccd1 vccd1 _08561_/B
+ sky130_fd_sc_hd__o22a_1
X_08491_ _08491_/A _08491_/B vssd1 vssd1 vccd1 vccd1 _08524_/A sky130_fd_sc_hd__xor2_2
XANTENNA__10919__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07511_ _07512_/A _07512_/B vssd1 vssd1 vccd1 vccd1 _09243_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_76_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout18 _12786_/A vssd1 vssd1 vccd1 vccd1 fanout18/X sky130_fd_sc_hd__clkbuf_8
Xfanout29 _07006_/Y vssd1 vssd1 vccd1 vccd1 fanout29/X sky130_fd_sc_hd__buf_6
XFILLER_0_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07442_ fanout69/X fanout98/X fanout56/X _11431_/A vssd1 vssd1 vccd1 vccd1 _07443_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10638__B _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07373_ _10557_/B _09295_/B _10433_/A fanout14/X vssd1 vssd1 vccd1 vccd1 _07374_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09112_ _09200_/A _09200_/B _09202_/A _06859_/Y vssd1 vssd1 vccd1 vccd1 _09218_/B
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_17_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07805__A2 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09043_ _09043_/A _09043_/B vssd1 vssd1 vccd1 vccd1 _10104_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_32_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11117__A2 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09945_ _09793_/A _09793_/B _09791_/Y vssd1 vssd1 vccd1 vccd1 _09947_/B sky130_fd_sc_hd__a21boi_4
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _09876_/A _09876_/B vssd1 vssd1 vccd1 vccd1 _09940_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__06579__A _06898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08827_ _08828_/B _08827_/B vssd1 vssd1 vccd1 vccd1 _08891_/B sky130_fd_sc_hd__and2b_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _10557_/A _08758_/A2 fanout58/X _07134_/A vssd1 vssd1 vccd1 vccd1 _08759_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _08689_/A _08689_/B _08689_/C vssd1 vssd1 vccd1 vccd1 _08701_/A sky130_fd_sc_hd__and3_1
X_07709_ _07308_/A _07308_/B _08819_/B2 vssd1 vssd1 vccd1 vccd1 _07710_/C sky130_fd_sc_hd__a21o_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10720_ _10720_/A _10720_/B vssd1 vssd1 vccd1 vccd1 _10722_/B sky130_fd_sc_hd__xnor2_2
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10651_ _10603_/A _10603_/B _10601_/Y vssd1 vssd1 vccd1 vccd1 _10728_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10582_ _12782_/A fanout95/X fanout54/X fanout22/X vssd1 vssd1 vccd1 vccd1 _10583_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12321_ _06585_/B _12274_/X _06583_/X vssd1 vssd1 vccd1 vccd1 _12321_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_51_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12252_ _07278_/B fanout8/X fanout7/X _12301_/A vssd1 vssd1 vccd1 vccd1 _12253_/B
+ sky130_fd_sc_hd__o22a_1
X_11203_ hold239/A _12332_/B _11302_/B _11920_/C1 vssd1 vssd1 vccd1 vccd1 _11203_/X
+ sky130_fd_sc_hd__a31o_1
X_12183_ hold264/A hold286/A _12183_/C vssd1 vssd1 vccd1 vccd1 _12240_/B sky130_fd_sc_hd__or3_1
XANTENNA__10564__B1 fanout12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ _11347_/A fanout15/X fanout6/X _11134_/B2 vssd1 vssd1 vccd1 vccd1 _11135_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10316__B1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065_ _11067_/A _11067_/B _11067_/C vssd1 vssd1 vccd1 vccd1 _11068_/A sky130_fd_sc_hd__a21oi_2
X_10016_ _10016_/A _10016_/B vssd1 vssd1 vccd1 vccd1 _10018_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06809__A_N _07303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11967_ _11967_/A _11967_/B vssd1 vssd1 vccd1 vccd1 _11969_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10918_ _12776_/A fanout47/X _11603_/A _11935_/A vssd1 vssd1 vccd1 vccd1 _10919_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11898_ _11898_/A _11898_/B vssd1 vssd1 vccd1 vccd1 _11972_/D sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10849_ _10730_/B _10959_/A vssd1 vssd1 vccd1 vccd1 _10850_/B sky130_fd_sc_hd__and2b_1
X_12519_ _12529_/A _12519_/B vssd1 vssd1 vccd1 vccd1 new_PC[20] sky130_fd_sc_hd__xnor2_4
XANTENNA__07799__A1 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07799__B2 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08748__B1 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07991_ fanout70/X _08774_/A2 _08774_/B1 _12762_/A vssd1 vssd1 vccd1 vccd1 _07992_/B
+ sky130_fd_sc_hd__o22a_2
Xfanout208 _07763_/A vssd1 vssd1 vccd1 vccd1 _08775_/A sky130_fd_sc_hd__clkbuf_16
Xfanout219 _06780_/X vssd1 vssd1 vccd1 vccd1 _09392_/S sky130_fd_sc_hd__buf_4
XFILLER_0_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06774__A2 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06942_ _07087_/B _07087_/C _07086_/C _07165_/A vssd1 vssd1 vccd1 vccd1 _06956_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_5_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09730_ _09597_/A _09597_/C _09597_/B vssd1 vssd1 vccd1 vccd1 _09731_/B sky130_fd_sc_hd__a21boi_4
XANTENNA__07723__A1 _07073_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07723__B2 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06873_ _09198_/C _12357_/A vssd1 vssd1 vccd1 vccd1 _06873_/Y sky130_fd_sc_hd__nand2_1
X_09661_ _09329_/X _09504_/X _09505_/X vssd1 vssd1 vccd1 vccd1 _09661_/X sky130_fd_sc_hd__a21o_1
X_08612_ _08485_/A _08485_/B _08485_/C vssd1 vssd1 vccd1 vccd1 _09009_/B sky130_fd_sc_hd__o21ai_1
X_09592_ _09592_/A _09592_/B vssd1 vssd1 vccd1 vccd1 _09593_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_82_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08543_ _07004_/A _07004_/B _06864_/A vssd1 vssd1 vccd1 vccd1 _08546_/B sky130_fd_sc_hd__a21o_1
XANTENNA_fanout161_A _07154_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout259_A _06898_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07487__B1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08474_ _08480_/A _08480_/B vssd1 vssd1 vccd1 vccd1 _08474_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07425_ _08982_/A _08982_/B _07422_/X vssd1 vssd1 vccd1 vccd1 _07622_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09228__A1 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09228__B2 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07356_ _07356_/A _07356_/B vssd1 vssd1 vccd1 vccd1 _07376_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07287_ _11125_/A _07287_/B vssd1 vssd1 vccd1 vccd1 _07355_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12583__B _12583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09026_ _08641_/A _08641_/B _08633_/A _08633_/B vssd1 vssd1 vccd1 vccd1 _09026_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__06581__B _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11991__C1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11338__A2 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold262 hold262/A vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__buf_1
Xhold251 hold251/A vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 hold240/A vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__buf_1
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold295 hold295/A vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 hold284/A vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
X_09928_ _09928_/A _09928_/B vssd1 vssd1 vccd1 vccd1 _09929_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout74_A _12768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _10273_/D _10273_/C _10002_/B _10617_/A vssd1 vssd1 vccd1 vccd1 _09859_/X
+ sky130_fd_sc_hd__a31o_1
X_12870_ _13121_/A _13122_/A _13121_/B vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_87_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11943__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06922__C1 _09199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ _11739_/A _11737_/X _11756_/A vssd1 vssd1 vccd1 vccd1 _11821_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_68_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10559__A _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ _12187_/A1 _11835_/B hold221/A vssd1 vssd1 vccd1 vccd1 _11754_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12774__A _12774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13015__A2 _06537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09219__A1 _12726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11683_ _12206_/A _11683_/B vssd1 vssd1 vccd1 vccd1 _11684_/A sky130_fd_sc_hd__xnor2_1
X_10703_ _10584_/A _10584_/B _10581_/A vssd1 vssd1 vccd1 vccd1 _10707_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_125_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10634_ hold205/A _12187_/A1 _10755_/B _10633_/Y _12290_/C1 vssd1 vssd1 vccd1 vccd1
+ _10641_/A sky130_fd_sc_hd__a311o_1
XANTENNA__12223__B1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11026__B2 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11026__A1 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11577__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12304_ _12786_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _12305_/B sky130_fd_sc_hd__nor2_1
X_10565_ _10565_/A _10565_/B vssd1 vssd1 vccd1 vccd1 _10567_/B sky130_fd_sc_hd__xnor2_1
X_13284_ _13311_/CLK _13284_/D vssd1 vssd1 vccd1 vccd1 hold246/A sky130_fd_sc_hd__dfxtp_1
X_10496_ _06739_/A _10371_/Y _06739_/B vssd1 vssd1 vccd1 vccd1 _10496_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_51_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12235_ _12361_/B _12235_/B vssd1 vssd1 vccd1 vccd1 _12235_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07402__B1 _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12166_ _11973_/B _12221_/A _12221_/B _11973_/A vssd1 vssd1 vccd1 vccd1 _12166_/X
+ sky130_fd_sc_hd__a31o_1
X_11117_ fanout33/X _11935_/A _12776_/A _10553_/A vssd1 vssd1 vccd1 vccd1 _11118_/B
+ sky130_fd_sc_hd__o22a_1
X_12097_ _12097_/A vssd1 vssd1 vccd1 vccd1 _12099_/A sky130_fd_sc_hd__inv_2
XANTENNA__07108__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11048_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11062_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11501__A2 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11853__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06947__A _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12999_ hold128/A _13013_/A2 _13020_/A2 hold107/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold108/A sky130_fd_sc_hd__o221a_1
XANTENNA__09458__A1 _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09458__B2 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08130__A1 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08130__B2 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13006__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08190_ _08190_/A _08190_/B vssd1 vssd1 vccd1 vccd1 _08247_/A sky130_fd_sc_hd__xor2_1
X_07210_ _07632_/A _07223_/B vssd1 vssd1 vccd1 vccd1 _07210_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_6_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12765__A1 _11511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07141_ _08595_/A _07141_/B vssd1 vssd1 vccd1 vccd1 _07160_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09630__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09630__B2 _10553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07072_ _10155_/A _07080_/C vssd1 vssd1 vccd1 vccd1 _07073_/B sky130_fd_sc_hd__and2_1
XFILLER_0_23_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07974_ _07974_/A _07974_/B vssd1 vssd1 vccd1 vccd1 _07977_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10370__C _10370_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06925_ _12487_/S _06925_/B vssd1 vssd1 vccd1 vccd1 dest_mask[0] sky130_fd_sc_hd__nand2_8
X_09713_ _12005_/A _09998_/C vssd1 vssd1 vccd1 vccd1 _09713_/Y sky130_fd_sc_hd__nor2_1
X_06856_ _06856_/A _06856_/B vssd1 vssd1 vccd1 vccd1 _06858_/A sky130_fd_sc_hd__nor2_1
X_09644_ _09496_/A _09496_/B _09494_/Y vssd1 vssd1 vccd1 vccd1 _09651_/A sky130_fd_sc_hd__a21o_1
XANTENNA__12578__B _12578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12048__A3 _09079_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06787_ _12563_/A _09679_/S vssd1 vssd1 vccd1 vccd1 _06787_/X sky130_fd_sc_hd__and2_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09575_ _09575_/A _09575_/B _09575_/C vssd1 vssd1 vccd1 vccd1 _09576_/B sky130_fd_sc_hd__and3_1
X_08526_ _09011_/A _09011_/B vssd1 vssd1 vccd1 vccd1 _09010_/B sky130_fd_sc_hd__nand2_1
X_08457_ _08457_/A _08457_/B _08457_/C vssd1 vssd1 vccd1 vccd1 _08457_/X sky130_fd_sc_hd__and3_1
XFILLER_0_77_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07408_ _08896_/A _08896_/B vssd1 vssd1 vccd1 vccd1 _08897_/A sky130_fd_sc_hd__or2_1
XANTENNA__11008__A1 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11008__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08388_ _08821_/A _08854_/B2 _08748_/B1 _08420_/B vssd1 vssd1 vccd1 vccd1 _08389_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_52_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08424__A2 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07339_ _07335_/A _07335_/B _07381_/A vssd1 vssd1 vccd1 vccd1 _07349_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_103_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10350_ _10216_/A _10216_/B _10214_/Y vssd1 vssd1 vccd1 vccd1 _10351_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_103_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09009_ _09009_/A _09009_/B vssd1 vssd1 vccd1 vccd1 _09009_/X sky130_fd_sc_hd__and2_1
XANTENNA__12533__S _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10281_ _10281_/A _10551_/B _10281_/C vssd1 vssd1 vccd1 vccd1 _10283_/A sky130_fd_sc_hd__and3_1
XFILLER_0_20_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08188__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08188__B2 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09408__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12020_ _12020_/A _12020_/B vssd1 vssd1 vccd1 vccd1 _12023_/A sky130_fd_sc_hd__nor2_1
X_12922_ _13116_/A hold181/X vssd1 vssd1 vccd1 vccd1 hold182/A sky130_fd_sc_hd__and2_1
XANTENNA__11673__A _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11495__A1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10298__A2 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12853_ hold9/X hold274/X vssd1 vssd1 vccd1 vccd1 _13082_/B sky130_fd_sc_hd__nand2b_1
X_12784_ _12784_/A _12786_/B vssd1 vssd1 vccd1 vccd1 _12784_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _11805_/A _11805_/B vssd1 vssd1 vccd1 vccd1 _11888_/B sky130_fd_sc_hd__or2_1
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _12332_/B _09069_/X _09073_/D _11184_/A _11734_/Y vssd1 vssd1 vccd1 vccd1
+ _11735_/X sky130_fd_sc_hd__a311o_1
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12747__A1 _10551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11666_ hold277/A _12119_/B1 _11748_/B _11665_/Y _11400_/A vssd1 vssd1 vccd1 vccd1
+ _11668_/C sky130_fd_sc_hd__a311o_1
XFILLER_0_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10617_ _10617_/A _10617_/B _10617_/C vssd1 vssd1 vccd1 vccd1 _10618_/B sky130_fd_sc_hd__or3_1
XFILLER_0_52_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11597_ _12022_/A _11597_/B vssd1 vssd1 vccd1 vccd1 _11598_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12009__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10548_ _10551_/B _10548_/B vssd1 vssd1 vccd1 vccd1 _10550_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_12_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13267_ _13277_/CLK _13267_/D vssd1 vssd1 vccd1 vccd1 hold116/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13172__B2 _06537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ _11968_/Y _12101_/X _12100_/Y vssd1 vssd1 vccd1 vccd1 _12218_/Y sky130_fd_sc_hd__a21oi_1
X_10479_ _10479_/A _10479_/B vssd1 vssd1 vccd1 vccd1 _10481_/B sky130_fd_sc_hd__xnor2_4
X_13198_ _13310_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_20_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12149_ _12087_/A _12088_/A _09252_/B vssd1 vssd1 vccd1 vccd1 _12151_/B sky130_fd_sc_hd__a21o_1
X_06710_ _06708_/Y _06710_/B vssd1 vssd1 vccd1 vccd1 _10972_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__10289__A2 _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07690_ _07690_/A _07690_/B vssd1 vssd1 vccd1 vccd1 _08969_/B sky130_fd_sc_hd__xor2_2
X_06641_ _06641_/A _12593_/B vssd1 vssd1 vccd1 vccd1 _06641_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06572_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06572_/X sky130_fd_sc_hd__or4bb_2
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09360_ _09207_/X _09359_/X _09679_/S vssd1 vssd1 vccd1 vccd1 _09360_/X sky130_fd_sc_hd__mux2_1
X_08311_ _08311_/A _08311_/B vssd1 vssd1 vccd1 vccd1 _08362_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09291_ _09291_/A _09291_/B vssd1 vssd1 vccd1 vccd1 _09292_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08242_ _08242_/A _08242_/B vssd1 vssd1 vccd1 vccd1 _08250_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_74_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10927__A _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_13 reg1_val[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_46 reg2_val[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 reg2_val[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_57 reg2_val[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07301__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 reg1_val[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08173_ _08857_/A _08173_/B vssd1 vssd1 vccd1 vccd1 _08243_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout124_A _07319_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_68 _10135_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 _12768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07124_ _12563_/A _07124_/B vssd1 vssd1 vccd1 vccd1 _08695_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11410__A1 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11410__B2 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07055_ _07111_/B _07055_/B vssd1 vssd1 vccd1 vccd1 _07055_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_684 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06601__A2_N _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ _08857_/A _07957_/B vssd1 vssd1 vccd1 vccd1 _07958_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07971__A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ instruction[19] _06552_/X _06907_/X _06678_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[1]
+ sky130_fd_sc_hd__o211a_4
X_07888_ _07888_/A _07888_/B vssd1 vssd1 vccd1 vccd1 _07939_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__06587__A _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06839_ reg1_val[25] _07157_/A vssd1 vssd1 vccd1 vccd1 _06839_/X sky130_fd_sc_hd__and2_1
X_09627_ _09628_/A _09628_/B vssd1 vssd1 vccd1 vccd1 _09629_/A sky130_fd_sc_hd__or2_1
X_09558_ _09402_/Y _09557_/X _12005_/A vssd1 vssd1 vccd1 vccd1 dest_val[2] sky130_fd_sc_hd__mux2_8
XANTENNA__09898__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08509_ _08509_/A _08509_/B vssd1 vssd1 vccd1 vccd1 _08527_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout37_A _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08645__A2 _08774_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11520_ _12019_/A _11520_/B vssd1 vssd1 vccd1 vccd1 _11522_/B sky130_fd_sc_hd__xnor2_1
X_09489_ _09489_/A _09489_/B vssd1 vssd1 vccd1 vccd1 _09502_/A sky130_fd_sc_hd__xor2_4
XANTENNA__12729__A1 _09283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10452__A2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11451_ _11451_/A _11451_/B vssd1 vssd1 vccd1 vccd1 _11453_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11382_ _06691_/Y _11287_/Y _06693_/B vssd1 vssd1 vccd1 vccd1 _11382_/X sky130_fd_sc_hd__a21o_1
X_10402_ _10523_/A _10523_/B _10523_/C vssd1 vssd1 vccd1 vccd1 _10524_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_33_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13121_ _13121_/A _13121_/B vssd1 vssd1 vccd1 vccd1 _13122_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_104_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07081__A1 _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10333_ _10333_/A _10333_/B vssd1 vssd1 vccd1 vccd1 _10334_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08042__A _08853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13052_ _13052_/A _13052_/B vssd1 vssd1 vccd1 vccd1 _13053_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_103_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10264_ reg1_val[7] curr_PC[7] vssd1 vssd1 vccd1 vccd1 _10265_/B sky130_fd_sc_hd__nand2_1
X_12003_ curr_PC[24] _12070_/C vssd1 vssd1 vccd1 vccd1 _12003_/X sky130_fd_sc_hd__or2_1
X_10195_ _10553_/A _12760_/A _11134_/B2 fanout33/X vssd1 vssd1 vccd1 vccd1 _10196_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13094__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12905_ hold189/X _12947_/A2 _12947_/B1 hold228/A vssd1 vssd1 vccd1 vccd1 hold190/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06928__C _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12836_ _13034_/A _13035_/A _13034_/B vssd1 vssd1 vccd1 vccd1 _13039_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__10691__A2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08097__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12968__A1 _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12767_ hold23/X _12778_/B _12766_/Y _13147_/A vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__o211a_1
XFILLER_0_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08217__A _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ _12698_/A _12698_/B _12698_/C vssd1 vssd1 vccd1 vccd1 _12700_/C sky130_fd_sc_hd__or3_1
XANTENNA__10443__A2 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11718_ _11719_/B _11719_/A vssd1 vssd1 vccd1 vccd1 _11809_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_126_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11649_ _06661_/C _11647_/X _11648_/Y vssd1 vssd1 vccd1 vccd1 _11668_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13319_ instruction[11] vssd1 vssd1 vccd1 vccd1 loadstore_dest[0] sky130_fd_sc_hd__buf_12
XFILLER_0_110_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08860_ _08860_/A _08860_/B vssd1 vssd1 vccd1 vccd1 _08861_/B sky130_fd_sc_hd__nand2_1
X_07811_ _08777_/A _07811_/B vssd1 vssd1 vccd1 vccd1 _07846_/B sky130_fd_sc_hd__xnor2_1
X_08791_ _08791_/A _08791_/B vssd1 vssd1 vccd1 vccd1 _08792_/B sky130_fd_sc_hd__xor2_2
X_07742_ _07821_/B _07821_/C _08544_/C vssd1 vssd1 vccd1 vccd1 _07744_/C sky130_fd_sc_hd__and3_1
XFILLER_0_74_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07673_ _10557_/A _08588_/B _09273_/A1 _07119_/Y vssd1 vssd1 vccd1 vccd1 _07674_/B
+ sky130_fd_sc_hd__o22a_1
X_06624_ _12713_/A _12370_/B vssd1 vssd1 vccd1 vccd1 _12357_/A sky130_fd_sc_hd__xnor2_4
X_09412_ _09412_/A _09412_/B vssd1 vssd1 vccd1 vccd1 _09413_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09511__A _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09343_ _09341_/X _09342_/X _09676_/S vssd1 vssd1 vccd1 vccd1 _09343_/X sky130_fd_sc_hd__mux2_1
X_06555_ instruction[20] _06915_/B vssd1 vssd1 vccd1 vccd1 _06555_/X sky130_fd_sc_hd__or2_1
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10657__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08127__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09274_ _09622_/A _09274_/B vssd1 vssd1 vccd1 vccd1 _09280_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_16_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08225_ _08692_/A2 fanout84/X fanout82/X _08692_/B1 vssd1 vssd1 vccd1 vccd1 _08226_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08156_ _08211_/A _08211_/B vssd1 vssd1 vccd1 vccd1 _08212_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07966__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11395__B1 _11838_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ _08589_/A _07115_/B vssd1 vssd1 vccd1 vccd1 _09764_/A sky130_fd_sc_hd__nand2_2
XANTENNA__07063__A1 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08087_ _08772_/B2 fanout82/X _08672_/B _08772_/A2 vssd1 vssd1 vccd1 vccd1 _08088_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07063__B2 _12768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07038_ _07105_/A _07038_/B vssd1 vssd1 vccd1 vccd1 _07039_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_30_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12895__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07366__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09392__S _09392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08989_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _09102_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11935__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08315__A1 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08315__B2 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__B1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ _10951_/A _10951_/B vssd1 vssd1 vccd1 vccd1 _10953_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10882_ _10863_/A _09383_/B _10878_/Y _10879_/X _10881_/X vssd1 vssd1 vccd1 vccd1
+ _10882_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12621_ _12629_/A _12621_/B vssd1 vssd1 vccd1 vccd1 _12623_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_109_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12552_ _12552_/A _12552_/B vssd1 vssd1 vccd1 vccd1 _12554_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_109_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08037__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07826__B1 _08692_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12782__A _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12483_ _12490_/A _12483_/B vssd1 vssd1 vccd1 vccd1 _12485_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11503_ _11504_/B _11503_/B vssd1 vssd1 vccd1 vccd1 _11618_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_124_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09579__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11434_ _11434_/A _11434_/B _11434_/C vssd1 vssd1 vccd1 vccd1 _11435_/B sky130_fd_sc_hd__or3_1
XANTENNA__13089__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10506__S _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11365_ _11365_/A _11365_/B vssd1 vssd1 vccd1 vccd1 _11367_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13104_ hold294/A _13103_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13104_/X sky130_fd_sc_hd__mux2_1
X_11296_ hold258/A _11296_/B vssd1 vssd1 vccd1 vccd1 _11397_/B sky130_fd_sc_hd__or2_1
XFILLER_0_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10316_ _10677_/A fanout95/X fanout54/X fanout58/X vssd1 vssd1 vccd1 vccd1 _10317_/B
+ sky130_fd_sc_hd__o22a_1
X_13035_ _13035_/A _13035_/B vssd1 vssd1 vccd1 vccd1 _13035_/Y sky130_fd_sc_hd__xnor2_1
X_10247_ _09673_/X _09678_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _10247_/X sky130_fd_sc_hd__mux2_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07357__A2 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10178_ _10894_/A _10178_/B vssd1 vssd1 vccd1 vccd1 _10182_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12022__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11861__A _11861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12819_ hold284/X hold77/X vssd1 vssd1 vccd1 vccd1 _13047_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08010_ _08011_/A _08011_/B vssd1 vssd1 vccd1 vccd1 _08010_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_72_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11377__B1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09961_ _09664_/B _09960_/X _09959_/Y vssd1 vssd1 vccd1 vccd1 _09962_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_100_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08912_ _08912_/A _08912_/B _08912_/C vssd1 vssd1 vccd1 vccd1 _08914_/B sky130_fd_sc_hd__or3_1
XFILLER_0_0_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _10030_/B _09892_/B vssd1 vssd1 vccd1 vccd1 _09917_/A sky130_fd_sc_hd__or2_1
XFILLER_0_85_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08843_ _08844_/A _08844_/B vssd1 vssd1 vccd1 vccd1 _08899_/B sky130_fd_sc_hd__nand2_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout289_A _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13028__A _13028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ _12768_/A _08774_/A2 _08774_/B1 _12766_/A vssd1 vssd1 vccd1 vccd1 _08775_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07725_ _07726_/B vssd1 vssd1 vccd1 vccd1 _07725_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_95_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06859__A1 _12713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ _08588_/A fanout36/X _08825_/A2 _08821_/B vssd1 vssd1 vccd1 vccd1 _07657_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07520__A2 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06607_ _06649_/A _12620_/B vssd1 vssd1 vccd1 vccd1 _06607_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06584__B _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ _07587_/A _07587_/B vssd1 vssd1 vccd1 vccd1 _07588_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_75_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06538_ instruction[3] vssd1 vssd1 vccd1 vccd1 _09198_/B sky130_fd_sc_hd__inv_2
XFILLER_0_48_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09326_ _09327_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09326_/X sky130_fd_sc_hd__and2_1
XFILLER_0_63_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09257_ _09256_/B _09256_/C _09256_/A vssd1 vssd1 vccd1 vccd1 _09258_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__07284__A1 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09273__A2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08208_ _08255_/A _08255_/B _08168_/Y vssd1 vssd1 vccd1 vccd1 _08630_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_106_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07284__B2 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09188_ _09200_/A _09200_/B _09188_/C vssd1 vssd1 vccd1 vccd1 _09188_/X sky130_fd_sc_hd__or3_4
XFILLER_0_16_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08139_ _08748_/B1 fanout55/X _12730_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08140_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08233__B1 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07036__A1 _07023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07036__B2 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09981__B1 _09198_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11011__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _11150_/A _11150_/B vssd1 vssd1 vccd1 vccd1 _11151_/B sky130_fd_sc_hd__and2_1
XFILLER_0_101_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10101_ _10003_/X _10273_/B _09110_/X vssd1 vssd1 vccd1 vccd1 _10101_/Y sky130_fd_sc_hd__a21oi_1
X_11081_ _06812_/Y _11080_/Y _11738_/S vssd1 vssd1 vccd1 vccd1 _11081_/X sky130_fd_sc_hd__mux2_1
X_10032_ _10033_/A _10033_/B vssd1 vssd1 vccd1 vccd1 _10212_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06759__B _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_4_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13305_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11983_ _11910_/B _11912_/B _11910_/A vssd1 vssd1 vccd1 vccd1 _11987_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11843__B2 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10934_ _10934_/A _10934_/B _10934_/C vssd1 vssd1 vccd1 vccd1 _10935_/B sky130_fd_sc_hd__and3_1
X_10865_ _11089_/A _10865_/B vssd1 vssd1 vccd1 vccd1 _10865_/X sky130_fd_sc_hd__or2_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12604_ _12609_/B _12611_/A vssd1 vssd1 vccd1 vccd1 _12605_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12535_ _12527_/B _12532_/B _12525_/X vssd1 vssd1 vccd1 vccd1 _12536_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10796_ fanout37/X _11431_/A _11347_/A fanout35/X vssd1 vssd1 vccd1 vccd1 _10797_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09264__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12466_ reg1_val[13] curr_PC[13] _12524_/S vssd1 vssd1 vccd1 vccd1 _12468_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_22_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11559__C _11559_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12397_ _12573_/B _12398_/B vssd1 vssd1 vccd1 vccd1 _12408_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11417_ fanout32/X _12150_/B _12776_/A fanout29/X vssd1 vssd1 vccd1 vccd1 _11418_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12017__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11348_ _11347_/A _12304_/B _11347_/C vssd1 vssd1 vccd1 vccd1 _11349_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__10582__A1 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10582__B2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11856__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11279_ _11279_/A _11279_/B vssd1 vssd1 vccd1 vccd1 _11279_/Y sky130_fd_sc_hd__nand2_1
X_13018_ _07277_/B _12744_/B hold49/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__a21oi_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07510_ _10180_/A _07510_/B vssd1 vssd1 vccd1 vccd1 _07512_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11591__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08490_ _08491_/A _08491_/B vssd1 vssd1 vccd1 vccd1 _08490_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07441_ _07441_/A _07441_/B vssd1 vssd1 vccd1 vccd1 _07464_/A sky130_fd_sc_hd__xnor2_4
Xfanout19 _12784_/A vssd1 vssd1 vccd1 vccd1 fanout19/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_119_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07372_ _07372_/A _07372_/B vssd1 vssd1 vccd1 vccd1 _07655_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09111_ _09559_/A _09108_/B _09108_/Y _12223_/B1 vssd1 vssd1 vccd1 vccd1 _09111_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08463__B1 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09042_ _09966_/B _09966_/C vssd1 vssd1 vccd1 vccd1 _10104_/B sky130_fd_sc_hd__and2_1
XFILLER_0_25_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08215__B1 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout204_A _08311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09963__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10022__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09944_ _09781_/A _09781_/B _09779_/Y vssd1 vssd1 vccd1 vccd1 _09947_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__08140__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09875_ _09875_/A _09875_/B vssd1 vssd1 vccd1 vccd1 _09876_/B sky130_fd_sc_hd__xnor2_4
X_08826_ _10306_/A _08826_/B vssd1 vssd1 vccd1 vccd1 _08827_/B sky130_fd_sc_hd__xnor2_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08757_ _09622_/A _08757_/B vssd1 vssd1 vccd1 vccd1 _08761_/A sky130_fd_sc_hd__xnor2_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _08678_/Y _08679_/X _08685_/X _08686_/Y vssd1 vssd1 vccd1 vccd1 _08689_/C
+ sky130_fd_sc_hd__a211o_1
X_07708_ _12734_/A _09752_/B vssd1 vssd1 vccd1 vccd1 _07710_/B sky130_fd_sc_hd__or2_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07639_ _09580_/A _07639_/B vssd1 vssd1 vccd1 vccd1 _08906_/B sky130_fd_sc_hd__xnor2_1
X_10650_ _11000_/A _10774_/A _12278_/A vssd1 vssd1 vccd1 vccd1 _10650_/X sky130_fd_sc_hd__o21a_1
X_09309_ _09309_/A _09309_/B vssd1 vssd1 vccd1 vccd1 _09310_/B sky130_fd_sc_hd__xor2_2
X_10581_ _10581_/A _10581_/B vssd1 vssd1 vccd1 vccd1 _10584_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_91_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12320_ _12319_/A _12319_/B _09110_/X vssd1 vssd1 vccd1 vccd1 _12320_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12002__A1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ _12249_/X _12250_/X _12345_/A vssd1 vssd1 vccd1 vccd1 dest_val[28] sky130_fd_sc_hd__a21oi_4
XFILLER_0_16_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11379__C _11379_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11202_ _12332_/B _11302_/B hold239/A vssd1 vssd1 vccd1 vccd1 _11202_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12182_ _12179_/Y _12180_/X _12181_/X _09851_/B vssd1 vssd1 vccd1 vccd1 _12182_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10564__B2 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10564__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11676__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11133_ _12255_/A _11133_/B vssd1 vssd1 vccd1 vccd1 _11142_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09706__B1 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10316__A1 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11064_ _11064_/A _11064_/B vssd1 vssd1 vccd1 vccd1 _11067_/C sky130_fd_sc_hd__xor2_1
XANTENNA__09182__A1 _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10316__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _10015_/A _10015_/B vssd1 vssd1 vccd1 vccd1 _10016_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11966_ _11808_/A _11890_/A _11889_/A vssd1 vssd1 vccd1 vccd1 _11966_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10917_ _10917_/A _10917_/B vssd1 vssd1 vccd1 vccd1 _10920_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_128_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11897_ _11179_/B _11552_/X _11893_/Y _11896_/X vssd1 vssd1 vccd1 vccd1 _11898_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_27_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10848_ _10959_/B _10959_/C vssd1 vssd1 vccd1 vccd1 _11070_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_54_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10779_ _12255_/A _10779_/B vssd1 vssd1 vccd1 vccd1 _10783_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12518_ _12519_/B vssd1 vssd1 vccd1 vccd1 _12518_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07799__A2 _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12449_ _12450_/A _12450_/B _12450_/C vssd1 vssd1 vccd1 vccd1 _12457_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_42_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08748__A1 _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__B2 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07990_ _09621_/A _07990_/B vssd1 vssd1 vccd1 vccd1 _07994_/A sky130_fd_sc_hd__xnor2_4
Xfanout209 _06918_/X vssd1 vssd1 vccd1 vccd1 _09205_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__06774__A3 _12573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06941_ reg1_val[24] reg1_val[25] vssd1 vssd1 vccd1 vccd1 _07086_/C sky130_fd_sc_hd__or2_2
XFILLER_0_5_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09660_ _09660_/A _09660_/B _09660_/C _09816_/A vssd1 vssd1 vccd1 vccd1 _10230_/B
+ sky130_fd_sc_hd__or4_2
XANTENNA__07723__A2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06872_ _06632_/X _06872_/B _06872_/C _06872_/D vssd1 vssd1 vccd1 vccd1 _06872_/X
+ sky130_fd_sc_hd__and4b_1
X_08611_ _09010_/B _09049_/A _09049_/B _08525_/Y _09052_/A vssd1 vssd1 vccd1 vccd1
+ _08611_/X sky130_fd_sc_hd__a311o_1
X_09591_ _09592_/A _09592_/B vssd1 vssd1 vccd1 vccd1 _09591_/Y sky130_fd_sc_hd__nand2_1
X_08542_ _08550_/B _08550_/A vssd1 vssd1 vccd1 vccd1 _08542_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_49_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08473_ _08473_/A _08473_/B vssd1 vssd1 vccd1 vccd1 _08480_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07487__A1 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08684__B1 _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07424_ _07424_/A _07424_/B vssd1 vssd1 vccd1 vccd1 _08982_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_15_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07487__B2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09228__A2 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07355_ _07355_/A _07355_/B vssd1 vssd1 vccd1 vccd1 _07356_/B sky130_fd_sc_hd__and2_1
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07286_ _07179_/Y fanout95/X _07553_/A fanout54/X vssd1 vssd1 vccd1 vccd1 _07287_/B
+ sky130_fd_sc_hd__o22a_1
X_09025_ _08163_/Y _08628_/X _08634_/X vssd1 vssd1 vccd1 vccd1 _09025_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07974__A _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold252 hold252/A vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold241 hold241/A vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold230 hold230/A vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold274 hold274/A vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold285 hold285/A vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 hold296/A vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
X_09927_ _09928_/A _09928_/B vssd1 vssd1 vccd1 vccd1 _09929_/A sky130_fd_sc_hd__and2_1
XANTENNA_fanout67_A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09858_ _10400_/S _09856_/Y _09857_/X _09855_/X vssd1 vssd1 vccd1 vccd1 dest_val[4]
+ sky130_fd_sc_hd__a31o_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08809_ _09032_/A _09077_/B vssd1 vssd1 vccd1 vccd1 _08933_/B sky130_fd_sc_hd__or2_1
X_09789_ _09913_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09792_/A sky130_fd_sc_hd__nor2_2
X_11820_ _11820_/A _11820_/B _11820_/C vssd1 vssd1 vccd1 vccd1 _11820_/X sky130_fd_sc_hd__and3_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ hold234/A _13236_/Q _11751_/C vssd1 vssd1 vccd1 vccd1 _11835_/B sky130_fd_sc_hd__or3_1
XANTENNA__06583__A_N _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08675__B1 _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10702_ _10832_/B _10702_/B vssd1 vssd1 vccd1 vccd1 _10708_/A sky130_fd_sc_hd__nand2_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09219__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11682_ _12205_/A _11935_/A _12776_/A _07389_/B vssd1 vssd1 vccd1 vccd1 _11683_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10633_ _12187_/A1 _10755_/B hold205/A vssd1 vssd1 vccd1 vccd1 _10633_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11026__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06772__B _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10564_ fanout77/X fanout46/X fanout12/X _11704_/A vssd1 vssd1 vccd1 vccd1 _10565_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12303_ fanout8/X _12301_/C _12302_/Y vssd1 vssd1 vccd1 vccd1 _12348_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13283_ _13311_/CLK _13283_/D vssd1 vssd1 vccd1 vccd1 hold250/A sky130_fd_sc_hd__dfxtp_1
X_10495_ _11973_/A _09048_/X _09050_/X _11381_/A vssd1 vssd1 vccd1 vccd1 _10495_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__11734__B1 _09073_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12234_ reg1_val[28] _12281_/C vssd1 vssd1 vccd1 vccd1 _12234_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07402__A1 _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12165_ _12215_/B _12165_/B vssd1 vssd1 vccd1 vccd1 _12221_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11116_ _11116_/A _11116_/B vssd1 vssd1 vccd1 vccd1 _11119_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12096_ _12098_/A _12098_/B _12098_/C vssd1 vssd1 vccd1 vccd1 _12097_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07108__B _07115_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11047_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11047_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_36_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06947__B _12370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12998_ _07317_/B _13020_/B2 hold129/X vssd1 vssd1 vccd1 vccd1 _13269_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_59_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07124__A _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09458__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08130__A2 _08672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11949_ _11950_/A _11950_/B vssd1 vssd1 vccd1 vccd1 _12025_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06963__A _11194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12765__A2 _12781_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07140_ _06864_/A _12782_/A _08758_/A2 fanout22/X vssd1 vssd1 vccd1 vccd1 _07141_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09630__A2 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07071_ _10155_/A _07080_/C vssd1 vssd1 vccd1 vccd1 _07073_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_100_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09933__A3 _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12205__A _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07973_ _12730_/A _07322_/A _07322_/B fanout47/X _08819_/B2 vssd1 vssd1 vccd1 vccd1
+ _07974_/B sky130_fd_sc_hd__o32a_1
X_09712_ curr_PC[3] _09712_/B vssd1 vssd1 vccd1 vccd1 _09998_/C sky130_fd_sc_hd__and2_1
X_06924_ instruction[24] _11823_/S is_load _06923_/X vssd1 vssd1 vccd1 vccd1 _06925_/B
+ sky130_fd_sc_hd__a31o_2
XANTENNA_fanout271_A _06537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06855_ _12276_/A _06854_/Y _06835_/Y vssd1 vssd1 vccd1 vccd1 _06856_/B sky130_fd_sc_hd__o21a_1
X_09643_ _09489_/A _09488_/B _09486_/Y vssd1 vssd1 vccd1 vccd1 _09653_/A sky130_fd_sc_hd__a21o_1
X_09574_ _09575_/A _09575_/B _09575_/C vssd1 vssd1 vccd1 vccd1 _09576_/A sky130_fd_sc_hd__a21oi_1
X_06786_ _06864_/A _09362_/S vssd1 vssd1 vccd1 vccd1 _09380_/B sky130_fd_sc_hd__nand2_1
X_08525_ _09011_/A _09011_/B vssd1 vssd1 vccd1 vccd1 _08525_/Y sky130_fd_sc_hd__nor2_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08456_ _08456_/A _08456_/B vssd1 vssd1 vccd1 vccd1 _08457_/C sky130_fd_sc_hd__xor2_1
XANTENNA__07969__A _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08387_ _08358_/A _08358_/B _08358_/C vssd1 vssd1 vccd1 vccd1 _08390_/B sky130_fd_sc_hd__o21ai_1
X_07407_ _10458_/A _07407_/B vssd1 vssd1 vccd1 vccd1 _08896_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11008__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07338_ _07380_/A _07380_/B vssd1 vssd1 vccd1 vccd1 _07381_/A sky130_fd_sc_hd__and2_1
XFILLER_0_45_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10767__B2 _06918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07269_ _11125_/A _07269_/B vssd1 vssd1 vccd1 vccd1 _07270_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_33_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09008_ _09008_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _09057_/A sky130_fd_sc_hd__xnor2_2
X_10280_ _10280_/A _10280_/B vssd1 vssd1 vccd1 vccd1 _10281_/C sky130_fd_sc_hd__xor2_1
XANTENNA__08188__A2 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12921_ hold215/A _12947_/A2 _12947_/B1 hold180/X vssd1 vssd1 vccd1 vccd1 hold181/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09424__A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12852_ _13077_/A _13078_/A _13077_/B vssd1 vssd1 vccd1 vccd1 _13083_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_68_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12783_ hold7/X _12786_/B _12782_/Y _13166_/A vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__o211a_1
XFILLER_0_95_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11247__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11803_ _11713_/A _11713_/B _11711_/X vssd1 vssd1 vccd1 vccd1 _11805_/B sky130_fd_sc_hd__a21oi_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11734_ _11559_/A _09069_/X _09073_/D vssd1 vssd1 vccd1 vccd1 _11734_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10455__B1 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11665_ _12119_/B1 _11748_/B hold277/A vssd1 vssd1 vccd1 vccd1 _11665_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12747__A2 _12980_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10616_ _10617_/A _10617_/B _10617_/C vssd1 vssd1 vccd1 vccd1 _10618_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11596_ fanout37/X _12150_/B _12776_/A fanout35/X vssd1 vssd1 vccd1 vccd1 _11597_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10547_ _07278_/B fanout83/X fanout81/X fanout7/X vssd1 vssd1 vccd1 vccd1 _10548_/B
+ sky130_fd_sc_hd__o22a_2
X_13266_ _13277_/CLK hold115/X vssd1 vssd1 vccd1 vccd1 hold113/A sky130_fd_sc_hd__dfxtp_1
X_10478_ _10479_/B _10479_/A vssd1 vssd1 vccd1 vccd1 _10478_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_121_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13172__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09376__A1 _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12217_ _12097_/A _12159_/A _12161_/B vssd1 vssd1 vccd1 vccd1 _12217_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_20_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13197_ _13296_/CLK _13197_/D vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12148_ _12148_/A _12148_/B vssd1 vssd1 vccd1 vccd1 _12154_/A sky130_fd_sc_hd__xor2_1
XANTENNA__06958__A _11780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12079_ _06965_/X _12349_/A _12078_/Y _10169_/A vssd1 vssd1 vccd1 vccd1 _12081_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11486__A2 _11838_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ instruction[32] _06678_/B vssd1 vssd1 vccd1 vccd1 _12593_/B sky130_fd_sc_hd__and2_4
XFILLER_0_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06571_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06898_/B sky130_fd_sc_hd__and4bb_1
XFILLER_0_87_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08310_ _07149_/Y _10551_/A _07325_/Y _07155_/X vssd1 vssd1 vccd1 vccd1 _08311_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09290_ _09291_/A _09291_/B vssd1 vssd1 vccd1 vccd1 _09290_/X sky130_fd_sc_hd__and2_1
XFILLER_0_117_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08241_ _08264_/A _08264_/B _08230_/Y vssd1 vssd1 vccd1 vccd1 _08250_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10927__B _12349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_14 reg1_val[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 reg2_val[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_47 reg2_val[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 reg1_val[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12199__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_69 instruction[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ _08748_/B1 _08217_/B fanout55/X _08821_/A vssd1 vssd1 vccd1 vccd1 _08173_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_58 reg2_val[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07301__B _11429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07123_ _12563_/A _07124_/B vssd1 vssd1 vccd1 vccd1 _09620_/A sky130_fd_sc_hd__xor2_4
XANTENNA__11410__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07054_ _07112_/B _07055_/B vssd1 vssd1 vccd1 vccd1 _11793_/A sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout117_A _07364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07029__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07956_ _08841_/A1 fanout55/X _08835_/B1 _08217_/B vssd1 vssd1 vccd1 vccd1 _07957_/B
+ sky130_fd_sc_hd__o22a_1
X_06907_ instruction[26] _06915_/B vssd1 vssd1 vccd1 vccd1 _06907_/X sky130_fd_sc_hd__or2_1
X_07887_ _07887_/A _07887_/B vssd1 vssd1 vccd1 vccd1 _08019_/A sky130_fd_sc_hd__xor2_4
XANTENNA__06587__B _12626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06838_ _06956_/A _07153_/A vssd1 vssd1 vccd1 vccd1 _06838_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07550__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09626_ _10578_/A _09626_/B vssd1 vssd1 vccd1 vccd1 _09628_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06769_ reg1_val[3] _11194_/S vssd1 vssd1 vccd1 vccd1 _06771_/B sky130_fd_sc_hd__nand2_1
X_09557_ _11381_/A _09515_/X _09556_/X _09513_/Y vssd1 vssd1 vccd1 vccd1 _09557_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_77_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08508_ _08509_/A _08509_/B vssd1 vssd1 vccd1 vccd1 _08508_/X sky130_fd_sc_hd__or2_1
XANTENNA__10437__B1 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09488_ _09486_/Y _09488_/B vssd1 vssd1 vccd1 vccd1 _09489_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07302__B1 _07303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08439_ _08841_/A1 _08758_/A2 _08835_/B1 _06864_/A vssd1 vssd1 vccd1 vccd1 _08440_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_38_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12729__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11450_ _11451_/A _11451_/B vssd1 vssd1 vccd1 vccd1 _11544_/B sky130_fd_sc_hd__and2_1
XFILLER_0_104_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11381_ _11381_/A _11381_/B _11381_/C vssd1 vssd1 vccd1 vccd1 _11381_/X sky130_fd_sc_hd__and3_2
X_10401_ curr_PC[9] _10646_/C vssd1 vssd1 vccd1 vccd1 _10401_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_116_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13120_ _13147_/A hold278/X vssd1 vssd1 vccd1 vccd1 _13301_/D sky130_fd_sc_hd__and2_1
XFILLER_0_33_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10332_ _10333_/A _10333_/B vssd1 vssd1 vccd1 vccd1 _10334_/A sky130_fd_sc_hd__and2_1
X_13051_ _13086_/A hold267/X vssd1 vssd1 vccd1 vccd1 _13287_/D sky130_fd_sc_hd__and2_1
X_10263_ reg1_val[7] curr_PC[7] vssd1 vssd1 vccd1 vccd1 _10263_/Y sky130_fd_sc_hd__nor2_1
X_12002_ _12223_/B1 _11974_/Y _11975_/X _11978_/X _12001_/X vssd1 vssd1 vccd1 vccd1
+ _12002_/X sky130_fd_sc_hd__a311o_1
XANTENNA__12901__A2 _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10194_ _10194_/A _10194_/B vssd1 vssd1 vccd1 vccd1 _10208_/A sky130_fd_sc_hd__nand2_1
X_12904_ _13169_/A hold225/X vssd1 vssd1 vccd1 vccd1 _13222_/D sky130_fd_sc_hd__and2_1
XANTENNA__10676__B1 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12835_ hold105/X hold250/X vssd1 vssd1 vccd1 vccd1 _13034_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08097__A1 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12968__A2 _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12766_ _12766_/A _12778_/B vssd1 vssd1 vccd1 vccd1 _12766_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08097__B2 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08217__B _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12697_ _12708_/B _12697_/B vssd1 vssd1 vccd1 vccd1 _12700_/B sky130_fd_sc_hd__nand2_1
X_11717_ _11622_/A _11622_/B _11623_/X vssd1 vssd1 vccd1 vccd1 _11719_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_126_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11648_ _06661_/C _11647_/X _12228_/B1 vssd1 vssd1 vccd1 vccd1 _11648_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11579_ _09115_/X _10867_/Y _10883_/Y _09184_/X _11578_/X vssd1 vssd1 vccd1 vccd1
+ _11579_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_52_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13318_ _13318_/CLK hold164/X vssd1 vssd1 vccd1 vccd1 hold163/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13249_ _13289_/CLK _13249_/D vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_110_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09048__B _10370_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07810_ _08477_/B fanout84/X fanout82/X _08776_/B1 vssd1 vssd1 vccd1 vccd1 _07811_/B
+ sky130_fd_sc_hd__o22a_1
X_08790_ _08791_/A _08791_/B vssd1 vssd1 vccd1 vccd1 _08790_/Y sky130_fd_sc_hd__nor2_1
X_07741_ _07062_/A _07062_/B _07134_/A vssd1 vssd1 vccd1 vccd1 _07744_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07672_ _07676_/A _07676_/B vssd1 vssd1 vccd1 vccd1 _07672_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09999__A _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10667__B1 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06623_ instruction[41] _06898_/A _06579_/B _06621_/X vssd1 vssd1 vccd1 vccd1 _12370_/B
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_90_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09411_ _09412_/A _09412_/B vssd1 vssd1 vccd1 vccd1 _09413_/A sky130_fd_sc_hd__or2_1
X_06554_ instruction[16] _06552_/X _06553_/X _06678_/B vssd1 vssd1 vccd1 vccd1 reg1_idx[5]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__12959__A2 _06537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09511__B _09511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09342_ _09120_/X _09123_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09342_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09285__B1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout234_A _09384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09273_ _09273_/A1 fanout18/X fanout9/X _08588_/B vssd1 vssd1 vccd1 vccd1 _09274_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ _08228_/A _08228_/B vssd1 vssd1 vccd1 vccd1 _08224_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_90_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08155_ _08155_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _08211_/B sky130_fd_sc_hd__and2_1
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07106_ reg1_val[4] _07106_/B vssd1 vssd1 vccd1 vccd1 _07115_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_43_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08086_ _08089_/A _08089_/B vssd1 vssd1 vccd1 vccd1 _08091_/A sky130_fd_sc_hd__or2_1
XANTENNA__08143__A _08853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07063__A2 _07055_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07037_ _10658_/A _07037_/B vssd1 vssd1 vccd1 vccd1 _07066_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07771__B1 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _08990_/B sky130_fd_sc_hd__nand2_1
X_07939_ _07939_/A _07939_/B vssd1 vssd1 vccd1 vccd1 _08021_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_98_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08315__A2 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__A _12349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10950_ _10951_/A _10951_/B vssd1 vssd1 vccd1 vccd1 _11067_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_98_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10881_ _06715_/B _09188_/X _09191_/X _06713_/Y _10880_/X vssd1 vssd1 vccd1 vccd1
+ _10881_/X sky130_fd_sc_hd__o221a_1
X_09609_ _07058_/A _07132_/Y fanout20/X _08532_/B vssd1 vssd1 vccd1 vccd1 _09610_/B
+ sky130_fd_sc_hd__o22a_1
X_12620_ reg1_val[12] _12620_/B vssd1 vssd1 vccd1 vccd1 _12621_/B sky130_fd_sc_hd__or2_1
XFILLER_0_93_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09276__B1 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12551_ _12551_/A _12551_/B vssd1 vssd1 vccd1 vccd1 _12552_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_109_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07826__A1 _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07826__B2 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12280__C1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12482_ _12637_/B _12482_/B vssd1 vssd1 vccd1 vccd1 _12483_/B sky130_fd_sc_hd__or2_1
XFILLER_0_93_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ _11604_/A _11502_/B vssd1 vssd1 vccd1 vccd1 _11503_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09579__A1 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09579__B2 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11433_ _11434_/A _11434_/B _11434_/C vssd1 vssd1 vccd1 vccd1 _11435_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10583__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11364_ _11364_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11367_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_235 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13103_ _13103_/A _13103_/B vssd1 vssd1 vccd1 vccd1 _13103_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11295_ _11208_/X _11294_/Y _11831_/S vssd1 vssd1 vccd1 vccd1 _11295_/X sky130_fd_sc_hd__mux2_1
X_10315_ _10894_/A _10315_/B vssd1 vssd1 vccd1 vccd1 _10433_/C sky130_fd_sc_hd__xnor2_1
X_13034_ _13034_/A _13034_/B vssd1 vssd1 vccd1 vccd1 _13035_/B sky130_fd_sc_hd__nand2_1
X_10246_ _09670_/X _09672_/X _10246_/S vssd1 vssd1 vccd1 vccd1 _10246_/X sky130_fd_sc_hd__mux2_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_4_4_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07762__B1 _08774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10177_ fanout22/X fanout98/X fanout56/X _10677_/A vssd1 vssd1 vccd1 vccd1 _10178_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12818_ hold266/X hold56/X vssd1 vssd1 vccd1 vccd1 _13052_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__07132__A _12250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09331__B _09331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12749_ _10694_/A _12980_/A2 hold82/X _13086_/A vssd1 vssd1 vccd1 vccd1 _13196_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09960_ _10229_/A _10229_/B vssd1 vssd1 vccd1 vccd1 _09960_/X sky130_fd_sc_hd__or2_1
XFILLER_0_110_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08911_ _08910_/B _08910_/C _08910_/A vssd1 vssd1 vccd1 vccd1 _08912_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10888__B1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _09891_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _09892_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_85_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08842_ _08842_/A _08842_/B vssd1 vssd1 vccd1 vccd1 _08844_/B sky130_fd_sc_hd__xnor2_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _08773_/A _08773_/B vssd1 vssd1 vccd1 vccd1 _08780_/A sky130_fd_sc_hd__xnor2_2
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07724_ _08777_/A _07724_/B vssd1 vssd1 vccd1 vccd1 _07726_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout184_A _08415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07655_ _07655_/A _07655_/B vssd1 vssd1 vccd1 vccd1 _07687_/A sky130_fd_sc_hd__xor2_1
XANTENNA__06859__A2 _12370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06606_ instruction[37] _06633_/B vssd1 vssd1 vccd1 vccd1 _12620_/B sky130_fd_sc_hd__and2_4
XFILLER_0_95_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10668__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08138__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07586_ _07587_/A _07587_/B vssd1 vssd1 vccd1 vccd1 _07586_/Y sky130_fd_sc_hd__nor2_1
X_06537_ _06537_/A vssd1 vssd1 vccd1 vccd1 _06537_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09325_ _09325_/A _09325_/B vssd1 vssd1 vccd1 vccd1 _09327_/B sky130_fd_sc_hd__xnor2_2
X_09256_ _09256_/A _09256_/B _09256_/C vssd1 vssd1 vccd1 vccd1 _09258_/A sky130_fd_sc_hd__and3_1
XANTENNA__07284__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08207_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08255_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_118_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11499__A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09187_ _09198_/C _09200_/B _09188_/C vssd1 vssd1 vccd1 vccd1 wire201/A sky130_fd_sc_hd__nor3_1
XFILLER_0_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08138_ _08855_/A _08138_/B vssd1 vssd1 vccd1 vccd1 _08144_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08233__B2 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08233__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07036__A2 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08069_ _08069_/A _08069_/B vssd1 vssd1 vccd1 vccd1 _08070_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_3_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11080_ _10972_/A _10970_/X _06710_/B vssd1 vssd1 vccd1 vccd1 _11080_/Y sky130_fd_sc_hd__o21ai_1
X_10100_ _10361_/A _10100_/B vssd1 vssd1 vccd1 vccd1 _10273_/B sky130_fd_sc_hd__xnor2_4
X_10031_ _10212_/A _10031_/B vssd1 vssd1 vccd1 vccd1 _10033_/B sky130_fd_sc_hd__and2_1
XANTENNA__07217__A _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11982_ _06604_/X _11980_/X _11981_/Y vssd1 vssd1 vccd1 vccd1 _11982_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_98_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06775__B _07279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10933_ _10934_/B _10934_/C _10934_/A vssd1 vssd1 vccd1 vccd1 _11054_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__10578__A _10578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08048__A _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13045__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ _10863_/A _10863_/B _10863_/Y _12277_/B1 vssd1 vssd1 vccd1 vccd1 _10864_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12603_ reg1_val[9] _12603_/B vssd1 vssd1 vccd1 vccd1 _12611_/A sky130_fd_sc_hd__nand2_1
X_10795_ _10795_/A _10795_/B vssd1 vssd1 vccd1 vccd1 _10807_/A sky130_fd_sc_hd__xnor2_1
X_12534_ _12551_/A _12534_/B vssd1 vssd1 vccd1 vccd1 _12539_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_109_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10803__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12465_ _12471_/B _12465_/B vssd1 vssd1 vccd1 vccd1 new_PC[12] sky130_fd_sc_hd__and2_4
XFILLER_0_41_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12396_ reg1_val[3] curr_PC[3] _12556_/S vssd1 vssd1 vccd1 vccd1 _12398_/B sky130_fd_sc_hd__mux2_1
X_11416_ _11416_/A _11416_/B vssd1 vssd1 vccd1 vccd1 _11439_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09972__A1 _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11347_ _11347_/A _12304_/B _11347_/C vssd1 vssd1 vccd1 vccd1 _11349_/A sky130_fd_sc_hd__or3_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10582__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08511__A _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ _11069_/Y _11279_/B _11276_/Y vssd1 vssd1 vccd1 vccd1 _11638_/A sky130_fd_sc_hd__a21bo_1
X_13017_ hold48/X _06537_/A _13151_/A2 _06533_/Y rst vssd1 vssd1 vccd1 vccd1 hold49/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__07735__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10229_ _10229_/A _10229_/B _10229_/C _10361_/A vssd1 vssd1 vccd1 vccd1 _10230_/C
+ sky130_fd_sc_hd__or4_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07440_ _07440_/A _07440_/B vssd1 vssd1 vccd1 vccd1 _07441_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07371_ _07371_/A _07371_/B vssd1 vssd1 vccd1 vccd1 _07372_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_29_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09110_ _09188_/C _09199_/B vssd1 vssd1 vccd1 vccd1 _09110_/X sky130_fd_sc_hd__or2_4
XFILLER_0_45_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08463__A1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08463__B2 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09041_ _09041_/A _09041_/B vssd1 vssd1 vccd1 vccd1 _09966_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_744 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08215__A1 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08215__B2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11112__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10022__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10022__B2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09943_ _09781_/A _09781_/B _09779_/Y vssd1 vssd1 vccd1 vccd1 _09946_/A sky130_fd_sc_hd__o21a_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ _09875_/A _09875_/B vssd1 vssd1 vccd1 vccd1 _09874_/Y sky130_fd_sc_hd__nand2b_1
X_08825_ fanout30/X _08825_/A2 _12730_/A _07000_/X vssd1 vssd1 vccd1 vccd1 _08826_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07037__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11782__A _11782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08756_ fanout62/X _08588_/B _09273_/A1 _11794_/A vssd1 vssd1 vccd1 vccd1 _08757_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12597__B _12598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11286__B1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08687_ _08685_/X _08686_/Y _08678_/Y _08679_/X vssd1 vssd1 vccd1 vccd1 _08689_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_68_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07707_ _07707_/A _07707_/B vssd1 vssd1 vccd1 vccd1 _09660_/A sky130_fd_sc_hd__xnor2_4
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13027__B2 _06537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07638_ _08841_/A1 fanout14/X _08835_/B1 _09752_/B vssd1 vssd1 vccd1 vccd1 _07639_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11038__B1 _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07569_ _10280_/A _07569_/B vssd1 vssd1 vccd1 vccd1 _07573_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_48_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09308_ _09309_/A _09309_/B vssd1 vssd1 vccd1 vccd1 _09308_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout12_A _07322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10580_ _10580_/A _10580_/B vssd1 vssd1 vccd1 vccd1 _10581_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07500__A _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10261__A1 _06866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09239_ _09239_/A _09239_/B vssd1 vssd1 vccd1 vccd1 _09241_/B sky130_fd_sc_hd__xor2_1
X_12250_ _12250_/A _12250_/B vssd1 vssd1 vccd1 vccd1 _12250_/X sky130_fd_sc_hd__or2_1
XFILLER_0_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11022__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11201_ hold180/A hold215/A _11201_/C vssd1 vssd1 vccd1 vccd1 _11302_/B sky130_fd_sc_hd__or3_1
X_12181_ _12361_/B _12181_/B vssd1 vssd1 vccd1 vccd1 _12181_/X sky130_fd_sc_hd__or2_1
XANTENNA__07965__B1 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11761__A1 _11733_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10564__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11132_ fanout70/X fanout27/X fanout26/X _11431_/A vssd1 vssd1 vccd1 vccd1 _11133_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10316__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11063_ _11064_/B _11064_/A vssd1 vssd1 vccd1 vccd1 _11171_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__07717__B1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ _09295_/A fanout57/X _11222_/A _09294_/A vssd1 vssd1 vccd1 vccd1 _10015_/B
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__06786__A _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08142__B1 _07181_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11965_ _12101_/A _12101_/B vssd1 vssd1 vccd1 vccd1 _12102_/A sky130_fd_sc_hd__nand2_2
XANTENNA__13018__A1 _07277_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10916_ _10916_/A _10916_/B vssd1 vssd1 vccd1 vccd1 _10917_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_67_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11029__B1 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ _11551_/X _11893_/Y _11894_/Y _11895_/Y vssd1 vssd1 vccd1 vccd1 _11896_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_128_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10847_ _10847_/A _10847_/B vssd1 vssd1 vccd1 vccd1 _10959_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10778_ fanout27/X _11134_/B2 fanout57/X _12205_/A vssd1 vssd1 vccd1 vccd1 _10779_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_27_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12517_ _12539_/A _12541_/A vssd1 vssd1 vccd1 vccd1 _12519_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_82_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12448_ _12457_/A _12448_/B vssd1 vssd1 vccd1 vccd1 _12450_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08748__A2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11867__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12379_ _12560_/B _12380_/B vssd1 vssd1 vccd1 vccd1 _12387_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06940_ reg1_val[23] _06940_/B _12658_/B vssd1 vssd1 vccd1 vccd1 _07087_/C sky130_fd_sc_hd__or3_4
X_06871_ _06871_/A _06871_/B _06871_/C vssd1 vssd1 vccd1 vccd1 _06872_/D sky130_fd_sc_hd__and3_1
XANTENNA__08381__B1 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ _09010_/B _09049_/A _09049_/B _08525_/Y vssd1 vssd1 vccd1 vccd1 _09052_/B
+ sky130_fd_sc_hd__a31o_1
X_09590_ _09482_/A _09482_/B _09480_/X vssd1 vssd1 vccd1 vccd1 _09592_/B sky130_fd_sc_hd__a21o_1
X_08541_ _08541_/A _08541_/B vssd1 vssd1 vccd1 vccd1 _08550_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_77_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08472_ _08470_/Y _08492_/B _08467_/Y vssd1 vssd1 vccd1 vccd1 _08480_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07487__A2 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07423_ _07423_/A _07423_/B vssd1 vssd1 vccd1 vccd1 _08982_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout147_A _06952_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07354_ _07354_/A _07354_/B vssd1 vssd1 vccd1 vccd1 _07426_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_17_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10243__A1 _06866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07285_ _10894_/A _07285_/B vssd1 vssd1 vccd1 vccd1 _07355_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09024_ _09022_/A _09022_/B _09023_/Y _08641_/Y _08633_/Y vssd1 vssd1 vccd1 vccd1
+ _09028_/A sky130_fd_sc_hd__a2111o_2
XFILLER_0_115_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold220 hold220/A vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold287/A vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10681__A _11695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 hold264/A vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 hold286/A vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 hold297/A vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ _09926_/A _09926_/B vssd1 vssd1 vccd1 vccd1 _09928_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07990__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09857_ curr_PC[4] _09998_/C vssd1 vssd1 vccd1 vccd1 _09857_/X sky130_fd_sc_hd__or2_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10620__S _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08808_ _08806_/X _09029_/B vssd1 vssd1 vccd1 vccd1 _09077_/B sky130_fd_sc_hd__nand2b_2
X_09788_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__nor2_1
X_08739_ _08739_/A _08739_/B vssd1 vssd1 vccd1 vccd1 _08741_/B sky130_fd_sc_hd__xnor2_1
X_11750_ hold252/A _12119_/B1 _11832_/B _11400_/A vssd1 vssd1 vccd1 vccd1 _11750_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08124__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10701_ _10832_/A _10699_/C _10699_/A vssd1 vssd1 vccd1 vccd1 _10702_/B sky130_fd_sc_hd__a21o_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10880__A1_N _07303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11681_ _11777_/A _11681_/B vssd1 vssd1 vccd1 vccd1 _11686_/A sky130_fd_sc_hd__and2_1
XFILLER_0_119_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08326__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10632_ hold198/A _10632_/B vssd1 vssd1 vccd1 vccd1 _10755_/B sky130_fd_sc_hd__or2_1
XFILLER_0_64_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10563_ _10705_/B _10563_/B vssd1 vssd1 vccd1 vccd1 _10567_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12302_ _12206_/A _07277_/B fanout8/X _12349_/B vssd1 vssd1 vccd1 vccd1 _12302_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_24_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13282_ _13311_/CLK _13282_/D vssd1 vssd1 vccd1 vccd1 hold279/A sky130_fd_sc_hd__dfxtp_1
X_10494_ _11973_/A _09048_/X _09050_/X vssd1 vssd1 vccd1 vccd1 _10494_/Y sky130_fd_sc_hd__o21ai_1
X_12233_ _12179_/A _12176_/Y _12178_/B vssd1 vssd1 vccd1 vccd1 _12281_/C sky130_fd_sc_hd__o21ai_2
XFILLER_0_32_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07402__A2 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12164_ _12040_/B _12163_/Y _12162_/X vssd1 vssd1 vccd1 vccd1 _12165_/B sky130_fd_sc_hd__o21ai_1
X_12095_ _12160_/B _12095_/B vssd1 vssd1 vccd1 vccd1 _12098_/C sky130_fd_sc_hd__nand2_1
X_11115_ _11116_/A _11116_/B vssd1 vssd1 vccd1 vccd1 _11115_/X sky130_fd_sc_hd__and2_1
X_11046_ _11046_/A _11046_/B vssd1 vssd1 vccd1 vccd1 _11048_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07405__A _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12997_ hold110/X _13013_/A2 _13020_/A2 hold128/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold129/A sky130_fd_sc_hd__o221a_1
XANTENNA__09620__A _09620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ _12025_/A _11948_/B vssd1 vssd1 vccd1 vccd1 _11950_/B sky130_fd_sc_hd__and2_1
X_11879_ _11932_/A _11879_/B vssd1 vssd1 vccd1 vccd1 _11881_/B sky130_fd_sc_hd__or2_1
XFILLER_0_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07070_ reg1_val[8] _07070_/B vssd1 vssd1 vccd1 vccd1 _07080_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_54_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11597__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12205__B fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07972_ _07971_/B _07971_/C _09580_/A vssd1 vssd1 vccd1 vccd1 _07977_/B sky130_fd_sc_hd__a21o_1
X_09711_ curr_PC[3] _09712_/B vssd1 vssd1 vccd1 vccd1 _09711_/X sky130_fd_sc_hd__or2_1
X_06923_ _06923_/A _06923_/B _06923_/C vssd1 vssd1 vccd1 vccd1 _06923_/X sky130_fd_sc_hd__and3_1
XANTENNA__08354__B1 _08695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06854_ _06592_/Y _12225_/B _06845_/A vssd1 vssd1 vccd1 vccd1 _06854_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09514__B _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09642_ _09642_/A _09642_/B vssd1 vssd1 vccd1 vccd1 _09655_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_117_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06785_ reg2_val[0] _06778_/B _06649_/A _06783_/X vssd1 vssd1 vccd1 vccd1 _06785_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07315__A _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09573_ _09573_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09575_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08524_ _08524_/A _08524_/B vssd1 vssd1 vccd1 vccd1 _09011_/B sky130_fd_sc_hd__xor2_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07969__B _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08455_ _08484_/A _08484_/B vssd1 vssd1 vccd1 vccd1 _08457_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08386_ _08399_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08401_/A sky130_fd_sc_hd__and2b_1
X_07406_ _10156_/B2 fanout69/X _10156_/A1 _12762_/A vssd1 vssd1 vccd1 vccd1 _07407_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_46_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07337_ _10306_/A _07337_/B vssd1 vssd1 vccd1 vccd1 _07380_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07268_ _11134_/B2 fanout95/X fanout54/X fanout57/X vssd1 vssd1 vccd1 vccd1 _07269_/B
+ sky130_fd_sc_hd__o22a_1
X_09007_ _08621_/A _09007_/B vssd1 vssd1 vccd1 vccd1 _09007_/X sky130_fd_sc_hd__and2b_1
X_07199_ _08857_/A _07199_/B vssd1 vssd1 vccd1 vccd1 _07631_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08593__B1 _08544_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ _09909_/A _09909_/B _09909_/C vssd1 vssd1 vccd1 vccd1 _10037_/A sky130_fd_sc_hd__nand3_1
XANTENNA_clkbuf_4_9_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12920_ _12946_/A hold216/X vssd1 vssd1 vccd1 vccd1 _13230_/D sky130_fd_sc_hd__and2_1
XFILLER_0_88_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12131__A _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__B1 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12851_ hold61/X hold291/X vssd1 vssd1 vccd1 vccd1 _13077_/B sky130_fd_sc_hd__nand2b_1
X_11802_ _11802_/A _11802_/B vssd1 vssd1 vccd1 vccd1 _11805_/A sky130_fd_sc_hd__xnor2_1
X_12782_ _12782_/A _12786_/B vssd1 vssd1 vccd1 vccd1 _12782_/Y sky130_fd_sc_hd__nand2_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09845__B1 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06783__B _12563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07320__A1 _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ _11767_/B _11731_/Y _11732_/Y vssd1 vssd1 vccd1 vccd1 _11733_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_37_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10455__A1 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10455__B2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11664_ hold280/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11748_/B sky130_fd_sc_hd__or2_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10615_ _12278_/A _11000_/A _10774_/A _09110_/X vssd1 vssd1 vccd1 vccd1 _10615_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11595_ _11595_/A _11595_/B vssd1 vssd1 vccd1 vccd1 _11599_/B sky130_fd_sc_hd__xor2_1
X_10546_ _10454_/Y _10459_/B _10457_/X vssd1 vssd1 vccd1 vccd1 _10550_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_121_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13265_ _13277_/CLK hold44/X vssd1 vssd1 vccd1 vccd1 _13265_/Q sky130_fd_sc_hd__dfxtp_1
X_10477_ _10477_/A _10477_/B vssd1 vssd1 vccd1 vccd1 _10479_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12216_ _12216_/A _12216_/B _12216_/C _12313_/A vssd1 vssd1 vccd1 vccd1 _12216_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_20_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13196_ _13296_/CLK _13196_/D vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfxtp_1
X_12147_ _12206_/A _12147_/B vssd1 vssd1 vccd1 vccd1 _12148_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12078_ _12078_/A _12349_/A vssd1 vssd1 vccd1 vccd1 _12078_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06958__B _06965_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11029_ fanout32/X _11794_/A _11704_/A fanout29/X vssd1 vssd1 vccd1 vccd1 _11030_/B
+ sky130_fd_sc_hd__o22a_1
X_06570_ instruction[0] instruction[1] instruction[2] instruction[41] pred_val vssd1
+ vssd1 vccd1 vccd1 _12658_/A sky130_fd_sc_hd__o311a_4
XANTENNA__09836__B1 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08240_ _08240_/A _08240_/B vssd1 vssd1 vccd1 vccd1 _08264_/B sky130_fd_sc_hd__xor2_2
X_08171_ _08733_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _08243_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_48 reg2_val[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_37 reg2_val[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09203__A2_N _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_26 reg1_val[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_15 reg1_val[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12199__A1 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12199__B2 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_59 reg2_val[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07122_ reg1_val[0] reg1_val[31] _09968_/A vssd1 vssd1 vccd1 vccd1 _07124_/B sky130_fd_sc_hd__and3_4
XFILLER_0_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07053_ _07128_/B _07111_/C _07135_/B vssd1 vssd1 vccd1 vccd1 _07055_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10382__B1 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ _07955_/A _07955_/B vssd1 vssd1 vccd1 vccd1 _07958_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06906_ instruction[18] _06552_/X _06905_/X _06678_/B vssd1 vssd1 vccd1 vccd1 reg2_idx[0]
+ sky130_fd_sc_hd__o211a_4
XANTENNA__09093__B1_N _12230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ _07887_/A _07887_/B vssd1 vssd1 vccd1 vccd1 _07886_/X sky130_fd_sc_hd__and2_1
XANTENNA__06889__B1 _09199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07045__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09625_ fanout69/X _08134_/B fanout51/X _12762_/A vssd1 vssd1 vccd1 vccd1 _09626_/B
+ sky130_fd_sc_hd__o22a_1
X_06837_ reg1_val[27] _06837_/B vssd1 vssd1 vccd1 vccd1 _06837_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07550__B2 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07550__A1 _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06768_ reg1_val[3] _11194_/S vssd1 vssd1 vccd1 vccd1 _06768_/Y sky130_fd_sc_hd__nor2_1
X_09556_ _06919_/X _09551_/X _09552_/X _09555_/Y vssd1 vssd1 vccd1 vccd1 _09556_/X
+ sky130_fd_sc_hd__a211o_1
X_06699_ reg2_val[14] _06729_/B vssd1 vssd1 vccd1 vccd1 _06699_/X sky130_fd_sc_hd__and2_1
XFILLER_0_78_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08507_ _08529_/A _08507_/B vssd1 vssd1 vccd1 vccd1 _08509_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09260__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10437__A1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10437__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09487_ _09487_/A _09487_/B vssd1 vssd1 vccd1 vccd1 _09488_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08438_ _09898_/A _08438_/B vssd1 vssd1 vccd1 vccd1 _08445_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_65_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08369_ _08367_/A _08367_/B _08368_/X vssd1 vssd1 vccd1 vccd1 _08619_/B sky130_fd_sc_hd__o21bai_4
XANTENNA__11014__B _11014_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11380_ _11379_/A _11379_/B _11379_/C vssd1 vssd1 vccd1 vccd1 _11381_/C sky130_fd_sc_hd__o21ai_1
X_10400_ _10396_/X _10399_/Y _10400_/S vssd1 vssd1 vccd1 vccd1 dest_val[8] sky130_fd_sc_hd__mux2_8
XFILLER_0_104_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10331_ _11604_/A _10331_/B vssd1 vssd1 vccd1 vccd1 _10333_/B sky130_fd_sc_hd__xnor2_1
X_13050_ hold266/X _12721_/B _13049_/X _12722_/A vssd1 vssd1 vccd1 vccd1 hold267/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10262_ _10132_/A _10129_/Y _10131_/B vssd1 vssd1 vccd1 vccd1 _10266_/A sky130_fd_sc_hd__o21a_1
XANTENNA__11030__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12001_ _09851_/B _11988_/X _12000_/X _11982_/X vssd1 vssd1 vccd1 vccd1 _12001_/X
+ sky130_fd_sc_hd__a211o_1
X_10193_ _10193_/A _10193_/B vssd1 vssd1 vccd1 vccd1 _10209_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08318__B1 _07182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06778__B _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12903_ hold224/X _12947_/A2 _12947_/B1 hold189/X vssd1 vssd1 vccd1 vccd1 hold225/A
+ sky130_fd_sc_hd__a22o_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12834_ _13029_/A _13030_/A _13029_/B vssd1 vssd1 vccd1 vccd1 _13035_/A sky130_fd_sc_hd__a21bo_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ _11511_/A _12781_/A2 hold89/X _13116_/A vssd1 vssd1 vccd1 vccd1 _13204_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08097__A2 _08348_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13090__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11716_ _11809_/A _11716_/B vssd1 vssd1 vccd1 vccd1 _11719_/A sky130_fd_sc_hd__and2_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12705_/A _12696_/B vssd1 vssd1 vccd1 vccd1 _12700_/A sky130_fd_sc_hd__or2_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11647_ _06824_/X _11646_/X _11647_/S vssd1 vssd1 vccd1 vccd1 _11647_/X sky130_fd_sc_hd__mux2_1
X_11578_ _06666_/Y _12243_/B1 _11576_/X _06668_/B _11577_/X vssd1 vssd1 vccd1 vccd1
+ _11578_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_64_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06596__A_N _07157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13317_ _13318_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09329__B _09331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10529_ _10445_/A _10445_/B _10441_/X vssd1 vssd1 vccd1 vccd1 _10531_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_24_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13248_ _13248_/CLK hold151/X vssd1 vssd1 vccd1 vccd1 hold149/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08557__B1 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13179_ _13179_/A _13179_/B hold155/X vssd1 vssd1 vccd1 vccd1 hold156/A sky130_fd_sc_hd__and3_1
X_07740_ _08821_/A _10553_/A vssd1 vssd1 vccd1 vccd1 _08004_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_74_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07671_ _08595_/A _07671_/B vssd1 vssd1 vccd1 vccd1 _07676_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10667__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10667__A1 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06622_ _06541_/Y _06688_/B1 _06621_/X vssd1 vssd1 vccd1 vccd1 _06622_/X sky130_fd_sc_hd__o21ba_2
X_09410_ _10306_/A _09410_/B vssd1 vssd1 vccd1 vccd1 _09412_/B sky130_fd_sc_hd__xor2_1
X_06553_ instruction[23] _06915_/B vssd1 vssd1 vccd1 vccd1 _06553_/X sky130_fd_sc_hd__or2_1
XFILLER_0_87_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09341_ _09116_/X _09119_/X _09359_/S vssd1 vssd1 vccd1 vccd1 _09341_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09285__A1 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09285__B2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09272_ _09438_/B _09272_/B vssd1 vssd1 vccd1 vccd1 _09281_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08223_ _09621_/A _08223_/B vssd1 vssd1 vccd1 vccd1 _08228_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08154_ _08154_/A _08154_/B vssd1 vssd1 vccd1 vccd1 _08155_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout227_A _07001_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12041__B1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08085_ _08777_/A _08085_/B vssd1 vssd1 vccd1 vccd1 _08089_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11395__A2 wire201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07105_ _07105_/A _07105_/B vssd1 vssd1 vccd1 vccd1 _07106_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_101_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07036_ _07023_/Y _10452_/B2 _07034_/Y _10527_/A vssd1 vssd1 vccd1 vccd1 _07037_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_113_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11785__A _11861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12895__A2 _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09255__A _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__A1 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07771__B2 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _08990_/A sky130_fd_sc_hd__or2_1
XANTENNA__06598__B _07157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07938_ _07937_/A _08068_/A vssd1 vssd1 vccd1 vccd1 _08021_/A sky130_fd_sc_hd__and2b_1
X_07869_ _12762_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07871_/C sky130_fd_sc_hd__or2_1
XANTENNA__11855__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10880_ _07303_/A _06928_/X _11099_/B reg1_val[12] vssd1 vssd1 vccd1 vccd1 _10880_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_09608_ _10658_/A _09608_/B vssd1 vssd1 vccd1 vccd1 _09612_/A sky130_fd_sc_hd__xnor2_1
X_09539_ _11197_/S _09539_/B vssd1 vssd1 vccd1 vccd1 _09539_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout42_A _11147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09276__A1 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09276__B2 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12550_ _12551_/A _12551_/B vssd1 vssd1 vccd1 vccd1 _12552_/A sky130_fd_sc_hd__and2_1
XANTENNA__07826__A2 _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12481_ _12637_/B _12482_/B vssd1 vssd1 vccd1 vccd1 _12490_/A sky130_fd_sc_hd__nand2_1
X_11501_ _12301_/A _11603_/A fanout8/X fanout47/X vssd1 vssd1 vccd1 vccd1 _11502_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_19_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09579__A2 _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11432_ _11509_/A _11432_/B vssd1 vssd1 vccd1 vccd1 _11434_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_123_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13102_ _13102_/A _13102_/B vssd1 vssd1 vccd1 vccd1 _13103_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_104_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11363_ _11364_/A _11364_/B vssd1 vssd1 vccd1 vccd1 _11457_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11294_ _11294_/A _11294_/B vssd1 vssd1 vccd1 vccd1 _11294_/Y sky130_fd_sc_hd__xnor2_1
X_10314_ _12782_/A fanout98/X fanout56/X fanout22/X vssd1 vssd1 vccd1 vccd1 _10315_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_21_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13033_ _13086_/A hold251/X vssd1 vssd1 vccd1 vccd1 _13283_/D sky130_fd_sc_hd__and2_1
X_10245_ _10251_/S _10244_/X _09214_/A vssd1 vssd1 vccd1 vccd1 _10245_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11695__A _11695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07211__B1 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ _10013_/B _10016_/B _10013_/A vssd1 vssd1 vccd1 vccd1 _10190_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__07762__A1 _07023_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07762__B2 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 _06946_/X vssd1 vssd1 vccd1 vccd1 _07303_/B sky130_fd_sc_hd__buf_6
XFILLER_0_88_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10649__A1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12817_ hold292/A hold73/X vssd1 vssd1 vccd1 vccd1 _13057_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_97_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12748_ hold81/X _12788_/B vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__or2_1
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11074__A1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10821__A1 _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12679_ _12660_/B _12678_/X _12714_/A _07087_/C vssd1 vssd1 vccd1 vccd1 _12681_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_115_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09059__B _09059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08910_ _08910_/A _08910_/B _08910_/C vssd1 vssd1 vccd1 vccd1 _08912_/B sky130_fd_sc_hd__and3_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09890_ _09891_/A _09891_/B vssd1 vssd1 vccd1 vccd1 _10030_/B sky130_fd_sc_hd__and2_1
X_08841_ _08841_/A1 _07301_/Y fanout14/X _08841_/B2 vssd1 vssd1 vccd1 vccd1 _08842_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _07023_/Y _08772_/A2 fanout69/X _08772_/B2 vssd1 vssd1 vccd1 vccd1 _08773_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06961__C1 _12370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07307__B _11429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07723_ _07073_/X fanout94/X _12752_/A _10156_/A1 vssd1 vssd1 vccd1 vccd1 _07724_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_fanout177_A _12781_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11301__A2 _11838_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07654_ _07690_/A _07690_/B vssd1 vssd1 vccd1 vccd1 _07654_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06605_ _12276_/A _06605_/B _12045_/A _06604_/X vssd1 vssd1 vccd1 vccd1 _06632_/A
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_125_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07585_ _07585_/A _07585_/B vssd1 vssd1 vccd1 vccd1 _07587_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06536_ hold40/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__inv_2
XFILLER_0_48_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09324_ _09325_/B _09325_/A vssd1 vssd1 vccd1 vccd1 _09324_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_62_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09255_ _09610_/A _09255_/B _09255_/C vssd1 vssd1 vccd1 vccd1 _09256_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_35_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08206_ _08213_/A _08213_/B _08197_/X vssd1 vssd1 vccd1 vccd1 _08255_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_90_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09186_ _09202_/A _09199_/B vssd1 vssd1 vccd1 vccd1 _11184_/A sky130_fd_sc_hd__or2_4
X_08137_ _08837_/B2 _08420_/B _08854_/B2 _07969_/A vssd1 vssd1 vccd1 vccd1 _08138_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08233__A2 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08068_ _08068_/A _08068_/B vssd1 vssd1 vccd1 vccd1 _08070_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_101_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07019_ _07178_/A _07192_/A _07197_/A _07303_/A vssd1 vssd1 vccd1 vccd1 _07021_/B
+ sky130_fd_sc_hd__or4_1
XANTENNA__12404__A _12578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10328__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10030_ _10030_/A _10030_/B _10030_/C vssd1 vssd1 vccd1 vccd1 _10031_/B sky130_fd_sc_hd__or3_1
XANTENNA__10541__A1_N fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _06604_/X _11980_/X _12277_/B1 vssd1 vssd1 vccd1 vccd1 _11981_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09713__A _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10932_ _10805_/A _10805_/B _10802_/A vssd1 vssd1 vccd1 vccd1 _10937_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13045__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10863_ _10863_/A _10863_/B vssd1 vssd1 vccd1 vccd1 _10863_/Y sky130_fd_sc_hd__nor2_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12602_ reg1_val[9] _12603_/B vssd1 vssd1 vccd1 vccd1 _12609_/B sky130_fd_sc_hd__or2_1
X_10794_ _10795_/A _10795_/B vssd1 vssd1 vccd1 vccd1 _10943_/A sky130_fd_sc_hd__and2_1
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12533_ reg1_val[23] curr_PC[23] _12556_/S vssd1 vssd1 vccd1 vccd1 _12534_/B sky130_fd_sc_hd__mux2_4
XFILLER_0_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10803__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10803__A1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06791__B _06964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12464_ _12464_/A _12464_/B _12464_/C vssd1 vssd1 vccd1 vccd1 _12465_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12395_ _12401_/B _12395_/B vssd1 vssd1 vccd1 vccd1 new_PC[2] sky130_fd_sc_hd__and2_4
XFILLER_0_61_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11415_ _11416_/A _11416_/B vssd1 vssd1 vccd1 vccd1 _11415_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07432__B1 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11346_ _12206_/A _11346_/B vssd1 vssd1 vccd1 vccd1 _11347_/C sky130_fd_sc_hd__xnor2_1
X_13016_ _07090_/X _12744_/B hold53/X vssd1 vssd1 vccd1 vccd1 _13278_/D sky130_fd_sc_hd__a21oi_1
X_11277_ _11462_/A _11462_/B vssd1 vssd1 vccd1 vccd1 _11279_/B sky130_fd_sc_hd__nor2_1
XANTENNA__07735__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ _10229_/C _10361_/A vssd1 vssd1 vccd1 vccd1 _10487_/A sky130_fd_sc_hd__nor2_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07735__B2 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10159_ _10160_/A _10160_/B vssd1 vssd1 vccd1 vccd1 _10159_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11819__B1 _11820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07499__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06982__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12244__B1 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07370_ _07371_/A _07371_/B vssd1 vssd1 vccd1 vccd1 _07372_/A sky130_fd_sc_hd__and2_1
XFILLER_0_29_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08463__A2 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09040_ _09821_/B _09040_/B vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_45_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_756 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08215__A2 _07181_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap110 _07974_/A vssd1 vssd1 vccd1 vccd1 _11695_/A sky130_fd_sc_hd__buf_6
XFILLER_0_40_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10558__B1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10022__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09942_ _09731_/A _09731_/B _09732_/Y vssd1 vssd1 vccd1 vccd1 _09948_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_110_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout294_A _13028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ _09873_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _09875_/B sky130_fd_sc_hd__xnor2_4
X_08824_ _08824_/A _08824_/B vssd1 vssd1 vccd1 vccd1 _08828_/B sky130_fd_sc_hd__xnor2_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ _08754_/B _08754_/C _08754_/A vssd1 vssd1 vccd1 vccd1 _08768_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__11782__B fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11286__A1 _11285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ _07707_/A _07707_/B vssd1 vssd1 vccd1 vccd1 _07706_/X sky130_fd_sc_hd__and2_1
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _08685_/B _08685_/C _08685_/A vssd1 vssd1 vccd1 vccd1 _08686_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09252__B _09252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13027__A2 _13151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07637_ _07637_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _08906_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11038__A1 _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09679__S _09679_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07568_ _09478_/B2 _07389_/B fanout26/X _09476_/A vssd1 vssd1 vccd1 vccd1 _07569_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_91_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09307_ _09362_/S _09775_/A _07539_/B _07537_/X vssd1 vssd1 vccd1 vccd1 _09309_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_36_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07499_ _08532_/B _10677_/A fanout58/X _07058_/A vssd1 vssd1 vccd1 vccd1 _07500_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10261__A2 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09238_ _07496_/A _07496_/B _07495_/A vssd1 vssd1 vccd1 vccd1 _09239_/B sky130_fd_sc_hd__a21o_1
X_09169_ reg1_val[20] reg1_val[11] _09172_/S vssd1 vssd1 vccd1 vccd1 _09169_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09403__A1 _09559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11200_ _11398_/B _11296_/B hold258/A vssd1 vssd1 vccd1 vccd1 _11200_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11210__A1 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12180_ _12179_/A _12179_/B _11197_/S vssd1 vssd1 vccd1 vccd1 _12180_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07965__B2 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11131_ _11131_/A _11131_/B vssd1 vssd1 vccd1 vccd1 _11143_/B sky130_fd_sc_hd__and2_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07717__A1 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09706__A2 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11062_ _11062_/A _11062_/B vssd1 vssd1 vccd1 vccd1 _11064_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07717__B2 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ _10013_/A _10013_/B vssd1 vssd1 vccd1 vccd1 _10016_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12788__B _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06786__B _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08142__A1 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11964_ _11964_/A _11964_/B _11964_/C vssd1 vssd1 vccd1 vccd1 _12101_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08142__B2 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10915_ _10916_/A _10916_/B vssd1 vssd1 vccd1 vccd1 _10917_/A sky130_fd_sc_hd__and2_1
X_11895_ _11721_/A _11808_/A _11810_/B vssd1 vssd1 vccd1 vccd1 _11895_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11029__A1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11029__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10846_ _10847_/A _10847_/B vssd1 vssd1 vccd1 vccd1 _10846_/X sky130_fd_sc_hd__and2_1
XFILLER_0_82_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10777_ _10720_/A _10720_/B _10721_/Y vssd1 vssd1 vccd1 vccd1 _10843_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_333 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12516_ _12516_/A _12516_/B _12516_/C vssd1 vssd1 vccd1 vccd1 _12541_/A sky130_fd_sc_hd__and3_1
X_12447_ _12607_/B _12447_/B vssd1 vssd1 vccd1 vccd1 _12448_/B sky130_fd_sc_hd__or2_1
XFILLER_0_2_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07956__B2 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07956__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12378_ _09180_/A curr_PC[0] _12556_/S vssd1 vssd1 vccd1 vccd1 _12380_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_50_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11329_ _11328_/A _11328_/B _11328_/C vssd1 vssd1 vccd1 vccd1 _11330_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06870_ _06870_/A _09383_/A _06870_/C _06870_/D vssd1 vssd1 vccd1 vccd1 _06871_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_0_66_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08381__B2 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__A1 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06696__B _07178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08540_ _08540_/A _08540_/B vssd1 vssd1 vccd1 vccd1 _08550_/A sky130_fd_sc_hd__xor2_1
X_08471_ _08471_/A _08471_/B vssd1 vssd1 vccd1 vccd1 _08492_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07422_ _07424_/A _07424_/B vssd1 vssd1 vccd1 vccd1 _07422_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07353_ _07353_/A _07353_/B vssd1 vssd1 vccd1 vccd1 _07354_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07644__B1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07284_ _11347_/A fanout98/X fanout56/X _11134_/B2 vssd1 vssd1 vccd1 vccd1 _07285_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11123__A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09023_ _09070_/C _09070_/D vssd1 vssd1 vccd1 vccd1 _09023_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_115_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold210 hold210/A vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 hold243/A vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__buf_1
Xhold221 hold221/A vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 hold232/A vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold276 hold301/X vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__buf_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold254 hold254/A vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 hold287/A vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07048__A _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09925_ _09925_/A1 _07322_/A _07322_/B fanout46/X _12760_/A vssd1 vssd1 vccd1 vccd1
+ _09926_/B sky130_fd_sc_hd__o32a_1
X_09856_ curr_PC[4] _09998_/C vssd1 vssd1 vccd1 vccd1 _09856_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__11793__A _11793_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _08806_/A _08806_/B _08806_/C vssd1 vssd1 vccd1 vccd1 _09029_/B sky130_fd_sc_hd__a21o_1
XANTENNA__09263__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06922__A2 _06567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06999_ _06999_/A _07005_/C vssd1 vssd1 vccd1 vccd1 _11933_/A sky130_fd_sc_hd__nor2_1
X_09787_ _09788_/A _09788_/B vssd1 vssd1 vccd1 vccd1 _09913_/A sky130_fd_sc_hd__and2_1
XANTENNA__08124__A1 _08774_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08738_ _08739_/A _08739_/B vssd1 vssd1 vccd1 vccd1 _08815_/A sky130_fd_sc_hd__or2_1
XFILLER_0_68_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08124__B2 _08774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08669_ _08853_/A _08669_/B vssd1 vssd1 vccd1 vccd1 _08678_/A sky130_fd_sc_hd__xnor2_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08675__A2 _08674_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10700_ _10700_/A vssd1 vssd1 vccd1 vccd1 _10832_/B sky130_fd_sc_hd__inv_2
XANTENNA__12759__A1 _07168_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11680_ _11680_/A _11680_/B vssd1 vssd1 vccd1 vccd1 _11681_/B sky130_fd_sc_hd__or2_1
X_10631_ _10629_/X _10630_/X _11831_/S vssd1 vssd1 vccd1 vccd1 _10631_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07635__B1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10562_ _10562_/A _10562_/B _10562_/C _10562_/D vssd1 vssd1 vccd1 vccd1 _10563_/B
+ sky130_fd_sc_hd__or4_1
X_13281_ _13311_/CLK _13281_/D vssd1 vssd1 vccd1 vccd1 hold240/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ _12301_/A fanout8/X _12301_/C vssd1 vssd1 vccd1 vccd1 _12301_/X sky130_fd_sc_hd__or3_1
XFILLER_0_17_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10872__A _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12232_ _09092_/X _12230_/Y _12231_/Y vssd1 vssd1 vccd1 vccd1 _12232_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10493_ _10403_/X _10524_/B _10492_/Y vssd1 vssd1 vccd1 vccd1 _10493_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_31_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12163_ _12163_/A _12215_/A vssd1 vssd1 vccd1 vccd1 _12163_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12094_ _12094_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _12095_/B sky130_fd_sc_hd__nand2_1
X_11114_ _11604_/A _11114_/B vssd1 vssd1 vccd1 vccd1 _11116_/B sky130_fd_sc_hd__xnor2_1
X_11045_ _11045_/A _11045_/B vssd1 vssd1 vccd1 vccd1 _11046_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12996_ _11499_/A _13020_/B2 hold111/X vssd1 vssd1 vccd1 vccd1 hold112/A sky130_fd_sc_hd__o21a_1
XANTENNA__10112__A _10249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12998__A1 _07317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11947_ _11947_/A _11947_/B vssd1 vssd1 vccd1 vccd1 _11948_/B sky130_fd_sc_hd__or2_1
XANTENNA__11670__A1 _07068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11878_ _11878_/A _11878_/B _11878_/C vssd1 vssd1 vccd1 vccd1 _11879_/B sky130_fd_sc_hd__and3_1
X_10829_ _10664_/A _10664_/B _10663_/A vssd1 vssd1 vccd1 vccd1 _10834_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_82_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09067__B _11559_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07971_ _09580_/A _07971_/B _07971_/C vssd1 vssd1 vccd1 vccd1 _07977_/A sky130_fd_sc_hd__nand3_1
X_06922_ instruction[3] _06567_/B _06572_/X instruction[40] _09199_/B vssd1 vssd1
+ vccd1 vccd1 _06923_/C sky130_fd_sc_hd__o221a_1
X_09710_ _12223_/B1 _09665_/X _09666_/Y _09709_/X vssd1 vssd1 vccd1 vccd1 _09710_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_93_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06853_ _06843_/A _06852_/X _06837_/Y vssd1 vssd1 vccd1 vccd1 _12225_/B sky130_fd_sc_hd__a21bo_1
X_09641_ _09641_/A _09641_/B vssd1 vssd1 vccd1 vccd1 _09642_/B sky130_fd_sc_hd__and2_2
X_06784_ reg2_val[0] _06778_/B _06649_/A _06783_/X vssd1 vssd1 vccd1 vccd1 _06784_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__11118__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09572_ _10301_/A _09572_/B vssd1 vssd1 vccd1 vccd1 _09573_/B sky130_fd_sc_hd__xnor2_1
X_08523_ _08527_/A _08527_/B _08508_/X vssd1 vssd1 vccd1 vccd1 _09011_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__11110__B1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08454_ _08488_/A _08460_/B _08447_/X vssd1 vssd1 vccd1 vccd1 _08484_/B sky130_fd_sc_hd__a21o_1
X_08385_ _08385_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _08399_/B sky130_fd_sc_hd__xnor2_1
X_07405_ _09610_/A _07405_/B vssd1 vssd1 vccd1 vccd1 _08896_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07336_ _08680_/B _12736_/A fanout30/X _09772_/A vssd1 vssd1 vccd1 vccd1 _07337_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09006_ _08619_/B _08619_/A _08339_/B _08339_/A vssd1 vssd1 vccd1 vccd1 _09006_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_103_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07267_ _07267_/A _07267_/B vssd1 vssd1 vccd1 vccd1 _07270_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10692__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07198_ _08217_/B fanout94/X fanout55/X _12752_/A vssd1 vssd1 vccd1 vccd1 _07199_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08593__B2 _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12412__A _12583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ _10819_/A _09908_/B vssd1 vssd1 vccd1 vccd1 _09909_/C sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout72_A _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ _12124_/B _10119_/C hold224/A vssd1 vssd1 vccd1 vccd1 _09839_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09542__B1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__A1 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10152__B2 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12850_ _13072_/A _13073_/A _13072_/B vssd1 vssd1 vccd1 vccd1 _13078_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09721__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11801_ _11802_/A _11802_/B vssd1 vssd1 vccd1 vccd1 _11888_/A sky130_fd_sc_hd__nand2_1
X_12781_ _09252_/B _12781_/A2 hold69/X _13166_/A vssd1 vssd1 vccd1 vccd1 _13212_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11101__B1 _11838_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09845__A1 _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07320__A2 _07317_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11732_ _11767_/B _11731_/Y _09110_/X vssd1 vssd1 vccd1 vccd1 _11732_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10455__A2 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11663_ _09115_/X _10752_/X _10765_/Y _09184_/X _11662_/X vssd1 vssd1 vccd1 vccd1
+ _11663_/X sky130_fd_sc_hd__o221a_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10614_ _12278_/A _11000_/A _10774_/A vssd1 vssd1 vccd1 vccd1 _10614_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11594_ _11595_/A _11595_/B vssd1 vssd1 vccd1 vccd1 _11706_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_122_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10545_ _10662_/B _10545_/B vssd1 vssd1 vccd1 vccd1 _10571_/A sky130_fd_sc_hd__or2_2
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13264_ _13264_/CLK _13264_/D vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_51_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10476_ _10476_/A _10476_/B vssd1 vssd1 vccd1 vccd1 _10477_/B sky130_fd_sc_hd__xor2_4
X_13195_ _13296_/CLK _13195_/D vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__dfxtp_1
X_12215_ _12215_/A _12215_/B vssd1 vssd1 vccd1 vccd1 _12313_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_121_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12146_ _12205_/A _12301_/A fanout8/X fanout27/X vssd1 vssd1 vccd1 vccd1 _12147_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12077_ _12206_/A _12077_/B vssd1 vssd1 vccd1 vccd1 _12081_/A sky130_fd_sc_hd__xor2_1
X_11028_ _11028_/A _11028_/B vssd1 vssd1 vccd1 vccd1 _11045_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09631__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12979_ hold144/A _13013_/A2 _13170_/B hold95/X _13066_/A vssd1 vssd1 vccd1 vccd1
+ hold96/A sky130_fd_sc_hd__o221a_1
XANTENNA__09836__A1 _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08170_ _08819_/B2 _08348_/B _07181_/Y _12730_/A vssd1 vssd1 vccd1 vccd1 _08171_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_103_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_38 reg2_val[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_16 reg1_val[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 reg1_val[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12199__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 reg2_val[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07121_ _09467_/A _07121_/B vssd1 vssd1 vccd1 vccd1 _07160_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07052_ _07068_/A _07052_/B vssd1 vssd1 vccd1 vccd1 _07111_/C sky130_fd_sc_hd__and2_1
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12371__A2 _12370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10382__A1 _09201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07954_ _07955_/A _07955_/B vssd1 vssd1 vccd1 vccd1 _07954_/X sky130_fd_sc_hd__or2_1
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06905_ instruction[25] _06915_/B vssd1 vssd1 vccd1 vccd1 _06905_/X sky130_fd_sc_hd__or2_1
X_07885_ _07885_/A _07885_/B vssd1 vssd1 vccd1 vccd1 _07887_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__06889__A1 _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07045__B _07046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06836_ reg1_val[28] _12250_/A vssd1 vssd1 vccd1 vccd1 _06845_/A sky130_fd_sc_hd__and2_1
XANTENNA__11331__B1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09624_ _10894_/A _09624_/B vssd1 vssd1 vccd1 vccd1 _09628_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07550__A2 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06884__B _06898_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09555_ _09541_/Y _09542_/X _09547_/Y _09554_/X vssd1 vssd1 vccd1 vccd1 _09555_/Y
+ sky130_fd_sc_hd__o211ai_1
X_06767_ _06783_/A _06649_/A _12578_/B _06765_/X vssd1 vssd1 vccd1 vccd1 _06767_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__12378__S _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06698_ _06696_/Y _06698_/B vssd1 vssd1 vccd1 vccd1 _11187_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_93_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08506_ _08506_/A _08506_/B vssd1 vssd1 vccd1 vccd1 _08509_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_38_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10437__A2 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09486_ _09487_/A _09487_/B vssd1 vssd1 vccd1 vccd1 _09486_/Y sky130_fd_sc_hd__nor2_1
X_08437_ _07969_/A _09618_/B2 _09618_/A1 _12734_/A vssd1 vssd1 vccd1 vccd1 _08438_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08368_ _08403_/B _08403_/A vssd1 vssd1 vccd1 vccd1 _08368_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_46_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08299_ _08299_/A _08299_/B vssd1 vssd1 vccd1 vccd1 _08301_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_104_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07319_ _07319_/A _07319_/B vssd1 vssd1 vccd1 vccd1 _07319_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10330_ _11688_/A fanout47/X _11603_/A fanout70/X vssd1 vssd1 vccd1 vccd1 _10331_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10261_ _06866_/D _09383_/B _10253_/Y _10254_/X _10260_/X vssd1 vssd1 vccd1 vccd1
+ _10261_/X sky130_fd_sc_hd__o221a_1
X_12000_ _12000_/A _12000_/B _11991_/X vssd1 vssd1 vccd1 vccd1 _12000_/X sky130_fd_sc_hd__or3b_1
X_10192_ _10192_/A _10192_/B vssd1 vssd1 vccd1 vccd1 _10193_/B sky130_fd_sc_hd__or2_1
XANTENNA__08318__A1 _09283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12142__A _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08318__B2 _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07236__A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ _13169_/A hold238/X vssd1 vssd1 vccd1 vccd1 _13221_/D sky130_fd_sc_hd__and2_1
XANTENNA__11322__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12833_ hold29/X hold279/A vssd1 vssd1 vccd1 vccd1 _13029_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ hold88/X _12778_/B vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__or2_1
XFILLER_0_84_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11715_ _11715_/A _11715_/B vssd1 vssd1 vccd1 vccd1 _11716_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ reg1_val[28] _12708_/B vssd1 vssd1 vccd1 vccd1 _12696_/B sky130_fd_sc_hd__nor2_1
X_11646_ _06865_/A _11560_/X _06668_/A vssd1 vssd1 vccd1 vccd1 _11646_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_71_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11577_ _07077_/A _12250_/B _11099_/B reg1_val[19] vssd1 vssd1 vccd1 vccd1 _11577_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07057__A1 _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13316_ _13318_/CLK hold156/X vssd1 vssd1 vccd1 vccd1 hold154/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_52_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10528_ _10658_/A _10528_/B vssd1 vssd1 vccd1 vccd1 _10705_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_122_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13247_ _13248_/CLK hold233/X vssd1 vssd1 vccd1 vccd1 hold231/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08557__B2 _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08557__A1 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ _10459_/A _10459_/B vssd1 vssd1 vccd1 vccd1 _10461_/C sky130_fd_sc_hd__xnor2_2
X_13178_ hold186/A hold298/A hold137/X hold154/X vssd1 vssd1 vccd1 vccd1 hold155/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__09626__A _10578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12129_ _09198_/X _12123_/X _12124_/Y _12128_/X vssd1 vssd1 vccd1 vccd1 _12129_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07146__A _08695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07670_ _06864_/A _10677_/A _07157_/Y _08758_/A2 vssd1 vssd1 vccd1 vccd1 _07671_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10667__A2 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ reg2_val[31] _06752_/A vssd1 vssd1 vccd1 vccd1 _06621_/X sky130_fd_sc_hd__and2_1
XFILLER_0_59_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06552_ _06881_/C _06881_/B instruction[2] vssd1 vssd1 vccd1 vccd1 _06552_/X sky130_fd_sc_hd__or3b_4
XFILLER_0_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09340_ _08594_/B _12131_/A _09338_/X _09339_/Y _11381_/A vssd1 vssd1 vccd1 vccd1
+ _09340_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_75_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09271_ _09271_/A _09271_/B vssd1 vssd1 vccd1 vccd1 _09272_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09285__A2 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08222_ _07134_/A fanout94/X _12752_/A _08758_/A2 vssd1 vssd1 vccd1 vccd1 _08223_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08153_ _08153_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _08211_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout122_A _07324_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08084_ _08841_/A1 _08776_/B1 _10433_/A _08477_/B vssd1 vssd1 vccd1 vccd1 _08085_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_70_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07104_ reg1_val[3] _07104_/B vssd1 vssd1 vccd1 vccd1 _08311_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_43_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07035_ _07031_/A _07031_/B _08855_/A vssd1 vssd1 vccd1 vccd1 _07035_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08440__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12344__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08986_ _08986_/A _08986_/B vssd1 vssd1 vccd1 vccd1 _08989_/B sky130_fd_sc_hd__xor2_2
X_07937_ _07937_/A _07937_/B _07937_/C vssd1 vssd1 vccd1 vccd1 _08068_/A sky130_fd_sc_hd__or3_2
XANTENNA__07771__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07056__A _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07868_ _07079_/A _07079_/B _07134_/A vssd1 vssd1 vccd1 vccd1 _07871_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_3_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11855__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07799_ _08819_/B2 _09752_/B fanout14/X _12730_/A vssd1 vssd1 vccd1 vccd1 _07800_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06819_ reg1_val[17] _07049_/C vssd1 vssd1 vccd1 vccd1 _06819_/Y sky130_fd_sc_hd__nand2_1
X_09607_ _10527_/A _10557_/A fanout58/X _10452_/B2 vssd1 vssd1 vccd1 vccd1 _09608_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09538_ _09538_/A _09538_/B vssd1 vssd1 vccd1 vccd1 _09539_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_66_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09276__A2 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout35_A fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12280__A1 _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09469_ _09620_/A _09469_/B vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__xnor2_2
X_11500_ _11618_/A _11500_/B vssd1 vssd1 vccd1 vccd1 _11504_/B sky130_fd_sc_hd__or2_1
X_12480_ reg1_val[15] curr_PC[15] _12524_/S vssd1 vssd1 vccd1 vccd1 _12482_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_81_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08236__B1 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11431_ _11431_/A _12304_/B vssd1 vssd1 vccd1 vccd1 _11432_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09984__B1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ _11362_/A _11362_/B vssd1 vssd1 vccd1 vccd1 _11364_/B sky130_fd_sc_hd__xnor2_1
X_13101_ _13166_/A _13101_/B vssd1 vssd1 vccd1 vccd1 _13297_/D sky130_fd_sc_hd__and2_1
XFILLER_0_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10313_ _10201_/B _10204_/B _10201_/A vssd1 vssd1 vccd1 vccd1 _10323_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_21_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11293_ _11291_/Y _11293_/B vssd1 vssd1 vccd1 vccd1 _11294_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_21_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13032_ hold250/X _12721_/B _13031_/X _12722_/A vssd1 vssd1 vccd1 vccd1 hold251/A
+ sky130_fd_sc_hd__a22o_1
X_10244_ _10750_/S _09161_/X _11195_/C vssd1 vssd1 vccd1 vccd1 _10244_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09446__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06789__B _10249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07211__B2 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07211__A1 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10175_ _10175_/A _10175_/B vssd1 vssd1 vccd1 vccd1 _10192_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07762__A2 _08774_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout180 _12742_/B vssd1 vssd1 vccd1 vccd1 _12786_/B sky130_fd_sc_hd__clkbuf_4
Xfanout191 _13170_/B vssd1 vssd1 vccd1 vccd1 _13020_/A2 sky130_fd_sc_hd__buf_4
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12816_ hold268/X hold63/X vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_56_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12747_ _10551_/A _12980_/A2 hold55/X _13179_/A vssd1 vssd1 vccd1 vccd1 _13195_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08475__B1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12678_ _12678_/A _12678_/B _12678_/C _12678_/D vssd1 vssd1 vccd1 vccd1 _12678_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_72_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11629_ _11629_/A _11629_/B vssd1 vssd1 vccd1 vccd1 _11632_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_108_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09727__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09075__B _11820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08840_ _08840_/A _08840_/B vssd1 vssd1 vccd1 vccd1 _08844_/A sky130_fd_sc_hd__xor2_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _10306_/A _08685_/A _08685_/X vssd1 vssd1 vccd1 vccd1 _08784_/A sky130_fd_sc_hd__o21bai_2
XFILLER_0_85_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06961__B1 _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07307__C _10180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07722_ _07722_/A _07722_/B vssd1 vssd1 vccd1 vccd1 _07726_/A sky130_fd_sc_hd__xor2_2
X_07653_ _07632_/A _07632_/B _07651_/B _07652_/X vssd1 vssd1 vccd1 vccd1 _07690_/B
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_79_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06604_ reg1_val[24] _07126_/B vssd1 vssd1 vccd1 vccd1 _06604_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07584_ _07584_/A _07584_/B vssd1 vssd1 vccd1 vccd1 _07587_/A sky130_fd_sc_hd__xnor2_4
X_09323_ _09323_/A _09323_/B vssd1 vssd1 vccd1 vccd1 _09325_/B sky130_fd_sc_hd__xnor2_2
X_06535_ hold51/X vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__inv_2
XFILLER_0_48_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09254_ _09255_/B _09255_/C _09610_/A vssd1 vssd1 vccd1 vccd1 _09256_/B sky130_fd_sc_hd__a21o_1
X_08205_ _08205_/A _08205_/B vssd1 vssd1 vccd1 vccd1 _08213_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_118_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09185_ _09202_/A _09199_/B vssd1 vssd1 vccd1 vccd1 _11381_/A sky130_fd_sc_hd__nor2_8
XFILLER_0_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08136_ _08146_/A _08146_/B vssd1 vssd1 vccd1 vccd1 _08136_/X sky130_fd_sc_hd__and2_1
X_08067_ _07937_/A _07937_/B _07937_/C vssd1 vssd1 vccd1 vccd1 _08068_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07018_ _07018_/A _07319_/A vssd1 vssd1 vccd1 vccd1 _07175_/D sky130_fd_sc_hd__or2_1
XANTENNA__10328__A1 _12774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10328__B2 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08969_ _08969_/A _08969_/B vssd1 vssd1 vccd1 vccd1 _08970_/B sky130_fd_sc_hd__xor2_1
X_11980_ _06833_/B _11979_/Y _12322_/S vssd1 vssd1 vccd1 vccd1 _11980_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_98_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07514__A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ _10929_/Y _10931_/B vssd1 vssd1 vccd1 vccd1 _10938_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10862_ _06808_/Y _10861_/Y _11738_/S vssd1 vssd1 vccd1 vccd1 _10863_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12601_ _12600_/A _12597_/Y _12599_/B vssd1 vssd1 vccd1 vccd1 _12605_/A sky130_fd_sc_hd__o21a_2
X_10793_ _10793_/A _10793_/B vssd1 vssd1 vccd1 vccd1 _10795_/B sky130_fd_sc_hd__xor2_1
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ _12539_/B _12532_/B vssd1 vssd1 vccd1 vccd1 new_PC[22] sky130_fd_sc_hd__xnor2_4
XFILLER_0_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10803__A2 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12463_ _12464_/A _12464_/B _12464_/C vssd1 vssd1 vccd1 vccd1 _12471_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_53_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11414_ _11414_/A _11414_/B vssd1 vssd1 vccd1 vccd1 _11416_/B sky130_fd_sc_hd__xor2_2
X_12394_ _12394_/A _12394_/B _12394_/C vssd1 vssd1 vccd1 vccd1 _12395_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07432__B2 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07432__A1 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11345_ _11704_/A fanout27/X _12205_/A _11688_/A vssd1 vssd1 vccd1 vccd1 _11346_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09709__B1 _09708_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11276_ _11068_/A _11170_/Y _11172_/B vssd1 vssd1 vccd1 vccd1 _11276_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_120_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13015_ hold52/X _06537_/A _13151_/A2 hold48/X rst vssd1 vssd1 vccd1 vccd1 hold53/A
+ sky130_fd_sc_hd__a221o_1
X_10227_ _10227_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10486_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07735__A2 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09904__A _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10158_ _10158_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _10160_/B sky130_fd_sc_hd__xnor2_2
X_10089_ _10090_/A _10090_/B vssd1 vssd1 vccd1 vccd1 _10089_/X sky130_fd_sc_hd__and2_1
XFILLER_0_89_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07499__A1 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07499__B2 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08448__B1 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10785__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06982__B _06987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10255__B1 _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07120__B1 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10007__B1 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11755__B1 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10558__A1 _07308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_768 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09941_ _09797_/A _09796_/B _09794_/Y vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12180__B1 _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10025__A _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09872_ _10306_/A _09872_/B vssd1 vssd1 vccd1 vccd1 _09873_/B sky130_fd_sc_hd__xor2_4
X_08823_ _08824_/A _08824_/B vssd1 vssd1 vccd1 vccd1 _08891_/A sky130_fd_sc_hd__and2_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07854__A_N _07855_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08754_ _08754_/A _08754_/B _08754_/C vssd1 vssd1 vccd1 vccd1 _08768_/A sky130_fd_sc_hd__and3_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ _07707_/A _07707_/B vssd1 vssd1 vccd1 vccd1 _07705_/X sky130_fd_sc_hd__or2_1
XANTENNA__07334__A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _08685_/A _08685_/B _08685_/C vssd1 vssd1 vccd1 vccd1 _08685_/X sky130_fd_sc_hd__and3_1
XFILLER_0_68_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _11604_/A _07636_/B vssd1 vssd1 vccd1 vccd1 _07637_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08439__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07567_ _07250_/A _07250_/B _07248_/Y vssd1 vssd1 vccd1 vccd1 _07573_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09306_ _09306_/A _09306_/B vssd1 vssd1 vccd1 vccd1 _09309_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_8_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11994__B1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09237_ _09237_/A _09237_/B vssd1 vssd1 vccd1 vccd1 _09239_/A sky130_fd_sc_hd__nand2_1
X_07498_ _10658_/A _07498_/B vssd1 vssd1 vccd1 vccd1 _07502_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09168_ _09164_/X _09167_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09168_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08119_ _08059_/A _08058_/C _08058_/B vssd1 vssd1 vccd1 vccd1 _08120_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_102_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ _08935_/X _08979_/Y _09082_/B _09098_/X _08998_/X vssd1 vssd1 vccd1 vccd1
+ _09100_/B sky130_fd_sc_hd__o221ai_4
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11130_ _11131_/A _11131_/B vssd1 vssd1 vccd1 vccd1 _11262_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12171__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11061_ _11062_/A _11062_/B vssd1 vssd1 vccd1 vccd1 _11171_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07717__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ _10012_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _10013_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12150__A _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08142__A2 _08348_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11963_ _11964_/A _11964_/B _11964_/C vssd1 vssd1 vccd1 vccd1 _12101_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10914_ _11499_/A _10914_/B vssd1 vssd1 vccd1 vccd1 _10916_/B sky130_fd_sc_hd__xnor2_1
X_11894_ _11894_/A _11894_/B vssd1 vssd1 vccd1 vccd1 _11894_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11029__A2 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10845_ _10847_/A _10847_/B vssd1 vssd1 vccd1 vccd1 _10959_/B sky130_fd_sc_hd__or2_1
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10776_ _10776_/A vssd1 vssd1 vccd1 vccd1 _10776_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_27_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12515_ _12515_/A _12515_/B _12515_/C vssd1 vssd1 vccd1 vccd1 _12539_/A sky130_fd_sc_hd__or3_1
XFILLER_0_42_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12446_ _12607_/B _12447_/B vssd1 vssd1 vccd1 vccd1 _12457_/A sky130_fd_sc_hd__nand2_1
X_12377_ _12370_/B _12250_/B _12376_/X _12382_/S vssd1 vssd1 vccd1 vccd1 dest_val[31]
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_2_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07956__A2 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11328_ _11328_/A _11328_/B _11328_/C vssd1 vssd1 vccd1 vccd1 _11444_/B sky130_fd_sc_hd__and3_1
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09158__A1 _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11259_ _11160_/A _11159_/B _11159_/A vssd1 vssd1 vccd1 vccd1 _11266_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__08381__A2 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08470_ _08492_/A vssd1 vssd1 vccd1 vccd1 _08470_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06695__A2 _12658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07421_ _07421_/A _07421_/B vssd1 vssd1 vccd1 vccd1 _07424_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07352_ _07353_/A _07353_/B vssd1 vssd1 vccd1 vccd1 _07352_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11976__B1 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07644__B2 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07644__A1 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08841__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07283_ _07205_/A _07205_/B _07208_/Y vssd1 vssd1 vccd1 vccd1 _07293_/A sky130_fd_sc_hd__o21ai_1
X_09022_ _09022_/A _09022_/B vssd1 vssd1 vccd1 vccd1 _09066_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_115_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold200 hold200/A vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_3_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13312_/CLK sky130_fd_sc_hd__clkbuf_8
Xhold211 hold211/A vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09397__A1 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09397__B2 _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold244 hold244/A vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold222 hold222/A vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 hold233/A vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12235__A _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold277 hold277/A vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 hold255/A vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 hold266/A vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__buf_1
XANTENNA__06988__C_N _06987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold299 hold299/A vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 hold288/A vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ _10180_/A _09924_/B vssd1 vssd1 vccd1 vccd1 _09928_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09855_ _09820_/X _09823_/X _09827_/X _09854_/X _12382_/S vssd1 vssd1 vccd1 vccd1
+ _09855_/X sky130_fd_sc_hd__o41a_1
XANTENNA__11793__B _12255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _08806_/A _08806_/B _08806_/C vssd1 vssd1 vccd1 vccd1 _08806_/X sky130_fd_sc_hd__and3_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07064__A _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06998_ _06999_/A _07005_/C vssd1 vssd1 vccd1 vccd1 _07000_/A sky130_fd_sc_hd__and2_1
X_09786_ _10565_/A _09786_/B vssd1 vssd1 vccd1 vccd1 _09788_/B sky130_fd_sc_hd__xnor2_1
X_08737_ _08857_/A _08737_/B vssd1 vssd1 vccd1 vccd1 _08739_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08124__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _07173_/Y _10811_/A _10694_/A _07182_/X vssd1 vssd1 vccd1 vccd1 _08669_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07619_ _07619_/A _07619_/B vssd1 vssd1 vccd1 vccd1 _07620_/B sky130_fd_sc_hd__xor2_4
XANTENNA__12759__A2 _12781_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ _10630_/A _10630_/B vssd1 vssd1 vccd1 vccd1 _10630_/X sky130_fd_sc_hd__xor2_1
XANTENNA__10629__S _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ _08599_/A vssd1 vssd1 vccd1 vccd1 _08599_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07635__B2 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07635__A1 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10561_ _10562_/A _10562_/B _10562_/C _10562_/D vssd1 vssd1 vccd1 vccd1 _10705_/B
+ sky130_fd_sc_hd__o22a_1
X_13280_ _13280_/CLK hold39/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12300_ _12257_/A _12257_/B _12255_/Y fanout19/X vssd1 vssd1 vccd1 vccd1 _12307_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_10492_ _10403_/X _10524_/B _09110_/X vssd1 vssd1 vccd1 vccd1 _10492_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09388__A1 _09679_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12231_ _09092_/X _12230_/Y _11184_/A vssd1 vssd1 vccd1 vccd1 _12231_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12931__A2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07239__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ _12035_/A _12097_/A _12099_/B vssd1 vssd1 vccd1 vccd1 _12162_/X sky130_fd_sc_hd__a21o_1
X_12093_ _12094_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _12160_/B sky130_fd_sc_hd__or2_1
X_11113_ _12150_/A fanout47/X _11603_/A _12150_/B vssd1 vssd1 vccd1 vccd1 _11114_/B
+ sky130_fd_sc_hd__o22a_1
X_11044_ _11044_/A _11044_/B vssd1 vssd1 vccd1 vccd1 _11045_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07571__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12995_ hold116/A _13013_/A2 _13020_/A2 hold110/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold111/A sky130_fd_sc_hd__o221a_1
XFILLER_0_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12998__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11946_ _11947_/A _11947_/B vssd1 vssd1 vccd1 vccd1 _12025_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11670__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11877_ _11878_/A _11878_/B _11878_/C vssd1 vssd1 vccd1 vccd1 _11932_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10828_ _10708_/A _10708_/B _10711_/A vssd1 vssd1 vccd1 vccd1 _10839_/A sky130_fd_sc_hd__o21ai_2
X_10759_ _09385_/C _10877_/B hold291/A vssd1 vssd1 vccd1 vccd1 _10759_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12429_ _12429_/A _12429_/B _12429_/C vssd1 vssd1 vccd1 vccd1 _12430_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07970_ _07308_/A _07308_/B _09772_/A vssd1 vssd1 vccd1 vccd1 _07971_/C sky130_fd_sc_hd__a21o_1
X_06921_ instruction[17] _09205_/B _09184_/B _06752_/A vssd1 vssd1 vccd1 vccd1 _06923_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__06988__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06852_ _06620_/B _06851_/X _06838_/Y vssd1 vssd1 vccd1 vccd1 _06852_/X sky130_fd_sc_hd__a21o_1
X_09640_ _09640_/A _09640_/B vssd1 vssd1 vccd1 vccd1 _09641_/B sky130_fd_sc_hd__or2_1
X_06783_ _06783_/A _12563_/B vssd1 vssd1 vccd1 vccd1 _06783_/X sky130_fd_sc_hd__and2_1
X_09571_ fanout36/X _10144_/B2 _10433_/A _08821_/B vssd1 vssd1 vccd1 vccd1 _09572_/B
+ sky130_fd_sc_hd__o22a_1
X_08522_ _08522_/A vssd1 vssd1 vccd1 vccd1 _08527_/B sky130_fd_sc_hd__inv_2
XFILLER_0_89_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08453_ _08453_/A _08453_/B vssd1 vssd1 vccd1 vccd1 _08460_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07314__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11661__A2 _06653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout152_A _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07404_ _08532_/B _12768_/A _12766_/A _07058_/A vssd1 vssd1 vccd1 vccd1 _07405_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_107_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08384_ _08418_/A _08418_/B _08380_/X vssd1 vssd1 vccd1 vccd1 _08399_/A sky130_fd_sc_hd__o21a_1
X_07335_ _07335_/A _07335_/B vssd1 vssd1 vccd1 vccd1 _07380_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_45_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09539__A _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07266_ _07265_/B _07266_/B vssd1 vssd1 vccd1 vccd1 _07267_/B sky130_fd_sc_hd__nand2b_1
X_09005_ _08258_/Y _08626_/B _08256_/Y vssd1 vssd1 vccd1 vccd1 _09022_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_115_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08443__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07197_ _07197_/A _07197_/B vssd1 vssd1 vccd1 vccd1 _07197_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__07059__A _07068_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08593__A2 _09283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__A1 _09600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06898__A _06898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12126__B1 _07153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09907_ fanout62/X fanout95/X fanout54/X fanout77/X vssd1 vssd1 vccd1 vccd1 _09908_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09274__A _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09838_ hold237/A hold297/A _13218_/Q hold211/A vssd1 vssd1 vccd1 vccd1 _10119_/C
+ sky130_fd_sc_hd__or4_2
XANTENNA__06628__A2_N _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout65_A _12774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10152__A2 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ _09770_/A _09770_/B vssd1 vssd1 vccd1 vccd1 _09769_/Y sky130_fd_sc_hd__nand2_1
X_11800_ _11800_/A _11800_/B vssd1 vssd1 vccd1 vccd1 _11802_/B sky130_fd_sc_hd__xnor2_1
X_12780_ hold68/X _12786_/B vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__or2_1
XFILLER_0_96_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _12230_/A _11731_/B vssd1 vssd1 vccd1 vccd1 _11731_/Y sky130_fd_sc_hd__nand2_1
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _06654_/A _12243_/B1 _11099_/B reg1_val[20] _11661_/Y vssd1 vssd1 vccd1 vccd1
+ _11662_/X sky130_fd_sc_hd__o221a_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10613_ _10730_/B _10613_/B vssd1 vssd1 vccd1 vccd1 _10774_/A sky130_fd_sc_hd__xnor2_2
X_11593_ _12019_/A _11593_/B vssd1 vssd1 vccd1 vccd1 _11595_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10544_ _10543_/B _10544_/B vssd1 vssd1 vccd1 vccd1 _10545_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_107_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08353__A _08544_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13263_ _13264_/CLK _13263_/D vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12365__B1 _09198_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10475_ _10475_/A _10475_/B vssd1 vssd1 vccd1 vccd1 _10476_/B sky130_fd_sc_hd__xor2_4
X_13194_ _13318_/CLK _13194_/D vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfxtp_1
X_12214_ _12214_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _12312_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09230__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12145_ _12148_/A vssd1 vssd1 vccd1 vccd1 _12145_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07792__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09184__A _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12117__B1 _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12076_ _12205_/A fanout19/X _12301_/A _07389_/B vssd1 vssd1 vccd1 vccd1 _12077_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10679__B1 _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11027_ _11604_/A _11027_/B vssd1 vssd1 vccd1 vccd1 _11028_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12978_ _07030_/B _12744_/B hold145/X vssd1 vssd1 vccd1 vccd1 _13259_/D sky130_fd_sc_hd__a21boi_1
XANTENNA__09836__A2 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09297__B1 _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11929_ curr_PC[22] curr_PC[23] _11929_/C vssd1 vssd1 vccd1 vccd1 _12070_/C sky130_fd_sc_hd__and3_2
XFILLER_0_86_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_39 reg2_val[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_17 reg1_val[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 reg1_val[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ _09618_/B2 _10557_/A _09618_/A1 _07119_/Y vssd1 vssd1 vccd1 vccd1 _07121_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07051_ _07051_/A _07051_/B _07050_/C vssd1 vssd1 vccd1 vccd1 _07129_/B sky130_fd_sc_hd__or3b_2
XANTENNA__09078__B _11820_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12371__A3 wire201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07953_ _10578_/A _07953_/B vssd1 vssd1 vccd1 vccd1 _07955_/B sky130_fd_sc_hd__xnor2_1
X_06904_ instruction[16] _06904_/B vssd1 vssd1 vccd1 vccd1 dest_idx[5] sky130_fd_sc_hd__and2_4
X_07884_ _07885_/A _07885_/B vssd1 vssd1 vccd1 vccd1 _08014_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11331__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06835_ reg1_val[29] _07243_/A vssd1 vssd1 vccd1 vccd1 _06835_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07535__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11331__B2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ fanout62/X fanout98/X fanout56/X fanout77/X vssd1 vssd1 vccd1 vccd1 _09624_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_78_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08438__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09554_ _06777_/B _12243_/B1 _09383_/B _06870_/A _09553_/X vssd1 vssd1 vccd1 vccd1
+ _09554_/X sky130_fd_sc_hd__o221a_1
X_06766_ _06783_/A _06649_/A _12578_/B _06765_/X vssd1 vssd1 vccd1 vccd1 _06964_/A
+ sky130_fd_sc_hd__a31oi_4
X_06697_ reg1_val[15] _07178_/A vssd1 vssd1 vccd1 vccd1 _06698_/B sky130_fd_sc_hd__nand2_1
X_08505_ _08505_/A _08505_/B vssd1 vssd1 vccd1 vccd1 _09052_/A sky130_fd_sc_hd__xnor2_2
X_09485_ _09485_/A _09485_/B vssd1 vssd1 vccd1 vccd1 _09487_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_4_13_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08436_ _08436_/A _08436_/B vssd1 vssd1 vccd1 vccd1 _08453_/A sky130_fd_sc_hd__xnor2_2
X_08367_ _08367_/A _08367_/B vssd1 vssd1 vccd1 vccd1 _08403_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07318_ _07318_/A _07319_/B vssd1 vssd1 vccd1 vccd1 _10551_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08173__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ _08298_/A _08298_/B vssd1 vssd1 vccd1 vccd1 _08301_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_104_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09269__A _10184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07249_ _07249_/A _07249_/B vssd1 vssd1 vccd1 vccd1 _07250_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10260_ _06742_/Y _09191_/X _10255_/X _10259_/X vssd1 vssd1 vccd1 vccd1 _10260_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_103_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11738__S _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _10192_/A _10192_/B vssd1 vssd1 vccd1 vccd1 _10193_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08318__A2 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12901_ hold217/X _12955_/A2 _13168_/B1 hold224/X vssd1 vssd1 vccd1 vccd1 hold238/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11322__A1 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11322__B2 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13075__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12832_ _13025_/A _13025_/B _12830_/A vssd1 vssd1 vccd1 vccd1 _13030_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08348__A _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ hold25/X _12778_/B _12762_/Y _13147_/A vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__o211a_1
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07252__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11714_ _11715_/A _11715_/B vssd1 vssd1 vccd1 vccd1 _11809_/A sky130_fd_sc_hd__or2_1
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ reg1_val[28] _12708_/B vssd1 vssd1 vccd1 vccd1 _12705_/A sky130_fd_sc_hd__and2_1
XFILLER_0_37_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11645_ _12332_/B _09069_/A _09073_/C _11184_/A vssd1 vssd1 vccd1 vccd1 _11645_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11502__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08083__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11576_ _06668_/A _09383_/B _09191_/X vssd1 vssd1 vccd1 vccd1 _11576_/X sky130_fd_sc_hd__o21a_1
XANTENNA__09179__A _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09451__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13315_ _13318_/CLK hold300/X vssd1 vssd1 vccd1 vccd1 hold186/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10527_ _10527_/A fanout9/X vssd1 vssd1 vccd1 vccd1 _10528_/B sky130_fd_sc_hd__nor2_2
X_13246_ _13248_/CLK hold167/X vssd1 vssd1 vccd1 vccd1 _13246_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09203__B1 _09198_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10458_ _10458_/A _10458_/B vssd1 vssd1 vccd1 vccd1 _10459_/B sky130_fd_sc_hd__xor2_2
XANTENNA__08557__A2 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13177_ hold154/X _12721_/B _12718_/Y _12722_/A vssd1 vssd1 vccd1 vccd1 _13179_/B
+ sky130_fd_sc_hd__a22o_1
X_10389_ reg1_val[8] curr_PC[8] vssd1 vssd1 vccd1 vccd1 _10389_/Y sky130_fd_sc_hd__nor2_1
X_12128_ _09183_/Y _09972_/Y _09978_/X _12373_/A1 _12127_/X vssd1 vssd1 vccd1 vccd1
+ _12128_/X sky130_fd_sc_hd__a221o_1
XANTENNA__09118__S _12726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07146__B _07148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12059_ hold173/A _12059_/B vssd1 vssd1 vccd1 vccd1 _12122_/B sky130_fd_sc_hd__or2_1
XANTENNA__11383__S _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06620_ _06843_/A _06620_/B vssd1 vssd1 vccd1 vccd1 _06632_/B sky130_fd_sc_hd__nand2_1
X_06551_ instruction[1] instruction[2] instruction[0] pred_val vssd1 vssd1 vccd1 vccd1
+ _06915_/B sky130_fd_sc_hd__and4b_4
XANTENNA__11077__B1 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09270_ _09271_/A _09271_/B vssd1 vssd1 vccd1 vccd1 _09438_/B sky130_fd_sc_hd__or2_1
X_08221_ _08775_/A _08221_/B vssd1 vssd1 vccd1 vccd1 _08228_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08152_ _08153_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _08157_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_7_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08083_ _08775_/A _08083_/B vssd1 vssd1 vccd1 vccd1 _08089_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09993__A1 _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ reg1_val[0] _12563_/A reg1_val[2] _07165_/A vssd1 vssd1 vccd1 vccd1 _07104_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_31_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07034_ _07049_/C _07034_/B vssd1 vssd1 vccd1 vccd1 _07034_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_43_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08985_ _08986_/B _08986_/A vssd1 vssd1 vccd1 vccd1 _08985_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__07337__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07936_ _07936_/A _07936_/B vssd1 vssd1 vccd1 vccd1 _07937_/C sky130_fd_sc_hd__nand2_1
X_07867_ _08775_/A _07867_/B vssd1 vssd1 vccd1 vccd1 _07872_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_98_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10512__C1 _12487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12389__S _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06895__B _06897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11855__A2 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07798_ _07798_/A _07798_/B vssd1 vssd1 vccd1 vccd1 _07801_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_97_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06818_ _11289_/A _06816_/Y _06817_/Y vssd1 vssd1 vccd1 vccd1 _06818_/X sky130_fd_sc_hd__o21a_1
X_09606_ _09606_/A _09606_/B vssd1 vssd1 vccd1 vccd1 _09637_/A sky130_fd_sc_hd__xnor2_2
X_06749_ reg1_val[6] _06996_/A vssd1 vssd1 vccd1 vccd1 _06750_/B sky130_fd_sc_hd__nand2_1
X_09537_ _09535_/Y _09537_/B vssd1 vssd1 vccd1 vccd1 _09538_/B sky130_fd_sc_hd__and2b_1
XANTENNA__07072__A _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07800__A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09468_ _09621_/A _09469_/B vssd1 vssd1 vccd1 vccd1 _09468_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout28_A _07098_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12418__A _12588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08419_ _08419_/A _08419_/B vssd1 vssd1 vccd1 vccd1 _08433_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09399_ _10400_/S _09222_/X _09223_/Y _09398_/X vssd1 vssd1 vccd1 vccd1 dest_val[1]
+ sky130_fd_sc_hd__a31o_4
XANTENNA__08236__B2 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08236__A1 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11430_ _07308_/B fanout9/X _11429_/X _10559_/A vssd1 vssd1 vccd1 vccd1 _11509_/A
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_73_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11361_ _11362_/B _11362_/A vssd1 vssd1 vccd1 vccd1 _11361_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11041__B _11041_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13100_ hold294/X _13151_/A2 _13099_/X _13146_/B2 vssd1 vssd1 vccd1 vccd1 _13101_/B
+ sky130_fd_sc_hd__a22o_1
X_10312_ _10312_/A _10312_/B vssd1 vssd1 vccd1 vccd1 _10325_/A sky130_fd_sc_hd__xor2_1
X_11292_ reg1_val[16] curr_PC[16] vssd1 vssd1 vccd1 vccd1 _11293_/B sky130_fd_sc_hd__nand2_1
X_13031_ hold279/A _13030_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13031_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10372__S _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ _06866_/D _10241_/X _10242_/Y vssd1 vssd1 vccd1 vccd1 _10269_/C sky130_fd_sc_hd__o21a_1
XANTENNA__07211__A2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07247__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10174_ _10174_/A _10174_/B vssd1 vssd1 vccd1 vccd1 _10175_/B sky130_fd_sc_hd__xnor2_2
Xfanout192 _06892_/Y vssd1 vssd1 vccd1 vccd1 _13170_/B sky130_fd_sc_hd__buf_4
Xfanout181 _12788_/B vssd1 vssd1 vccd1 vccd1 _12744_/B sky130_fd_sc_hd__buf_4
Xfanout170 _07047_/X vssd1 vssd1 vccd1 vccd1 _08532_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__08172__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08078__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12815_ hold272/X hold54/X vssd1 vssd1 vccd1 vccd1 _13067_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_97_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12746_ hold54/X _12788_/B vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__or2_1
XANTENNA__07710__A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08475__B2 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08475__A1 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10821__A3 _07435_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12677_ _12682_/A _12677_/B vssd1 vssd1 vccd1 vccd1 _12681_/A sky130_fd_sc_hd__nand2_2
XANTENNA__10282__A1 _10281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11628_ _11629_/B _11629_/A vssd1 vssd1 vccd1 vccd1 _11722_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10034__A1 _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__B1 _08692_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11559_ _11559_/A _11559_/B _11559_/C vssd1 vssd1 vccd1 vccd1 _11559_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09637__A _09637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13229_ _13241_/CLK hold197/X vssd1 vssd1 vccd1 vccd1 hold195/A sky130_fd_sc_hd__dfxtp_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09727__A1 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09727__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07157__A _07157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08770_ _08768_/Y _08770_/B vssd1 vssd1 vccd1 vccd1 _08785_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__06961__A1 _09392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09372__A _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11298__B1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07721_ _07722_/A _07722_/B vssd1 vssd1 vccd1 vccd1 _07721_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07652_ _08942_/B _08942_/A vssd1 vssd1 vccd1 vccd1 _07652_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06603_ reg1_val[24] _07126_/B vssd1 vssd1 vccd1 vccd1 _06603_/X sky130_fd_sc_hd__and2b_1
X_07583_ _07583_/A _07583_/B vssd1 vssd1 vccd1 vccd1 _07588_/A sky130_fd_sc_hd__and2_2
X_06534_ hold47/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__inv_2
XFILLER_0_88_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09322_ _07612_/A _07612_/B _07610_/Y vssd1 vssd1 vccd1 vccd1 _09323_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_87_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout232_A _09384_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09253_ _09253_/A _12087_/A vssd1 vssd1 vccd1 vccd1 _09255_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08204_ _08260_/A _08260_/B _08202_/A vssd1 vssd1 vccd1 vccd1 _08213_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_106_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09184_ _11823_/S _09184_/B vssd1 vssd1 vccd1 vccd1 _09184_/X sky130_fd_sc_hd__or2_4
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08135_ _08836_/A _08199_/A _08199_/B vssd1 vssd1 vccd1 vccd1 _08146_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08066_ _08066_/A _08066_/B vssd1 vssd1 vccd1 vccd1 _08633_/A sky130_fd_sc_hd__xor2_4
XANTENNA__08451__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11288__S _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07017_ _07175_/A _07175_/B _07175_/C vssd1 vssd1 vccd1 vccd1 _07051_/A sky130_fd_sc_hd__or3_1
XANTENNA__07729__B1 _07325_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10328__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08968_ _08954_/A _08954_/B _08952_/X vssd1 vssd1 vccd1 vccd1 _08970_/A sky130_fd_sc_hd__a21o_1
X_07919_ _07919_/A _07919_/B vssd1 vssd1 vccd1 vccd1 _08034_/B sky130_fd_sc_hd__xor2_2
X_08899_ _08899_/A _08899_/B _08899_/C vssd1 vssd1 vccd1 vccd1 _08900_/B sky130_fd_sc_hd__and3_1
XFILLER_0_98_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11317__A _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10930_ _10930_/A _10930_/B vssd1 vssd1 vccd1 vccd1 _10931_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07901__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10861_ _10743_/A _10741_/Y _06722_/B vssd1 vssd1 vccd1 vccd1 _10861_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _12600_/A _12600_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[8] sky130_fd_sc_hd__xor2_4
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ _10793_/A _10793_/B vssd1 vssd1 vccd1 vccd1 _10934_/C sky130_fd_sc_hd__nand2_1
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ _12518_/Y _12539_/C _12541_/B vssd1 vssd1 vccd1 vccd1 _12532_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_54_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12462_ _12471_/A _12462_/B vssd1 vssd1 vccd1 vccd1 _12464_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_47_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11413_ _12022_/A _11413_/B vssd1 vssd1 vccd1 vccd1 _11414_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12393_ _12394_/A _12394_/B _12394_/C vssd1 vssd1 vccd1 vccd1 _12401_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07432__A2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11344_ _12200_/A _11344_/B vssd1 vssd1 vccd1 vccd1 _11350_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09457__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09709__A1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11275_ _11275_/A _11275_/B vssd1 vssd1 vccd1 vccd1 _11460_/A sky130_fd_sc_hd__or2_1
X_13014_ _07097_/B _13020_/B2 hold143/X vssd1 vssd1 vccd1 vccd1 _13277_/D sky130_fd_sc_hd__o21a_1
X_10226_ _10227_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10226_/X sky130_fd_sc_hd__and2_1
XANTENNA__07196__A1 _07303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08393__B1 _07325_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_max_cap128_A _07894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09904__B _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ _10458_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _10158_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10088_ _10088_/A _10088_/B vssd1 vssd1 vccd1 vccd1 _10090_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07499__A2 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09893__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08448__B2 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08448__A1 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12729_ _09283_/A _13020_/B2 hold46/X _13066_/A vssd1 vssd1 vccd1 vccd1 _13186_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07120__A1 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07120__B2 _07119_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10007__B2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10007__A1 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07959__B1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10558__A2 _07308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09940_ _09940_/A _09940_/B vssd1 vssd1 vccd1 vccd1 _09954_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_111_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10306__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09871_ _08680_/B _07197_/Y fanout83/X fanout30/X vssd1 vssd1 vccd1 vccd1 _09872_/B
+ sky130_fd_sc_hd__o22a_1
X_08822_ _12143_/A _08822_/B vssd1 vssd1 vccd1 vccd1 _08824_/B sky130_fd_sc_hd__xnor2_2
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _08864_/B _08752_/C _08752_/A vssd1 vssd1 vccd1 vccd1 _08754_/C sky130_fd_sc_hd__a21o_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout182_A _12742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07704_ _08992_/A _08992_/B _07623_/X vssd1 vssd1 vccd1 vccd1 _07707_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__11137__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08684_ _08683_/B _08683_/C _10015_/A vssd1 vssd1 vccd1 vccd1 _08685_/C sky130_fd_sc_hd__a21o_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07635_ _08837_/B2 _07322_/A _07322_/B fanout46/X _08841_/B2 vssd1 vssd1 vccd1 vccd1
+ _07636_/B sky130_fd_sc_hd__o32a_1
XANTENNA__08439__B2 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08439__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11038__A3 _07435_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07566_ _07566_/A _07566_/B vssd1 vssd1 vccd1 vccd1 _07576_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_91_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09305_ _10565_/A _09305_/B vssd1 vssd1 vccd1 vccd1 _09306_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09976__S _10249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09236_ _09236_/A _09236_/B vssd1 vssd1 vccd1 vccd1 _09237_/B sky130_fd_sc_hd__nand2_1
X_07497_ _10452_/B2 fanout77/X fanout75/X _10527_/A vssd1 vssd1 vccd1 vccd1 _07498_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_90_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09167_ _09165_/X _09166_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09167_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_50_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08118_ _08118_/A _08118_/B vssd1 vssd1 vccd1 vccd1 _08635_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_114_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08181__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09098_ _09098_/A _09103_/A _09103_/B _09102_/A vssd1 vssd1 vccd1 vccd1 _09098_/X
+ sky130_fd_sc_hd__or4b_2
X_08049_ _11499_/A _08109_/B _08109_/A vssd1 vssd1 vccd1 vccd1 _08105_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_102_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout95_A _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11060_ _11060_/A _11060_/B vssd1 vssd1 vccd1 vccd1 _11062_/B sky130_fd_sc_hd__xnor2_1
X_10011_ _10012_/A _10012_/B vssd1 vssd1 vccd1 vccd1 _10013_/A sky130_fd_sc_hd__and2_1
XFILLER_0_98_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12150__B _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09740__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11962_ _12036_/B _11962_/B vssd1 vssd1 vccd1 vccd1 _11964_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06689__B1 _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11682__B1 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913_ _12150_/A _10557_/B fanout13/X _12150_/B vssd1 vssd1 vccd1 vccd1 _10914_/B
+ sky130_fd_sc_hd__o22a_1
X_11893_ _11893_/A _11894_/B vssd1 vssd1 vccd1 vccd1 _11893_/Y sky130_fd_sc_hd__nor2_1
X_10844_ _10725_/A _10725_/B _10723_/X vssd1 vssd1 vccd1 vccd1 _10847_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12514_ _12514_/A _12514_/B vssd1 vssd1 vccd1 vccd1 _12529_/A sky130_fd_sc_hd__nand2_2
X_10775_ _11000_/A _11316_/A _12278_/A vssd1 vssd1 vccd1 vccd1 _10776_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12445_ reg1_val[10] curr_PC[10] _12524_/S vssd1 vssd1 vccd1 vccd1 _12447_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_41_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12376_ _12353_/Y _12354_/X _12357_/Y _09192_/Y _12375_/X vssd1 vssd1 vccd1 vccd1
+ _12376_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_2_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11327_ _11327_/A _11327_/B vssd1 vssd1 vccd1 vccd1 _11328_/C sky130_fd_sc_hd__xor2_1
X_11258_ _11145_/B _11152_/B _11143_/Y vssd1 vssd1 vccd1 vccd1 _11268_/A sky130_fd_sc_hd__a21oi_1
X_11189_ reg1_val[15] curr_PC[15] vssd1 vssd1 vccd1 vccd1 _11191_/A sky130_fd_sc_hd__nand2_1
X_10209_ _10209_/A _10209_/B vssd1 vssd1 vccd1 vccd1 _10223_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_82_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09866__B1 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12487__S _12487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09618__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07420_ _07420_/A _07420_/B vssd1 vssd1 vccd1 vccd1 _07424_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08266__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07351_ _07349_/A _07349_/B _07350_/X vssd1 vssd1 vccd1 vccd1 _07353_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_18_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07644__A2 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08841__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08841__B2 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07282_ _07591_/A _07282_/B vssd1 vssd1 vccd1 vccd1 _07295_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09021_ _09020_/A _09020_/B _08256_/Y _08257_/X _09063_/A vssd1 vssd1 vccd1 vccd1
+ _09022_/B sky130_fd_sc_hd__a2111o_1
XFILLER_0_60_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12925__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11420__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 hold234/A vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold212 hold212/A vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 hold278/A vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 hold245/A vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 hold267/A vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 hold256/A vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_13_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold289 hold289/A vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ fanout75/X _08134_/B fanout51/X _10553_/B vssd1 vssd1 vccd1 vccd1 _09924_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09854_ _09158_/S _12181_/B _09835_/X _09837_/A _09853_/Y vssd1 vssd1 vccd1 vccd1
+ _09854_/X sky130_fd_sc_hd__a221o_1
XANTENNA__10164__B1 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _08805_/A _08805_/B vssd1 vssd1 vccd1 vccd1 _08806_/C sky130_fd_sc_hd__xor2_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06997_ reg1_val[24] _06997_/B vssd1 vssd1 vccd1 vccd1 _07005_/C sky130_fd_sc_hd__xnor2_4
X_09785_ _11134_/B2 fanout46/X fanout12/X _07179_/Y vssd1 vssd1 vccd1 vccd1 _09786_/B
+ sky130_fd_sc_hd__o22a_1
X_08736_ _08217_/B fanout82/X _08672_/B fanout55/X vssd1 vssd1 vccd1 vccd1 _08737_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08667_ _08667_/A _08667_/B vssd1 vssd1 vccd1 vccd1 _08689_/A sky130_fd_sc_hd__xor2_2
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ _07619_/A _07619_/B vssd1 vssd1 vccd1 vccd1 _07618_/X sky130_fd_sc_hd__and2_1
XANTENNA__09609__B1 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08176__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08598_ _08589_/A _08592_/A _08598_/S vssd1 vssd1 vccd1 vccd1 _08599_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_64_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07549_ _07549_/A _07549_/B vssd1 vssd1 vccd1 vccd1 _07599_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_119_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07635__A2 _07322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10560_ _10559_/B _10559_/C _10559_/A vssd1 vssd1 vccd1 vccd1 _10562_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12426__A _12593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ _12726_/A _12250_/B _06930_/Y _09218_/X vssd1 vssd1 vccd1 vccd1 _09219_/X
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10491_ _10730_/A _10491_/B vssd1 vssd1 vccd1 vccd1 _10524_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09388__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12230_ _12230_/A _12230_/B vssd1 vssd1 vccd1 vccd1 _12230_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12161_ _12161_/A _12161_/B vssd1 vssd1 vccd1 vccd1 _12215_/B sky130_fd_sc_hd__nor2_1
X_11112_ _12019_/A _11112_/B vssd1 vssd1 vccd1 vccd1 _11116_/A sky130_fd_sc_hd__xnor2_1
X_12092_ _12027_/A _12027_/B _12026_/A vssd1 vssd1 vccd1 vccd1 _12094_/B sky130_fd_sc_hd__a21oi_1
X_11043_ _11044_/B _11044_/A vssd1 vssd1 vccd1 vccd1 _11043_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_36_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07571__B2 _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__A1 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12994_ _11429_/B _13020_/B2 hold117/X vssd1 vssd1 vccd1 vccd1 _13267_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_99_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11945_ _12022_/A _11945_/B vssd1 vssd1 vccd1 vccd1 _11947_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11876_ _11952_/B _11876_/B vssd1 vssd1 vccd1 vccd1 _11878_/C sky130_fd_sc_hd__or2_1
X_10827_ _10827_/A _10827_/B vssd1 vssd1 vccd1 vccd1 _10842_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_125_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10758_ hold301/A _10758_/B vssd1 vssd1 vccd1 vccd1 _10877_/B sky130_fd_sc_hd__or2_1
XFILLER_0_109_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12428_ _12429_/A _12429_/B _12429_/C vssd1 vssd1 vccd1 vccd1 _12436_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_35_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11240__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10689_ _10927_/A _07278_/B fanout83/X fanout6/X vssd1 vssd1 vccd1 vccd1 _10690_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_77_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12359_ _12360_/A _12360_/B vssd1 vssd1 vccd1 vccd1 _12359_/X sky130_fd_sc_hd__or2_1
XFILLER_0_22_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06920_ instruction[3] instruction[6] instruction[5] instruction[4] vssd1 vssd1 vccd1
+ vccd1 _09184_/B sky130_fd_sc_hd__or4b_4
XANTENNA__12135__A1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06988__B _11695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ _12045_/A _06850_/X _06839_/X vssd1 vssd1 vccd1 vccd1 _06851_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_89_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06782_ _12563_/A _09392_/S vssd1 vssd1 vccd1 vccd1 _09383_/A sky130_fd_sc_hd__xnor2_2
X_09570_ _09570_/A _09570_/B vssd1 vssd1 vccd1 vccd1 _09573_/A sky130_fd_sc_hd__nand2_1
X_08521_ _08521_/A _08531_/A vssd1 vssd1 vccd1 vccd1 _08522_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08452_ _08487_/A _08487_/B vssd1 vssd1 vccd1 vccd1 _08488_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07314__B2 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07314__A1 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07403_ _07629_/A _07401_/A _07678_/A _07402_/X vssd1 vssd1 vccd1 vccd1 _07414_/B
+ sky130_fd_sc_hd__a31o_1
X_08383_ _08383_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _08418_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08724__A _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ _10169_/A _07334_/B vssd1 vssd1 vccd1 vccd1 _07335_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07265_ _07266_/B _07265_/B vssd1 vssd1 vccd1 vccd1 _07267_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09004_ _08018_/Y _09029_/B _08806_/X vssd1 vssd1 vccd1 vccd1 _09031_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_103_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12374__A1 _09200_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07196_ _07303_/A _07303_/C _07303_/B vssd1 vssd1 vccd1 vccd1 _07197_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08578__B1 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11582__C1 _11557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__A2 _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10924__A2 _10925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12126__B2 _06928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09906_ _10658_/A _09906_/B _09906_/C vssd1 vssd1 vccd1 vccd1 _09909_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10137__B1 _12345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09837_ _09837_/A vssd1 vssd1 vccd1 vccd1 _09837_/Y sky130_fd_sc_hd__inv_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ _09879_/A _09768_/B vssd1 vssd1 vccd1 vccd1 _09770_/B sky130_fd_sc_hd__or2_1
XFILLER_0_96_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08719_ _08009_/A _08009_/B _08010_/Y vssd1 vssd1 vccd1 vccd1 _08805_/A sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout58_A _07157_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11101__A2 wire201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09699_ hold237/A _09698_/X _12290_/C1 vssd1 vssd1 vccd1 vccd1 _09699_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ _11730_/A _11730_/B _11730_/C _11730_/D vssd1 vssd1 vccd1 vccd1 _11731_/B
+ sky130_fd_sc_hd__or4_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ reg1_val[20] _06653_/B _11660_/X vssd1 vssd1 vccd1 vccd1 _11661_/Y sky130_fd_sc_hd__o21ai_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12062__B1 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10612_ _10098_/X _10608_/Y _10609_/Y _09511_/B _10611_/Y vssd1 vssd1 vccd1 vccd1
+ _10613_/B sky130_fd_sc_hd__o221ai_4
X_11592_ fanout32/X _12203_/A _12150_/A fanout29/X vssd1 vssd1 vccd1 vccd1 _11593_/B
+ sky130_fd_sc_hd__o22a_1
X_10543_ _10544_/B _10543_/B vssd1 vssd1 vccd1 vccd1 _10662_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_24_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10612__B2 _09511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08353__B _10551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13262_ _13280_/CLK _13262_/D vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13011__C1 _13028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10474_ _10475_/A _10475_/B vssd1 vssd1 vccd1 vccd1 _10474_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13193_ _13289_/CLK _13193_/D vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfxtp_1
X_12213_ _12213_/A _12213_/B _12213_/C vssd1 vssd1 vccd1 vccd1 _12214_/B sky130_fd_sc_hd__or3_1
XANTENNA__09230__B2 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09230__A1 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07241__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12144_ _12144_/A _12144_/B vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__and2_1
XANTENNA__07792__B2 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07792__A1 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12603__B _12603_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12075_ _12023_/A _12023_/B _12020_/A vssd1 vssd1 vccd1 vccd1 _12083_/A sky130_fd_sc_hd__a21o_1
X_11026_ _12150_/B fanout47/X _11603_/A _12776_/A vssd1 vssd1 vccd1 vccd1 _11027_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA_max_cap110_A _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07713__A _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12977_ hold140/X _12723_/A _13170_/B hold144/X _13066_/A vssd1 vssd1 vccd1 vccd1
+ hold145/A sky130_fd_sc_hd__o221a_1
XFILLER_0_87_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11928_ curr_PC[21] curr_PC[22] _11764_/B curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11928_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10300__B1 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11859_ _11938_/B _11859_/B vssd1 vssd1 vccd1 vccd1 _11861_/B sky130_fd_sc_hd__or2_1
XFILLER_0_55_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_18 reg1_val[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_29 reg1_val[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07050_ _07050_/A _07050_/B _07050_/C vssd1 vssd1 vccd1 vccd1 _07128_/B sky130_fd_sc_hd__and3_2
XFILLER_0_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09221__A1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10367__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09375__A _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07952_ _08841_/B2 _08134_/B fanout51/X _09888_/B2 vssd1 vssd1 vccd1 vccd1 _07953_/B
+ sky130_fd_sc_hd__o22a_1
X_06903_ instruction[15] _06904_/B vssd1 vssd1 vccd1 vccd1 dest_idx[4] sky130_fd_sc_hd__and2_4
X_07883_ _07883_/A _07883_/B vssd1 vssd1 vccd1 vccd1 _07885_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07535__A1 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__B1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06834_ reg1_val[30] _06834_/B vssd1 vssd1 vccd1 vccd1 _06834_/Y sky130_fd_sc_hd__nand2_1
X_09622_ _09622_/A _09622_/B vssd1 vssd1 vccd1 vccd1 _09634_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__07535__B2 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11331__A2 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09553_ _10249_/S _12250_/B _09191_/X _09694_/A _09550_/X vssd1 vssd1 vccd1 vccd1
+ _09553_/X sky130_fd_sc_hd__o221a_1
XANTENNA_fanout262_A _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08504_ _08505_/A _08505_/B vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__or2_1
X_06765_ reg2_val[3] _06778_/B vssd1 vssd1 vccd1 vccd1 _06765_/X sky130_fd_sc_hd__and2_1
X_06696_ reg1_val[15] _07178_/A vssd1 vssd1 vccd1 vccd1 _06696_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12292__B1 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09484_ _09484_/A _09484_/B vssd1 vssd1 vccd1 vccd1 _09485_/B sky130_fd_sc_hd__xor2_1
X_08435_ _08435_/A _08435_/B vssd1 vssd1 vccd1 vccd1 _08484_/A sky130_fd_sc_hd__xnor2_1
X_08366_ _08373_/A _08373_/B _08351_/X vssd1 vssd1 vccd1 vccd1 _08403_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_92_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07317_ _09580_/A _07317_/B vssd1 vssd1 vccd1 vccd1 _07852_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_34_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08297_ _08297_/A _08297_/B vssd1 vssd1 vccd1 vccd1 _08298_/B sky130_fd_sc_hd__or2_1
XFILLER_0_46_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07248_ _07249_/A _07249_/B vssd1 vssd1 vccd1 vccd1 _07248_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07179_ _07179_/A vssd1 vssd1 vccd1 vccd1 _07179_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_42_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10190_ _10190_/A _10190_/B vssd1 vssd1 vccd1 vccd1 _10192_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08723__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12900_ _13169_/A hold218/X vssd1 vssd1 vccd1 vccd1 _13220_/D sky130_fd_sc_hd__and2_1
XANTENNA__11322__A2 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12831_ hold38/X hold36/X vssd1 vssd1 vccd1 vccd1 _13025_/B sky130_fd_sc_hd__nand2b_1
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13075__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08348__B _08348_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12762_/A _12778_/B vssd1 vssd1 vccd1 vccd1 _12762_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12283__B1 _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12693_ _12693_/A _12698_/C vssd1 vssd1 vccd1 vccd1 loadstore_address[27] sky130_fd_sc_hd__xnor2_4
XANTENNA__10894__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11713_ _11713_/A _11713_/B vssd1 vssd1 vccd1 vccd1 _11715_/B sky130_fd_sc_hd__xnor2_1
X_11644_ _12332_/B _09069_/A _09073_/C vssd1 vssd1 vccd1 vccd1 _11644_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11575_ _13236_/Q _11559_/A _11751_/C _11920_/C1 vssd1 vssd1 vccd1 vccd1 _11575_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09451__B2 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09451__A1 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13314_ _13318_/CLK hold172/X vssd1 vssd1 vccd1 vccd1 hold298/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10526_ _10477_/A _10477_/B _10478_/X vssd1 vssd1 vccd1 vccd1 _10603_/A sky130_fd_sc_hd__a21o_2
X_13245_ _13312_/CLK _13245_/D vssd1 vssd1 vccd1 vccd1 hold165/A sky130_fd_sc_hd__dfxtp_1
X_10457_ _10458_/B _10458_/A vssd1 vssd1 vccd1 vccd1 _10457_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07708__A _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07214__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11010__A1 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ _13179_/A _13176_/B hold299/X vssd1 vssd1 vccd1 vccd1 hold300/A sky130_fd_sc_hd__and3_1
X_10388_ _10266_/A _10263_/Y _10265_/B vssd1 vssd1 vccd1 vccd1 _10392_/A sky130_fd_sc_hd__o21a_1
XANTENNA__11010__B2 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _06617_/Y wire201/X _12125_/X _06619_/B _12126_/X vssd1 vssd1 vccd1 vccd1
+ _12127_/X sky130_fd_sc_hd__a221o_1
X_12058_ hold286/A _12119_/B1 _12183_/C _12057_/Y _11400_/A vssd1 vssd1 vccd1 vccd1
+ _12058_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_74_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11009_ _12349_/B _11009_/B vssd1 vssd1 vccd1 vccd1 _11017_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06689__A2_N _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07443__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06550_ instruction[0] instruction[1] instruction[2] pred_val vssd1 vssd1 vccd1 vccd1
+ _06550_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_75_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08220_ _08774_/A2 _08672_/B _08835_/B1 _08774_/B1 vssd1 vssd1 vccd1 vccd1 _08221_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08274__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08151_ _08151_/A _08151_/B vssd1 vssd1 vccd1 vccd1 _08153_/B sky130_fd_sc_hd__and2_1
XFILLER_0_43_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08082_ _08774_/A2 _12752_/A fanout84/X _08774_/B1 vssd1 vssd1 vccd1 vccd1 _08083_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09993__A2 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06627__A2_N _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07102_ _07162_/A _07162_/B vssd1 vssd1 vccd1 vccd1 _07164_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_43_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07453__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07033_ _07167_/A _07050_/A _07050_/B _07135_/B vssd1 vssd1 vccd1 vccd1 _07034_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout108_A _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08984_ _08984_/A _08984_/B vssd1 vssd1 vccd1 vccd1 _08986_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07935_ _07935_/A _07935_/B _07935_/C vssd1 vssd1 vccd1 vccd1 _07936_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07866_ _08572_/B _11147_/A _11012_/A _07117_/Y vssd1 vssd1 vccd1 vccd1 _07867_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10512__B1 _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08449__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09605_ _09605_/A _09605_/B vssd1 vssd1 vccd1 vccd1 _09606_/B sky130_fd_sc_hd__xnor2_2
X_07797_ _07797_/A _07797_/B vssd1 vssd1 vccd1 vccd1 _07798_/B sky130_fd_sc_hd__nor2_1
X_06817_ reg1_val[16] _07167_/A vssd1 vssd1 vccd1 vccd1 _06817_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06748_ reg1_val[6] _06996_/A vssd1 vssd1 vccd1 vccd1 _06748_/X sky130_fd_sc_hd__and2_1
X_09536_ reg1_val[2] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09537_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07072__B _07080_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09467_ _09467_/A _09467_/B vssd1 vssd1 vccd1 vccd1 _09469_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08418_ _08418_/A _08418_/B vssd1 vssd1 vccd1 vccd1 _08419_/B sky130_fd_sc_hd__xnor2_1
X_06679_ _06687_/A _12568_/B vssd1 vssd1 vccd1 vccd1 _06679_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_65_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11603__A _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09398_ _09336_/Y _09340_/X _09376_/X _09397_/X _12382_/S vssd1 vssd1 vccd1 vccd1
+ _09398_/X sky130_fd_sc_hd__o41a_1
XFILLER_0_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08236__A2 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08349_ _08853_/A _08385_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _08365_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11360_ _11360_/A _11360_/B vssd1 vssd1 vccd1 vccd1 _11362_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07444__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10311_ _10311_/A _10311_/B vssd1 vssd1 vccd1 vccd1 _10312_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13030_ _13030_/A _13030_/B vssd1 vssd1 vccd1 vccd1 _13030_/Y sky130_fd_sc_hd__xnor2_1
X_11291_ reg1_val[16] curr_PC[16] vssd1 vssd1 vccd1 vccd1 _11291_/Y sky130_fd_sc_hd__nor2_1
X_10242_ _06866_/D _10241_/X _12277_/B1 vssd1 vssd1 vccd1 vccd1 _10242_/Y sky130_fd_sc_hd__a21oi_1
X_10173_ _10174_/A _10174_/B vssd1 vssd1 vccd1 vccd1 _10173_/X sky130_fd_sc_hd__or2_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout182 _12742_/B vssd1 vssd1 vccd1 vccd1 _12788_/B sky130_fd_sc_hd__buf_4
Xfanout171 _07047_/X vssd1 vssd1 vccd1 vccd1 _08772_/B2 sky130_fd_sc_hd__buf_4
Xfanout160 _07154_/X vssd1 vssd1 vccd1 vccd1 _09273_/A1 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08172__A1 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08172__B2 _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout193 _13168_/B1 vssd1 vssd1 vccd1 vccd1 _12947_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_88_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12814_ hold276/X hold81/X vssd1 vssd1 vccd1 vccd1 _13072_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12745_ _07325_/Y _12980_/A2 hold64/X _13179_/A vssd1 vssd1 vccd1 vccd1 _13194_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_97_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08475__A2 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08094__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06607__A _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ reg1_val[24] _12708_/B vssd1 vssd1 vccd1 vccd1 _12677_/B sky130_fd_sc_hd__or2_1
XANTENNA__10282__A2 _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12008__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11627_ _11722_/A _11627_/B vssd1 vssd1 vccd1 vccd1 _11629_/B sky130_fd_sc_hd__or2_1
XFILLER_0_114_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11558_ _12332_/B _11559_/B _11559_/C vssd1 vssd1 vccd1 vccd1 _11558_/X sky130_fd_sc_hd__a21o_1
XANTENNA__07435__B1 _06622_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07986__B2 _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07986__A1 _12768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10509_ hold187/A _13224_/Q _10509_/C vssd1 vssd1 vccd1 vccd1 _10632_/B sky130_fd_sc_hd__or3_1
XANTENNA__08822__A _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10990__B1 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11489_ _09115_/X _10981_/Y _10992_/Y _09184_/X _11488_/X vssd1 vssd1 vccd1 vccd1
+ _11490_/C sky130_fd_sc_hd__o221a_1
X_13228_ _13243_/CLK _13228_/D vssd1 vssd1 vccd1 vccd1 hold219/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07438__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09727__A2 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13159_ hold270/A _13158_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13159_/X sky130_fd_sc_hd__mux2_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ _08773_/A _07720_/B vssd1 vssd1 vccd1 vccd1 _07722_/B sky130_fd_sc_hd__xor2_2
XANTENNA__06961__A2 _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10799__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_07651_ _07651_/A _07651_/B vssd1 vssd1 vccd1 vccd1 _08942_/B sky130_fd_sc_hd__xor2_1
X_06602_ _07126_/B reg1_val[24] vssd1 vssd1 vccd1 vccd1 _06602_/Y sky130_fd_sc_hd__nand2b_2
X_07582_ _07582_/A _07582_/B vssd1 vssd1 vccd1 vccd1 _07583_/B sky130_fd_sc_hd__or2_1
X_06533_ hold296/X vssd1 vssd1 vccd1 vccd1 _06533_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_87_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09321_ _09321_/A _09321_/B vssd1 vssd1 vccd1 vccd1 _09323_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__13114__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09663__A1 _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09252_ _09252_/A _09252_/B vssd1 vssd1 vccd1 vccd1 _09255_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08203_ _08203_/A _08203_/B vssd1 vssd1 vccd1 vccd1 _08260_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_105_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09183_ _11823_/S _09184_/B vssd1 vssd1 vccd1 vccd1 _09183_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08134_ _08821_/A _08134_/B vssd1 vssd1 vccd1 vccd1 _08199_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_71_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12970__A1 _07046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08065_ _08018_/Y _08064_/Y _08017_/X vssd1 vssd1 vccd1 vccd1 _08065_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07729__A1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07016_ _07175_/A _07175_/B _07175_/C vssd1 vssd1 vccd1 vccd1 _07050_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_101_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07729__B2 _07182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ _08946_/A _08946_/B _08945_/A vssd1 vssd1 vccd1 vccd1 _08972_/A sky130_fd_sc_hd__o21ai_2
X_07918_ _08034_/A vssd1 vssd1 vccd1 vccd1 _07918_/Y sky130_fd_sc_hd__inv_2
X_08898_ _08899_/A _08899_/B _08899_/C vssd1 vssd1 vccd1 vccd1 _08950_/A sky130_fd_sc_hd__a21oi_1
X_07849_ _07848_/B _07848_/C _07848_/A vssd1 vssd1 vccd1 vccd1 _07880_/A sky130_fd_sc_hd__o21ba_2
XANTENNA__07083__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07901__A1 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07901__B2 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ _11381_/A _10860_/B vssd1 vssd1 vccd1 vccd1 _10860_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07811__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12789__A1 _07435_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09519_ _11195_/A _09518_/Y _09214_/A vssd1 vssd1 vccd1 vccd1 _12284_/B sky130_fd_sc_hd__o21a_1
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12334__A2_N wire201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10791_ _11499_/A _10791_/B vssd1 vssd1 vccd1 vccd1 _10793_/B sky130_fd_sc_hd__xnor2_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ _12530_/A vssd1 vssd1 vccd1 vccd1 _12539_/C sky130_fd_sc_hd__inv_2
XFILLER_0_109_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12461_ _12620_/B _12461_/B vssd1 vssd1 vccd1 vccd1 _12462_/B sky130_fd_sc_hd__or2_1
XFILLER_0_47_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11412_ fanout37/X _11935_/A _12772_/A fanout35/X vssd1 vssd1 vccd1 vccd1 _11413_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12392_ _12401_/A _12392_/B vssd1 vssd1 vccd1 vccd1 _12394_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11343_ fanout70/X fanout15/X fanout6/X _11431_/A vssd1 vssd1 vccd1 vccd1 _11344_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07258__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11274_ _11274_/A _11274_/B _11274_/C vssd1 vssd1 vccd1 vccd1 _11275_/B sky130_fd_sc_hd__nor3_1
X_13013_ hold92/X _13013_/A2 _13020_/A2 hold51/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold143/A sky130_fd_sc_hd__o221a_1
X_10225_ _10227_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10225_/X sky130_fd_sc_hd__or2_1
XANTENNA__08393__A1 _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08393__B2 _08544_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ _10156_/A1 fanout18/X fanout9/X _10156_/B2 vssd1 vssd1 vccd1 vccd1 _10157_/B
+ sky130_fd_sc_hd__o22a_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11508__A _11509_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10087_ _10088_/B _10088_/A vssd1 vssd1 vccd1 vccd1 _10087_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_89_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09893__A1 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09893__B2 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10989_ _07197_/A _06928_/X _11099_/B reg1_val[13] vssd1 vssd1 vccd1 vccd1 _10989_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08448__A2 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12728_ hold45/X _12744_/B vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__or2_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07656__B1 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07120__A2 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12659_ _12660_/B _12660_/C _12678_/A vssd1 vssd1 vccd1 vccd1 _12661_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_5_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10007__A2 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07959__A1 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11755__A2 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07959__B2 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09870_ _09870_/A _09870_/B vssd1 vssd1 vccd1 vccd1 _09873_/A sky130_fd_sc_hd__nor2_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _08821_/A _08821_/B vssd1 vssd1 vccd1 vccd1 _08822_/B sky130_fd_sc_hd__nor2_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09581__B1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13109__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08752_ _08752_/A _08864_/B _08752_/C vssd1 vssd1 vccd1 vccd1 _08754_/B sky130_fd_sc_hd__nand3_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11418__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08683_ _10015_/A _08683_/B _08683_/C vssd1 vssd1 vccd1 vccd1 _08685_/B sky130_fd_sc_hd__nand3_1
X_07703_ _07703_/A _07703_/B vssd1 vssd1 vccd1 vccd1 _08992_/B sky130_fd_sc_hd__xor2_4
XANTENNA_fanout175_A _06963_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07634_ _08836_/A _07634_/B vssd1 vssd1 vccd1 vccd1 _07637_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07895__B1 _07182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08439__A2 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07565_ _10565_/A _07565_/B vssd1 vssd1 vccd1 vccd1 _07566_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09304_ _10927_/A fanout46/X fanout12/X fanout83/X vssd1 vssd1 vccd1 vccd1 _09305_/B
+ sky130_fd_sc_hd__o22a_1
X_07496_ _07496_/A _07496_/B vssd1 vssd1 vccd1 vccd1 _07542_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_118_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09235_ _09236_/A _09236_/B vssd1 vssd1 vccd1 vccd1 _09237_/A sky130_fd_sc_hd__or2_1
XFILLER_0_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09166_ reg1_val[19] reg1_val[12] _09172_/S vssd1 vssd1 vccd1 vccd1 _09166_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08117_ _08633_/A _08633_/B vssd1 vssd1 vccd1 vccd1 _08643_/A sky130_fd_sc_hd__or2_1
XANTENNA__08072__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09097_ _09102_/A _09097_/B vssd1 vssd1 vccd1 vccd1 _12279_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_44_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08048_ _08836_/A _08048_/B vssd1 vssd1 vccd1 vccd1 _08109_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11903__C1 _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout88_A _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10010_ _10565_/A _10010_/B vssd1 vssd1 vccd1 vccd1 _10012_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07806__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ _12005_/A _10138_/B vssd1 vssd1 vccd1 vccd1 _09999_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12150__C _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ _11961_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _11962_/B sky130_fd_sc_hd__nand2_1
X_10912_ _11853_/A _10912_/B vssd1 vssd1 vccd1 vccd1 _10916_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11682__B2 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11682__A1 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11892_ _11892_/A _11967_/A vssd1 vssd1 vccd1 vccd1 _11894_/B sky130_fd_sc_hd__nand2_1
X_10843_ _10843_/A _10843_/B vssd1 vssd1 vccd1 vccd1 _10847_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07638__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10774_ _10774_/A _10774_/B vssd1 vssd1 vccd1 vccd1 _11316_/A sky130_fd_sc_hd__or2_1
X_12513_ _12557_/A _12513_/B vssd1 vssd1 vccd1 vccd1 _12514_/B sky130_fd_sc_hd__or2_1
XFILLER_0_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12444_ _12450_/B _12444_/B vssd1 vssd1 vccd1 vccd1 new_PC[9] sky130_fd_sc_hd__and2_4
XFILLER_0_50_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09468__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12606__B _12607_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12375_ _11381_/A _12359_/X _12360_/Y _12363_/X _12374_/X vssd1 vssd1 vccd1 vccd1
+ _12375_/X sky130_fd_sc_hd__a311o_1
XANTENNA__10407__A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07810__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06604__B _07126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11326_ _11327_/A _11327_/B vssd1 vssd1 vccd1 vccd1 _11444_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11257_ _11257_/A _11257_/B vssd1 vssd1 vccd1 vccd1 _11270_/A sky130_fd_sc_hd__xor2_2
X_11188_ _11187_/A _11187_/B _11187_/Y _12277_/B1 vssd1 vssd1 vccd1 vccd1 _11188_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_66_48 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10208_ _10208_/A _10208_/B vssd1 vssd1 vccd1 vccd1 _10209_/B sky130_fd_sc_hd__xnor2_1
X_10139_ curr_PC[6] _10138_/B _10400_/S vssd1 vssd1 vccd1 vccd1 _10139_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__11238__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09931__A _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11122__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09866__B2 _09295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09866__A1 _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09618__A1 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09618__B2 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07350_ _07421_/B _07421_/A vssd1 vssd1 vccd1 vccd1 _07350_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_9_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11976__A2 _09076_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09020_ _09020_/A _09020_/B vssd1 vssd1 vccd1 vccd1 _09063_/B sky130_fd_sc_hd__and2_2
XFILLER_0_93_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08841__A2 _07301_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07281_ _10280_/A _07281_/B vssd1 vssd1 vccd1 vccd1 _07282_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_122_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold202 hold202/A vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10317__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold235 hold235/A vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 hold213/A vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 hold224/A vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold268 hold268/A vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__buf_1
Xhold257 hold257/A vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 hold246/A vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 hold279/A vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09922_ _09729_/A _09729_/B _09726_/A vssd1 vssd1 vccd1 vccd1 _09936_/A sky130_fd_sc_hd__o21ai_2
X_09853_ _06868_/C _09383_/B _09840_/X _09852_/X vssd1 vssd1 vccd1 vccd1 _09853_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__09554__B1 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10164__A1 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout292_A _13028_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08804_ _08801_/X _08804_/B vssd1 vssd1 vccd1 vccd1 _09032_/A sky130_fd_sc_hd__nand2b_2
X_09784_ _10555_/A _09784_/B vssd1 vssd1 vccd1 vccd1 _09788_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10164__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ _08855_/A _08735_/B vssd1 vssd1 vccd1 vccd1 _08739_/A sky130_fd_sc_hd__xnor2_1
X_06996_ _06996_/A _06996_/B vssd1 vssd1 vccd1 vccd1 _06996_/X sky130_fd_sc_hd__xor2_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11113__B1 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07868__B1 _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08666_ _09580_/A _08666_/B vssd1 vssd1 vccd1 vccd1 _08667_/B sky130_fd_sc_hd__xnor2_2
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08597_ _08597_/A _08597_/B vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__xnor2_1
X_07617_ _07617_/A _07617_/B vssd1 vssd1 vccd1 vccd1 _07619_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__09609__A1 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07080__B _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09609__B2 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07548_ _07548_/A _07548_/B vssd1 vssd1 vccd1 vccd1 _07549_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07635__A3 _07322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07479_ _07479_/A _07479_/B vssd1 vssd1 vccd1 vccd1 _07582_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_106_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08192__A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09218_ _09111_/X _09218_/B _09218_/C _09218_/D vssd1 vssd1 vccd1 vccd1 _09218_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_17_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10490_ _09962_/B _10487_/Y _10961_/B vssd1 vssd1 vccd1 vccd1 _10491_/B sky130_fd_sc_hd__o21ba_1
X_09149_ _09147_/X _09148_/X _09359_/S vssd1 vssd1 vccd1 vccd1 _09149_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12377__C1 _12382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10014__A2_N fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12160_ _12160_/A _12160_/B _12160_/C vssd1 vssd1 vccd1 vccd1 _12161_/B sky130_fd_sc_hd__and3_1
XFILLER_0_31_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11111_ fanout29/X _11794_/A _12772_/A fanout32/X vssd1 vssd1 vccd1 vccd1 _11112_/B
+ sky130_fd_sc_hd__o22a_1
X_12091_ _12160_/A _12091_/B vssd1 vssd1 vccd1 vccd1 _12094_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07536__A _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11042_ _11150_/A _11042_/B vssd1 vssd1 vccd1 vccd1 _11044_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07571__A2 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09751__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12993_ hold113/X _13013_/A2 _13020_/A2 hold116/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold117/A sky130_fd_sc_hd__o221a_1
XFILLER_0_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11944_ fanout35/X fanout19/X _12301_/A fanout37/X vssd1 vssd1 vccd1 vccd1 _11945_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11875_ _11875_/A _11875_/B vssd1 vssd1 vccd1 vccd1 _11876_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10826_ _10826_/A _10826_/B vssd1 vssd1 vccd1 vccd1 _10827_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10757_ hold219/A _12187_/A1 _10874_/B _11920_/C1 vssd1 vssd1 vccd1 vccd1 _10757_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10688_ _10688_/A _10688_/B vssd1 vssd1 vccd1 vccd1 _10698_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08036__B1 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12427_ _12436_/A _12427_/B vssd1 vssd1 vccd1 vccd1 _12429_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10918__B1 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10394__A1 _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10394__B2 _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12358_ _12278_/B _12279_/A _12326_/A _12278_/A vssd1 vssd1 vccd1 vccd1 _12360_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12289_ _12332_/B _12330_/B _13246_/Q vssd1 vssd1 vccd1 vccd1 _12289_/Y sky130_fd_sc_hd__a21oi_1
X_11309_ _11283_/X _11308_/X _12382_/S vssd1 vssd1 vccd1 vccd1 _11309_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_10_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06850_ _06604_/X _06833_/B _06840_/X vssd1 vssd1 vccd1 vccd1 _06850_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11343__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06781_ _12563_/A _09392_/S vssd1 vssd1 vccd1 vccd1 _09544_/A sky130_fd_sc_hd__or2_1
XFILLER_0_26_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08277__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08520_ _08521_/A _08520_/B _08520_/C vssd1 vssd1 vccd1 vccd1 _08531_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08451_ _08777_/A _08451_/B vssd1 vssd1 vccd1 vccd1 _08487_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07314__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07402_ _08588_/A _07389_/B _10280_/A vssd1 vssd1 vccd1 vccd1 _07402_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_92_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08382_ _08773_/A _08382_/B vssd1 vssd1 vccd1 vccd1 _08418_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12071__A1 _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07333_ _08821_/B _09478_/B2 fanout36/X _09476_/A vssd1 vssd1 vccd1 vccd1 _07334_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout138_A _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07264_ _10180_/A _07264_/B vssd1 vssd1 vccd1 vccd1 _07265_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11431__A _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08027__B1 _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09003_ _09968_/A _12357_/A vssd1 vssd1 vccd1 vccd1 _11379_/A sky130_fd_sc_hd__nand2_4
XFILLER_0_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13020__B1 _11147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07195_ _07195_/A _07195_/B vssd1 vssd1 vccd1 vccd1 _07195_/X sky130_fd_sc_hd__and2_2
XANTENNA__08578__A1 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__B2 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10047__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06898__C _06898_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire3 wire3/A vssd1 vssd1 vccd1 vccd1 wire3/X sky130_fd_sc_hd__buf_1
X_09905_ _09906_/B _09906_/C _10658_/A vssd1 vssd1 vccd1 vccd1 _09909_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_6_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09836_ _11197_/S _09851_/B _09183_/Y vssd1 vssd1 vccd1 vccd1 _09837_/A sky130_fd_sc_hd__a21o_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06979_ reg1_val[20] reg1_val[21] _07087_/B _12658_/B _07165_/A vssd1 vssd1 vccd1
+ vccd1 _06980_/B sky130_fd_sc_hd__o41a_2
X_09767_ _09766_/B _09767_/B vssd1 vssd1 vccd1 vccd1 _09768_/B sky130_fd_sc_hd__and2b_1
X_08718_ _08720_/A _08720_/B vssd1 vssd1 vccd1 vccd1 _08801_/A sky130_fd_sc_hd__nand2_1
X_09698_ hold297/A _13218_/Q hold211/A _12124_/B vssd1 vssd1 vccd1 vccd1 _09698_/X
+ sky130_fd_sc_hd__o31a_1
XANTENNA__08187__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08649_ _08650_/A _08650_/B vssd1 vssd1 vccd1 vccd1 _08766_/A sky130_fd_sc_hd__nor2_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07091__A _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11660_ _06654_/A _11838_/A2 _10638_/B vssd1 vssd1 vccd1 vccd1 _11660_/X sky130_fd_sc_hd__a21o_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11591_ _12206_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11595_/A sky130_fd_sc_hd__xnor2_1
X_10611_ _10363_/Y _10850_/A _10610_/Y vssd1 vssd1 vccd1 vccd1 _10611_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13330_ instruction[4] vssd1 vssd1 vccd1 vccd1 sign_extend sky130_fd_sc_hd__buf_12
X_10542_ _12143_/A _10542_/B vssd1 vssd1 vccd1 vccd1 _10543_/B sky130_fd_sc_hd__xnor2_1
X_13261_ _13264_/CLK _13261_/D vssd1 vssd1 vccd1 vccd1 hold161/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_36_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12212_ _12213_/A _12213_/B _12213_/C vssd1 vssd1 vccd1 vccd1 _12214_/A sky130_fd_sc_hd__o21ai_2
X_10473_ _10473_/A _10473_/B vssd1 vssd1 vccd1 vccd1 _10475_/B sky130_fd_sc_hd__nor2_2
X_13192_ _13289_/CLK _13192_/D vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09230__A2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07241__B2 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07241__A1 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ _12143_/A _12143_/B vssd1 vssd1 vccd1 vccd1 _12144_/B sky130_fd_sc_hd__or2_1
XANTENNA__07792__A2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ _12014_/A _12014_/B _12012_/A vssd1 vssd1 vccd1 vccd1 _12085_/A sky130_fd_sc_hd__o21ai_1
X_11025_ _11025_/A _11025_/B vssd1 vssd1 vccd1 vccd1 _11028_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_87_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12976_ _08777_/A _12744_/B hold141/X vssd1 vssd1 vccd1 vccd1 _13258_/D sky130_fd_sc_hd__a21boi_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11927_ _11900_/Y _11902_/X _11907_/X _11926_/X _12382_/S vssd1 vssd1 vccd1 vccd1
+ _11927_/X sky130_fd_sc_hd__o41a_1
XANTENNA__10300__A1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10300__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11858_ _11858_/A _11858_/B vssd1 vssd1 vccd1 vccd1 _11859_/B sky130_fd_sc_hd__and2_1
XANTENNA_19 reg1_val[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11789_ _12200_/A _11789_/B vssd1 vssd1 vccd1 vccd1 _11791_/C sky130_fd_sc_hd__xnor2_1
X_10809_ _10686_/B _10686_/C _10686_/A vssd1 vssd1 vccd1 vccd1 _10812_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10064__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06999__B _07005_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07951_ _08853_/A _07951_/B vssd1 vssd1 vccd1 vccd1 _07955_/A sky130_fd_sc_hd__xor2_1
X_06902_ instruction[14] _06904_/B vssd1 vssd1 vccd1 vccd1 dest_idx[3] sky130_fd_sc_hd__and2_4
XFILLER_0_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07882_ _07883_/B _07883_/A vssd1 vssd1 vccd1 vccd1 _08014_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08732__A1 _08348_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08732__B2 _07181_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06833_ _06632_/X _06833_/B vssd1 vssd1 vccd1 vccd1 _06833_/Y sky130_fd_sc_hd__nand2b_1
X_09621_ _09621_/A _09621_/B vssd1 vssd1 vccd1 vccd1 _09622_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__07535__A2 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06764_ _06762_/Y _06764_/B vssd1 vssd1 vccd1 vccd1 _06868_/C sky130_fd_sc_hd__nand2b_2
X_09552_ _12361_/B _09533_/X _09539_/X _09851_/B vssd1 vssd1 vccd1 vccd1 _09552_/X
+ sky130_fd_sc_hd__o211a_1
X_08503_ _08505_/A _08505_/B vssd1 vssd1 vccd1 vccd1 _08503_/Y sky130_fd_sc_hd__nand2_1
X_06695_ _06783_/A _12658_/A _06641_/A _06694_/X vssd1 vssd1 vccd1 vccd1 _07178_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout255_A _12487_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08496__B1 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09483_ _09484_/A _09484_/B vssd1 vssd1 vccd1 vccd1 _09483_/X sky130_fd_sc_hd__and2_1
XANTENNA__08735__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08434_ _08435_/A _08435_/B vssd1 vssd1 vccd1 vccd1 _08457_/A sky130_fd_sc_hd__or2_1
XFILLER_0_77_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08365_ _08365_/A _08365_/B vssd1 vssd1 vccd1 vccd1 _08373_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07316_ reg1_val[20] _07316_/B vssd1 vssd1 vccd1 vccd1 _07317_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_46_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08296_ _08296_/A _08296_/B vssd1 vssd1 vccd1 vccd1 _08339_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07247_ _08595_/A _07247_/B vssd1 vssd1 vccd1 vccd1 _07249_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07178_ _07178_/A _07178_/B vssd1 vssd1 vccd1 vccd1 _11147_/A sky130_fd_sc_hd__xor2_4
XANTENNA__11555__B1 _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06702__B _07192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08723__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08723__B2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06589__A_N _12250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09819_ _09716_/X _10002_/B _09110_/X vssd1 vssd1 vccd1 vccd1 _09819_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12830_ _12830_/A _12830_/B vssd1 vssd1 vccd1 vccd1 _13025_/A sky130_fd_sc_hd__nor2_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ hold11/X _12786_/B _12760_/Y _13166_/A vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__o211a_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12692_ reg1_val[27] _12708_/B vssd1 vssd1 vccd1 vccd1 _12698_/C sky130_fd_sc_hd__xnor2_2
X_11712_ _11712_/A _11712_/B vssd1 vssd1 vccd1 vccd1 _11713_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10386__S _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11643_ _11588_/Y _11730_/D _11642_/Y vssd1 vssd1 vccd1 vccd1 _11643_/X sky130_fd_sc_hd__a21o_2
XANTENNA__09987__B1 _11838_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10046__B1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11574_ _12187_/A1 _11751_/C _13236_/Q vssd1 vssd1 vccd1 vccd1 _11574_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09451__A2 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13313_ _13318_/CLK hold139/X vssd1 vssd1 vccd1 vccd1 hold137/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10525_ _10482_/A _10482_/B _10480_/X vssd1 vssd1 vccd1 vccd1 _10606_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_122_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13244_ _13248_/CLK hold185/X vssd1 vssd1 vccd1 vccd1 hold213/A sky130_fd_sc_hd__dfxtp_1
X_10456_ _10894_/A _10456_/B vssd1 vssd1 vccd1 vccd1 _10458_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__09476__A _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09739__B1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ hold171/X hold137/X hold176/X vssd1 vssd1 vccd1 vccd1 hold299/A sky130_fd_sc_hd__a21o_1
XANTENNA__07214__A1 _12774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07214__B2 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11010__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12614__B _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11204__A2_N _06928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07708__B _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10387_ _09198_/X _10376_/Y _10386_/X _09837_/A _10384_/X vssd1 vssd1 vccd1 vccd1
+ _10395_/B sky130_fd_sc_hd__a221o_1
X_12126_ reg1_val[26] _10377_/B _07153_/A _06928_/X vssd1 vssd1 vccd1 vccd1 _12126_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_58_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12057_ _12119_/B1 _12183_/C hold286/A vssd1 vssd1 vccd1 vccd1 _12057_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07724__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11008_ _11134_/B2 fanout15/X fanout7/X fanout57/X vssd1 vssd1 vccd1 vccd1 _11009_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11246__A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12959_ hold41/A _06537_/A rst vssd1 vssd1 vccd1 vccd1 _12959_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11077__A2 _09059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08150_ _08150_/A _08150_/B vssd1 vssd1 vccd1 vccd1 _08151_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_90_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12077__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07101_ _10280_/A _07101_/B vssd1 vssd1 vccd1 vccd1 _07162_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_43_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08081_ _08149_/A _08149_/B _08074_/X vssd1 vssd1 vccd1 vccd1 _08103_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07453__A1 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07453__B2 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07032_ _07050_/A _07050_/B _07135_/B vssd1 vssd1 vccd1 vccd1 _07168_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08983_ _08983_/A _08983_/B vssd1 vssd1 vccd1 vccd1 _08984_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07934_ _07933_/A _07933_/B _07933_/C vssd1 vssd1 vccd1 vccd1 _07937_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07865_ _07904_/A _07904_/B vssd1 vssd1 vccd1 vccd1 _07877_/B sky130_fd_sc_hd__or2_2
XANTENNA__07634__A _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09604_ _09605_/A _09605_/B vssd1 vssd1 vccd1 vccd1 _09604_/X sky130_fd_sc_hd__and2b_1
X_07796_ _07797_/A _07797_/B vssd1 vssd1 vccd1 vccd1 _07798_/A sky130_fd_sc_hd__and2_1
XFILLER_0_97_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06816_ _11187_/A _06814_/Y _06815_/X vssd1 vssd1 vccd1 vccd1 _06816_/Y sky130_fd_sc_hd__a21oi_1
X_06747_ reg1_val[6] _06996_/A vssd1 vssd1 vccd1 vccd1 _06750_/A sky130_fd_sc_hd__or2_1
X_09535_ reg1_val[2] curr_PC[2] vssd1 vssd1 vccd1 vccd1 _09535_/Y sky130_fd_sc_hd__nor2_1
X_06678_ instruction[27] _06678_/B vssd1 vssd1 vccd1 vccd1 _12568_/B sky130_fd_sc_hd__and2_4
X_09466_ _09618_/A1 fanout20/X fanout18/X _09618_/B2 vssd1 vssd1 vccd1 vccd1 _09467_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08417_ _08436_/A _08416_/Y _08412_/X vssd1 vssd1 vccd1 vccd1 _08419_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_66_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11603__B fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09397_ _09183_/Y _09370_/X _09396_/X _12373_/A1 _09391_/X vssd1 vssd1 vccd1 vccd1
+ _09397_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_46_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08348_ _08821_/A _08348_/B vssd1 vssd1 vccd1 vccd1 _08385_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_74_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08279_ _08331_/A _08331_/B _08275_/Y vssd1 vssd1 vccd1 vccd1 _08302_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07444__B2 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07444__A1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ _11193_/A _11193_/B _11191_/A vssd1 vssd1 vccd1 vccd1 _11294_/A sky130_fd_sc_hd__o21a_1
XANTENNA__09296__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10310_ _10311_/A _10311_/B vssd1 vssd1 vccd1 vccd1 _10310_/Y sky130_fd_sc_hd__nand2_1
X_10241_ _06798_/Y _10240_/Y _12322_/S vssd1 vssd1 vccd1 vccd1 _10241_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10172_ _10320_/B _10172_/B vssd1 vssd1 vccd1 vccd1 _10174_/B sky130_fd_sc_hd__nand2_1
Xfanout161 _07154_/X vssd1 vssd1 vccd1 vccd1 _08692_/B1 sky130_fd_sc_hd__buf_4
Xfanout172 _10658_/A vssd1 vssd1 vccd1 vccd1 _08855_/A sky130_fd_sc_hd__buf_12
Xfanout183 _08415_/A vssd1 vssd1 vccd1 vccd1 _10155_/A sky130_fd_sc_hd__buf_8
Xfanout150 _11379_/A vssd1 vssd1 vccd1 vccd1 _12131_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__07544__A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08172__A2 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout194 _13151_/A2 vssd1 vssd1 vccd1 vccd1 _13168_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_88_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12813_ hold291/X hold61/X vssd1 vssd1 vccd1 vccd1 _13077_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12256__A1 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12744_ hold63/X _12744_/B vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__or2_1
XFILLER_0_97_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12008__A1 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06607__B _12620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ reg1_val[24] _12714_/A vssd1 vssd1 vccd1 vccd1 _12682_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12008__B2 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11626_ _11626_/A _11626_/B vssd1 vssd1 vccd1 vccd1 _11627_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07435__A1 _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11557_ _11586_/B _11555_/X _11556_/Y vssd1 vssd1 vccd1 vccd1 _11557_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07986__A2 _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10508_ _10504_/Y _10507_/Y _11197_/S vssd1 vssd1 vccd1 vccd1 _10508_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11488_ _06674_/Y _09188_/X _11486_/Y _06676_/B _11487_/X vssd1 vssd1 vccd1 vccd1
+ _11488_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_40_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11519__B1 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13227_ _13243_/CLK _13227_/D vssd1 vssd1 vccd1 vccd1 hold205/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__10145__A _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10439_ _11704_/A fanout47/X _11603_/A _11688_/A vssd1 vssd1 vccd1 vccd1 _10440_/B
+ sky130_fd_sc_hd__o22a_1
X_13158_ _13158_/A _13158_/B vssd1 vssd1 vccd1 vccd1 _13158_/Y sky130_fd_sc_hd__xnor2_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13089_ hold295/A _13088_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13089_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_109_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12109_ _06851_/X _12108_/X _12322_/S vssd1 vssd1 vccd1 vccd1 _12109_/X sky130_fd_sc_hd__mux2_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07454__A _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07650_ _07648_/A _07648_/B _08889_/A vssd1 vssd1 vccd1 vccd1 _08942_/A sky130_fd_sc_hd__o21ai_1
X_06601_ reg2_val[24] _06752_/A _06688_/B1 _06600_/Y vssd1 vssd1 vccd1 vccd1 _07126_/B
+ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_34_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07581_ _07581_/A _07581_/B vssd1 vssd1 vccd1 vccd1 _07619_/A sky130_fd_sc_hd__xor2_4
X_06532_ hold244/X vssd1 vssd1 vccd1 vccd1 _13163_/A sky130_fd_sc_hd__inv_2
XFILLER_0_34_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09320_ _09320_/A _09320_/B vssd1 vssd1 vccd1 vccd1 _09321_/B sky130_fd_sc_hd__xor2_4
XANTENNA__11704__A _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09251_ _10453_/A _09251_/B vssd1 vssd1 vccd1 vccd1 _09256_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08202_ _08202_/A _08202_/B vssd1 vssd1 vccd1 vccd1 _08260_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_63_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09182_ _12361_/B _09178_/X _09181_/X _09851_/B vssd1 vssd1 vccd1 vccd1 _09217_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08133_ _08133_/A _08133_/B vssd1 vssd1 vccd1 vccd1 _08199_/A sky130_fd_sc_hd__xor2_1
XANTENNA_fanout120_A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08064_ _08641_/A _08641_/B vssd1 vssd1 vccd1 vccd1 _08064_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12970__A2 _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout218_A _09392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ _07324_/A _07015_/B vssd1 vssd1 vccd1 vccd1 _07175_/C sky130_fd_sc_hd__or2_1
XANTENNA__07729__A2 _10551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08966_ _08966_/A _08966_/B vssd1 vssd1 vccd1 vccd1 _08974_/A sky130_fd_sc_hd__xor2_4
XANTENNA__07364__A _07364_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07917_ _08443_/A _07917_/B vssd1 vssd1 vccd1 vccd1 _08034_/A sky130_fd_sc_hd__xor2_2
X_08897_ _08897_/A _08897_/B vssd1 vssd1 vccd1 vccd1 _08899_/C sky130_fd_sc_hd__nand2_1
X_07848_ _07848_/A _07848_/B _07848_/C vssd1 vssd1 vccd1 vccd1 _07933_/A sky130_fd_sc_hd__or3_1
XANTENNA__07901__A2 _08672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12789__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ _07775_/A _07775_/B _07789_/A vssd1 vssd1 vccd1 vccd1 _07780_/B sky130_fd_sc_hd__o21ba_2
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09518_ _11089_/A _09517_/A _09212_/Y vssd1 vssd1 vccd1 vccd1 _09518_/Y sky130_fd_sc_hd__a21oi_1
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11997__B1 _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10790_ _12150_/B _10557_/B fanout13/X _12776_/A vssd1 vssd1 vccd1 vccd1 _10791_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _09450_/A _09450_/B vssd1 vssd1 vccd1 vccd1 _09596_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_124_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12460_ _12620_/B _12461_/B vssd1 vssd1 vccd1 vccd1 _12471_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12391_ _12568_/B _12391_/B vssd1 vssd1 vccd1 vccd1 _12392_/B sky130_fd_sc_hd__or2_1
XFILLER_0_74_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11411_ _12200_/A _11411_/B vssd1 vssd1 vccd1 vccd1 _11414_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13040__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11342_ _11342_/A _11342_/B vssd1 vssd1 vccd1 vccd1 _11351_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_22_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06688__A2_N _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_590 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07258__B _07259_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11273_ _11274_/A _11274_/B _11274_/C vssd1 vssd1 vccd1 vccd1 _11275_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13012_ _10169_/A _13020_/B2 hold93/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__o21a_1
XANTENNA__09754__A _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _10224_/A _10224_/B vssd1 vssd1 vccd1 vccd1 _10227_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08393__A2 _10551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11921__B1 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09473__B _09474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ _10155_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10158_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06943__A3 _07087_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10086_ _10086_/A _10086_/B vssd1 vssd1 vccd1 vccd1 _10088_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09893__A2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11524__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10988_ hold295/A _09842_/B _11198_/C _12339_/B1 vssd1 vssd1 vccd1 vccd1 _10988_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12727_ hold36/X _12744_/B _12726_/Y _13013_/C1 vssd1 vssd1 vccd1 vccd1 hold37/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07656__B2 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07656__A1 _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12658_ _12658_/A _12658_/B vssd1 vssd1 vccd1 vccd1 _12660_/C sky130_fd_sc_hd__nand2_2
XANTENNA__08833__A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11609_ _11688_/A _12200_/A vssd1 vssd1 vccd1 vccd1 _11610_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07959__A2 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12589_ _12589_/A _12589_/B vssd1 vssd1 vccd1 vccd1 _12590_/B sky130_fd_sc_hd__or2_2
XANTENNA__10412__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _10015_/A _08820_/B vssd1 vssd1 vccd1 vccd1 _08824_/A sky130_fd_sc_hd__xnor2_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09581__A1 _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07184__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09383__B _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09581__B2 _09295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08751_ _08864_/A _08750_/B _08750_/C vssd1 vssd1 vccd1 vccd1 _08752_/C sky130_fd_sc_hd__a21o_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08682_ _06989_/A _11782_/A _08748_/B1 vssd1 vssd1 vccd1 vccd1 _08683_/C sky130_fd_sc_hd__a21o_1
X_07702_ _07700_/A _07700_/B _07701_/Y vssd1 vssd1 vccd1 vccd1 _08992_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__07912__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07895__A1 _10149_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07633_ _07260_/Y fanout81/X _09295_/B fanout51/X vssd1 vssd1 vccd1 vccd1 _07634_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07895__B2 _10035_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout168_A _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07564_ fanout83/X fanout46/X fanout12/X fanout81/X vssd1 vssd1 vccd1 vccd1 _07565_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09303_ _09301_/X _09303_/B vssd1 vssd1 vccd1 vccd1 _09306_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07495_ _07495_/A _07495_/B vssd1 vssd1 vccd1 vccd1 _07496_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_90_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09234_ _10301_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _09236_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09165_ reg1_val[18] reg1_val[13] _09173_/S vssd1 vssd1 vccd1 vccd1 _09165_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08116_ _08070_/A _08070_/B _08115_/X vssd1 vssd1 vccd1 vccd1 _08633_/B sky130_fd_sc_hd__o21bai_4
XFILLER_0_9_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08072__B2 _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08072__A1 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09096_ _09103_/A _09103_/B _09085_/X _09095_/X vssd1 vssd1 vccd1 vccd1 _09097_/B
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_9_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08047_ _08748_/B1 fanout51/X _12730_/A _08134_/B vssd1 vssd1 vccd1 vccd1 _08048_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09998_ curr_PC[4] curr_PC[5] _09998_/C vssd1 vssd1 vccd1 vccd1 _10138_/B sky130_fd_sc_hd__and3_1
XANTENNA__11609__A _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08949_ _08949_/A _08949_/B vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__nand2_1
X_11960_ _11961_/A _11961_/B vssd1 vssd1 vccd1 vccd1 _12036_/B sky130_fd_sc_hd__or2_1
X_10911_ fanout33/X _11794_/A _12772_/A _10553_/A vssd1 vssd1 vccd1 vccd1 _10912_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_86_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11682__A2 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11891_ _11898_/A vssd1 vssd1 vccd1 vccd1 _11967_/B sky130_fd_sc_hd__inv_2
XANTENNA__11344__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10890__B1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10842_ _10842_/A _10842_/B vssd1 vssd1 vccd1 vccd1 _10843_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_109_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08835__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07638__B2 _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07638__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10773_ _12005_/A _10769_/X _10770_/X _10772_/Y vssd1 vssd1 vccd1 vccd1 dest_val[11]
+ sky130_fd_sc_hd__a22o_4
X_12512_ _12557_/A _12513_/B vssd1 vssd1 vccd1 vccd1 _12514_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12443_ _12443_/A _12443_/B _12443_/C vssd1 vssd1 vccd1 vccd1 _12444_/B sky130_fd_sc_hd__nand3_1
X_12374_ _09200_/X _12368_/Y _12373_/X _12366_/Y vssd1 vssd1 vccd1 vccd1 _12374_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__07269__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07810__A1 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07810__B2 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325_ _11325_/A _11325_/B vssd1 vssd1 vccd1 vccd1 _11327_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11256_ _11256_/A _11256_/B vssd1 vssd1 vccd1 vccd1 _11257_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11187_ _11187_/A _11187_/B vssd1 vssd1 vccd1 vccd1 _11187_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10423__A _12255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ _10207_/A _10207_/B vssd1 vssd1 vccd1 vccd1 _10208_/B sky130_fd_sc_hd__nor2_1
X_10138_ curr_PC[6] _10138_/B vssd1 vssd1 vccd1 vccd1 _10397_/C sky130_fd_sc_hd__and2_2
X_10069_ _10069_/A _10069_/B vssd1 vssd1 vccd1 vccd1 _10071_/B sky130_fd_sc_hd__xor2_4
XANTENNA__07732__A _10578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__B1 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11122__B2 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11122__A1 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09866__A2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10881__B1 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09618__A2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07280_ _08825_/A2 fanout26/X _09476_/A _07389_/B vssd1 vssd1 vccd1 vccd1 _07281_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08563__A _09620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12925__A2 _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07179__A _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold203 hold239/X vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold214 hold214/A vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 hold225/A vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold258 hold258/A vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold269 hold269/A vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ _09921_/A _09921_/B vssd1 vssd1 vccd1 vccd1 _09938_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_1_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09852_ _06762_/Y _09191_/X _09850_/Y _09851_/Y _09845_/X vssd1 vssd1 vccd1 vccd1
+ _09852_/X sky130_fd_sc_hd__o221a_1
XANTENNA__11429__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10164__A2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _08804_/B vssd1 vssd1 vccd1 vccd1 _08803_/Y sky130_fd_sc_hd__inv_2
X_09783_ _08681_/A _07553_/A _10927_/A _09295_/A vssd1 vssd1 vccd1 vccd1 _09784_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11148__B _11148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout285_A _06633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _07031_/Y _07179_/Y fanout94/X _08854_/B2 vssd1 vssd1 vccd1 vccd1 _08735_/B
+ sky130_fd_sc_hd__o22a_1
X_06995_ _06996_/A _06996_/B vssd1 vssd1 vccd1 vccd1 _10035_/A sky130_fd_sc_hd__xnor2_4
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11113__A1 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11113__B2 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08665_ _08837_/B2 _09752_/B fanout14/X _12736_/A vssd1 vssd1 vccd1 vccd1 _08666_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08596_ _08596_/A _08596_/B vssd1 vssd1 vccd1 vccd1 _08597_/B sky130_fd_sc_hd__xor2_1
X_07616_ _07617_/A _07617_/B vssd1 vssd1 vccd1 vccd1 _09226_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__09609__A2 _07132_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07080__C _07080_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07547_ _07548_/A _07548_/B vssd1 vssd1 vccd1 vccd1 _07549_/A sky130_fd_sc_hd__and2_1
XFILLER_0_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07478_ _07270_/A _07270_/B _07267_/A vssd1 vssd1 vccd1 vccd1 _07582_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09217_ _09217_/A _09217_/B vssd1 vssd1 vccd1 vccd1 _09218_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_51_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09148_ reg1_val[25] reg1_val[6] _09172_/S vssd1 vssd1 vccd1 vccd1 _09148_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09079_ _09079_/A _09079_/B vssd1 vssd1 vccd1 vccd1 _12131_/B sky130_fd_sc_hd__nor2_1
XANTENNA__06815__A_N _07178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11110_ _11000_/X _11215_/C _12278_/A vssd1 vssd1 vccd1 vccd1 _11110_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_31_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07817__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12090_ _12090_/A _12090_/B vssd1 vssd1 vccd1 vccd1 _12091_/B sky130_fd_sc_hd__or2_1
XANTENNA__11339__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11041_ _11041_/A _11041_/B vssd1 vssd1 vccd1 vccd1 _11042_/B sky130_fd_sc_hd__and2_1
XANTENNA__07556__B1 _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08648__A _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12992_ _08836_/A _13020_/B2 hold114/X vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__o21a_1
XANTENNA__11104__A1 _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11943_ _12200_/A _11943_/B vssd1 vssd1 vccd1 vccd1 _11947_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11874_ _11875_/A _11875_/B vssd1 vssd1 vccd1 vccd1 _11952_/B sky130_fd_sc_hd__and2_1
XANTENNA__12065__C1 _12064_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10825_ _10825_/A _10825_/B vssd1 vssd1 vccd1 vccd1 _10826_/B sky130_fd_sc_hd__and2_1
XFILLER_0_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10615__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10756_ _12187_/A1 _10874_/B hold219/A vssd1 vssd1 vccd1 vccd1 _10756_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09479__A _09775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ _10686_/A _10686_/B _10686_/C vssd1 vssd1 vccd1 vccd1 _10688_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__08036__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08036__B2 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12426_ _12593_/B _12426_/B vssd1 vssd1 vccd1 vccd1 _12427_/B sky130_fd_sc_hd__or2_1
XANTENNA__09233__B1 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10918__A1 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10918__B2 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10394__A2 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_max_cap250_A _09620_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12357_ _12357_/A _12357_/B vssd1 vssd1 vccd1 vccd1 _12357_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11308_ _11285_/X _11286_/Y _11289_/X _12228_/B1 _11307_/X vssd1 vssd1 vccd1 vccd1
+ _11308_/X sky130_fd_sc_hd__a221o_2
X_12288_ hold165/A _12288_/B vssd1 vssd1 vccd1 vccd1 _12330_/B sky130_fd_sc_hd__or2_1
XFILLER_0_10_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11239_ _12203_/A fanout47/X _11603_/A _12150_/A vssd1 vssd1 vccd1 vccd1 _11240_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10153__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11343__B2 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11343__A1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10146__A2 _10147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06780_ _06783_/A _06649_/A _12568_/B _06778_/X vssd1 vssd1 vccd1 vccd1 _06780_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08558__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08450_ _08588_/A _08776_/B1 _08825_/A2 _08477_/B vssd1 vssd1 vccd1 vccd1 _08451_/B
+ sky130_fd_sc_hd__o22a_1
X_08381_ _07969_/A _08772_/B2 _08772_/A2 _12734_/A vssd1 vssd1 vccd1 vccd1 _08382_/B
+ sky130_fd_sc_hd__o22a_1
X_07401_ _07401_/A _07678_/A vssd1 vssd1 vccd1 vccd1 _07629_/B sky130_fd_sc_hd__nand2_1
X_07332_ _10015_/A _07332_/B vssd1 vssd1 vccd1 vccd1 _07335_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07263_ _07553_/A fanout52/X _10677_/B _10927_/A vssd1 vssd1 vccd1 vccd1 _07264_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11431__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07194_ _08733_/A _10819_/A _07194_/C vssd1 vssd1 vccd1 vccd1 _07195_/B sky130_fd_sc_hd__or3_2
XANTENNA__09224__B1 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09002_ _09968_/A _12357_/A vssd1 vssd1 vccd1 vccd1 _09002_/X sky130_fd_sc_hd__and2_1
XFILLER_0_26_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13020__B2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08578__A2 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11031__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11582__A1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout200_A _09188_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire4 wire4/A vssd1 vssd1 vccd1 vccd1 wire4/X sky130_fd_sc_hd__buf_1
X_09904_ _10527_/A _10677_/A vssd1 vssd1 vccd1 vccd1 _09906_/C sky130_fd_sc_hd__or2_1
XANTENNA__10063__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09835_ _09832_/X _09834_/X _10251_/S vssd1 vssd1 vccd1 vccd1 _09835_/X sky130_fd_sc_hd__mux2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06978_ reg1_val[21] _06978_/B vssd1 vssd1 vccd1 vccd1 _07974_/A sky130_fd_sc_hd__xnor2_4
X_09766_ _09767_/B _09766_/B vssd1 vssd1 vccd1 vccd1 _09879_/A sky130_fd_sc_hd__and2b_1
X_08717_ _08717_/A _08717_/B vssd1 vssd1 vccd1 vccd1 _08720_/B sky130_fd_sc_hd__xnor2_1
X_09697_ _06770_/X _09695_/X _09696_/Y vssd1 vssd1 vccd1 vccd1 _09707_/B sky130_fd_sc_hd__a21oi_1
X_08648_ _08777_/A _08648_/B vssd1 vssd1 vccd1 vccd1 _08650_/B sky130_fd_sc_hd__xnor2_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07091__B _12370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08579_ _08595_/A _08579_/B vssd1 vssd1 vccd1 vccd1 _08596_/A sky130_fd_sc_hd__xnor2_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09299__A _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09463__B1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11590_ fanout27/X _11935_/A _12772_/A _12205_/A vssd1 vssd1 vccd1 vccd1 _11591_/B
+ sky130_fd_sc_hd__o22a_1
X_10610_ _10358_/X _10483_/X _10484_/X vssd1 vssd1 vccd1 vccd1 _10610_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ fanout36/X fanout57/X _11222_/A _06959_/Y vssd1 vssd1 vccd1 vccd1 _10542_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13260_ _13264_/CLK hold97/X vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08931__A _08932_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ _12264_/B _12211_/B vssd1 vssd1 vccd1 vccd1 _12213_/C sky130_fd_sc_hd__nor2_1
X_10472_ _10312_/A _10312_/B _10310_/Y vssd1 vssd1 vccd1 vccd1 _10475_/A sky130_fd_sc_hd__o21a_2
X_13191_ _13310_/CLK _13191_/D vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12453__A _12614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07241__A2 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ _12143_/A _12143_/B vssd1 vssd1 vccd1 vccd1 _12144_/A sky130_fd_sc_hd__nand2_1
X_12073_ _11973_/B _12221_/A _11973_/A vssd1 vssd1 vccd1 vccd1 _12107_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07529__B1 _12713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11024_ _11024_/A _11024_/B vssd1 vssd1 vccd1 vccd1 _11025_/B sky130_fd_sc_hd__nor2_1
X_12975_ hold134/X _12723_/A _13170_/B hold140/X _13066_/A vssd1 vssd1 vccd1 vccd1
+ hold141/A sky130_fd_sc_hd__o221a_1
Xclkbuf_4_2_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13248_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_87_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11926_ _11926_/A _11926_/B _11926_/C _11920_/X vssd1 vssd1 vccd1 vccd1 _11926_/X
+ sky130_fd_sc_hd__or4b_1
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10300__A2 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11857_ _11858_/A _11858_/B vssd1 vssd1 vccd1 vccd1 _11938_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_28_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06626__A _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11788_ _11935_/A fanout15/X fanout6/X _12772_/A vssd1 vssd1 vccd1 vccd1 _11789_/B
+ sky130_fd_sc_hd__o22a_1
X_10808_ _10453_/A _10658_/B _10659_/Y vssd1 vssd1 vccd1 vccd1 _10813_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_125_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10739_ _10617_/A _10740_/B _10740_/C vssd1 vssd1 vccd1 vccd1 _10739_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__08544__C _08544_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09002__A _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10064__B2 _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10064__A1 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13002__A1 _06987_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07768__B1 _08692_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ _12415_/B _12409_/B vssd1 vssd1 vccd1 vccd1 new_PC[4] sky130_fd_sc_hd__and2_4
XFILLER_0_51_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07950_ _07173_/Y _10694_/A _10551_/A _07182_/X vssd1 vssd1 vccd1 vccd1 _07951_/B
+ sky130_fd_sc_hd__a22o_1
X_06901_ instruction[13] _06904_/B vssd1 vssd1 vccd1 vccd1 dest_idx[2] sky130_fd_sc_hd__and2_4
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07881_ _07888_/A _07888_/B _07860_/Y vssd1 vssd1 vccd1 vccd1 _07883_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08732__A2 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06832_ reg1_val[23] _07119_/A _06872_/B _06825_/Y _06831_/Y vssd1 vssd1 vccd1 vccd1
+ _06833_/B sky130_fd_sc_hd__a221o_1
X_09620_ _09620_/A _09621_/B vssd1 vssd1 vccd1 vccd1 _09620_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07192__A _07192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06763_ reg1_val[4] _07001_/C vssd1 vssd1 vccd1 vccd1 _06764_/B sky130_fd_sc_hd__nand2_1
X_09551_ _12284_/B _09533_/X _12322_/S vssd1 vssd1 vccd1 vccd1 _09551_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08502_ _08502_/A _08502_/B vssd1 vssd1 vccd1 vccd1 _08505_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_93_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06694_ reg2_val[15] _06729_/B vssd1 vssd1 vccd1 vccd1 _06694_/X sky130_fd_sc_hd__and2_1
XANTENNA__12292__A2 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08496__B2 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08496__A1 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09482_ _09482_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09484_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08433_ _08433_/A _08433_/B vssd1 vssd1 vccd1 vccd1 _08435_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout150_A _11379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08364_ _08406_/A _08406_/B _08361_/Y vssd1 vssd1 vccd1 vccd1 _08373_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_58_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout248_A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09445__B1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09996__A1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ _10559_/A _07315_/B vssd1 vssd1 vccd1 vccd1 _07329_/A sky130_fd_sc_hd__xnor2_1
X_08295_ _08295_/A _08295_/B _08295_/C vssd1 vssd1 vccd1 vccd1 _08295_/X sky130_fd_sc_hd__and3_1
XFILLER_0_104_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07246_ _08758_/A2 fanout20/X fanout18/X _06864_/A vssd1 vssd1 vccd1 vccd1 _07247_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_42_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07177_ _07192_/A _07197_/A _07303_/A _07303_/C _07303_/B vssd1 vssd1 vccd1 vccd1
+ _07178_/B sky130_fd_sc_hd__o41a_2
XFILLER_0_112_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07759__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07367__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__A1 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09582__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08723__A2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09818_ _10229_/B _09818_/B vssd1 vssd1 vccd1 vccd1 _10002_/B sky130_fd_sc_hd__xnor2_4
XANTENNA_fanout63_A _07119_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ _09881_/B _09749_/B vssd1 vssd1 vccd1 vccd1 _09771_/A sky130_fd_sc_hd__nor2_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10818__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _12760_/A _12786_/B vssd1 vssd1 vccd1 vccd1 _12760_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_96_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12687_/B _12690_/B _12685_/X vssd1 vssd1 vccd1 vccd1 _12693_/A sky130_fd_sc_hd__a21o_1
X_11711_ _11712_/B _11712_/A vssd1 vssd1 vccd1 vccd1 _11711_/X sky130_fd_sc_hd__and2b_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11642_ _11588_/Y _11730_/D _12223_/B1 vssd1 vssd1 vccd1 vccd1 _11642_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10046__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10046__A1 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13312_ _13312_/CLK _13312_/D vssd1 vssd1 vccd1 vccd1 hold103/A sky130_fd_sc_hd__dfxtp_1
X_11573_ hold168/A _11573_/B vssd1 vssd1 vccd1 vccd1 _11751_/C sky130_fd_sc_hd__or2_1
XFILLER_0_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10524_ _10524_/A _10524_/B vssd1 vssd1 vccd1 vccd1 _11000_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13243_ _13243_/CLK _13243_/D vssd1 vssd1 vccd1 vccd1 hold183/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09739__A1 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ _12782_/A fanout56/X fanout20/X fanout98/X vssd1 vssd1 vccd1 vccd1 _10456_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09476__B _12349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09739__B2 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ hold176/X _12721_/B _12716_/Y _12722_/A vssd1 vssd1 vccd1 vccd1 _13176_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07214__A2 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07277__A _12255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10386_ _10244_/X _10385_/X _10752_/S vssd1 vssd1 vccd1 vccd1 _10386_/X sky130_fd_sc_hd__mux2_1
X_12125_ _06619_/A _09194_/Y _10638_/B vssd1 vssd1 vccd1 vccd1 _12125_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_58_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08175__B1 _08672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ hold262/A _12056_/B vssd1 vssd1 vccd1 vccd1 _12183_/C sky130_fd_sc_hd__or2_1
XFILLER_0_74_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _11007_/A _11007_/B vssd1 vssd1 vccd1 vccd1 _11048_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10150__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12958_ rst _12958_/B vssd1 vssd1 vccd1 vccd1 _13249_/D sky130_fd_sc_hd__nor2_1
XANTENNA__08836__A _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12889_ _13162_/A _13162_/B vssd1 vssd1 vccd1 vccd1 _12891_/C sky130_fd_sc_hd__or2_1
XANTENNA__07740__A _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11909_ reg1_val[23] curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11910_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_114_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07989__B1 _07869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07100_ _08825_/A2 _07389_/B fanout26/X _08588_/A vssd1 vssd1 vccd1 vccd1 _07101_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08080_ _08080_/A _08080_/B vssd1 vssd1 vccd1 vccd1 _08149_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_113_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08571__A _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07453__A2 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07031_ _07031_/A _07031_/B vssd1 vssd1 vccd1 vccd1 _07031_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_3_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08982_ _08982_/A _08982_/B vssd1 vssd1 vccd1 vccd1 _08984_/A sky130_fd_sc_hd__xor2_1
X_07933_ _07933_/A _07933_/B _07933_/C vssd1 vssd1 vccd1 vccd1 _07937_/A sky130_fd_sc_hd__and3_1
X_07864_ _08777_/A _07864_/B vssd1 vssd1 vccd1 vccd1 _07904_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07913__B1 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06815_ _07178_/A reg1_val[15] vssd1 vssd1 vccd1 vccd1 _06815_/X sky130_fd_sc_hd__and2b_1
X_09603_ _10551_/B _09603_/B vssd1 vssd1 vccd1 vccd1 _09605_/B sky130_fd_sc_hd__xnor2_2
X_07795_ _11604_/A _07795_/B vssd1 vssd1 vccd1 vccd1 _07797_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06746_ _06783_/A _06649_/A _12593_/B _06745_/X vssd1 vssd1 vccd1 vccd1 _06996_/A
+ sky130_fd_sc_hd__a31o_4
X_09534_ _09374_/A _09373_/A _09373_/B vssd1 vssd1 vccd1 vccd1 _09538_/A sky130_fd_sc_hd__o21ba_1
X_06677_ _06865_/B vssd1 vssd1 vccd1 vccd1 _06677_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09465_ _09465_/A _09465_/B vssd1 vssd1 vccd1 vccd1 _09474_/A sky130_fd_sc_hd__xnor2_1
X_08416_ _08436_/B vssd1 vssd1 vccd1 vccd1 _08416_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09969__A1 _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ _11195_/A _09395_/Y _09214_/A vssd1 vssd1 vccd1 vccd1 _09396_/X sky130_fd_sc_hd__o21a_1
XANTENNA__11225__B1 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08347_ _08855_/A _08347_/B vssd1 vssd1 vccd1 vccd1 _08385_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08278_ _08278_/A _08278_/B vssd1 vssd1 vccd1 vccd1 _08331_/B sky130_fd_sc_hd__xor2_1
XANTENNA__07444__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_750 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07229_ _09610_/A _07229_/B vssd1 vssd1 vccd1 vccd1 _07233_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06713__B _07303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10240_ _06750_/A _10106_/Y _06748_/X vssd1 vssd1 vccd1 vccd1 _10240_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07097__A _10169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10171_ _10170_/B _10171_/B vssd1 vssd1 vccd1 vccd1 _10172_/B sky130_fd_sc_hd__nand2b_1
Xfanout140 _09888_/B2 vssd1 vssd1 vccd1 vccd1 _08837_/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout173 _08232_/A vssd1 vssd1 vccd1 vccd1 _10658_/A sky130_fd_sc_hd__buf_12
Xfanout162 _08692_/A2 vssd1 vssd1 vccd1 vccd1 _08588_/B sky130_fd_sc_hd__clkbuf_8
Xfanout151 _12230_/A vssd1 vssd1 vccd1 vccd1 _12278_/A sky130_fd_sc_hd__buf_4
XANTENNA__11347__A _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout195 _13151_/A2 vssd1 vssd1 vccd1 vccd1 _13165_/A2 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06707__A1 _06898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout184 _08415_/A vssd1 vssd1 vccd1 vccd1 _09610_/A sky130_fd_sc_hd__buf_4
X_12812_ hold274/X hold9/X vssd1 vssd1 vccd1 vccd1 _13082_/A sky130_fd_sc_hd__nand2b_1
X_12743_ _10281_/A _12980_/A2 hold74/X _13066_/A vssd1 vssd1 vccd1 vccd1 _13193_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__10267__A1 _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12674_ _12674_/A _12678_/D vssd1 vssd1 vccd1 vccd1 loadstore_address[23] sky130_fd_sc_hd__xnor2_4
XANTENNA__09409__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12008__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11216__B1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11625_ _11626_/A _11626_/B vssd1 vssd1 vccd1 vccd1 _11722_/A sky130_fd_sc_hd__and2_1
XFILLER_0_107_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11556_ _11586_/B _11555_/X _09110_/X vssd1 vssd1 vccd1 vccd1 _11556_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10507_ _10507_/A vssd1 vssd1 vccd1 vccd1 _10507_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_69_16 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12625__B _12626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10990__A2 _09188_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11487_ _07075_/A _11923_/A2 _10377_/B reg1_val[18] vssd1 vssd1 vccd1 vccd1 _11487_/X
+ sky130_fd_sc_hd__o22a_1
X_13226_ _13243_/CLK _13226_/D vssd1 vssd1 vccd1 vccd1 hold198/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11519__A1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11519__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10438_ _12019_/A _10438_/B vssd1 vssd1 vccd1 vccd1 _10442_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13157_ _13157_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _13158_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10369_ _11973_/A _10370_/B _10370_/C vssd1 vssd1 vccd1 vccd1 _10369_/Y sky130_fd_sc_hd__o21ai_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12641__A _12641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13088_ _13088_/A _13088_/B vssd1 vssd1 vccd1 vccd1 _13088_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_85_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12108_ _12045_/A _12043_/X _06596_/Y vssd1 vssd1 vccd1 vccd1 _12108_/X sky130_fd_sc_hd__o21a_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12039_ _11898_/A _11898_/B _12102_/A _12038_/X vssd1 vssd1 vccd1 vccd1 _12040_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06600_ _06687_/A _12603_/B vssd1 vssd1 vccd1 vccd1 _06600_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07580_ _07578_/Y _07580_/B vssd1 vssd1 vccd1 vccd1 _07581_/B sky130_fd_sc_hd__and2b_1
X_06531_ hold242/X vssd1 vssd1 vccd1 vccd1 _13167_/A sky130_fd_sc_hd__inv_2
XANTENNA__11704__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09250_ _10527_/A _11794_/A fanout62/X _10452_/B2 vssd1 vssd1 vccd1 vccd1 _09251_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08201_ _08201_/A _08201_/B vssd1 vssd1 vccd1 vccd1 _08202_/B sky130_fd_sc_hd__and2_1
XANTENNA__06882__B1 _12345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09181_ _09374_/A _09180_/X _11197_/S vssd1 vssd1 vccd1 vccd1 _09181_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_16_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08132_ _08198_/A _08198_/B _08128_/X vssd1 vssd1 vccd1 vccd1 _08146_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__12955__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08063_ _08066_/A _08066_/B _08022_/X vssd1 vssd1 vccd1 vccd1 _08641_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_114_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07014_ _10658_/A vssd1 vssd1 vccd1 vccd1 _10453_/A sky130_fd_sc_hd__inv_4
XANTENNA__10336__A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07645__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08965_ _08955_/A _08955_/B _08956_/Y vssd1 vssd1 vccd1 vccd1 _08975_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__08139__B1 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07916_ _07149_/Y _07168_/Y _07179_/A _07155_/X vssd1 vssd1 vccd1 vccd1 _07917_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08896_ _08896_/A _08896_/B vssd1 vssd1 vccd1 vccd1 _08897_/B sky130_fd_sc_hd__nand2_1
X_07847_ _07847_/A _07847_/B vssd1 vssd1 vccd1 vccd1 _07848_/C sky130_fd_sc_hd__or2_1
XFILLER_0_98_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07778_ _07788_/B _07778_/B vssd1 vssd1 vccd1 vccd1 _07789_/A sky130_fd_sc_hd__and2b_1
XANTENNA__08476__A _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06729_ reg2_val[9] _06729_/B vssd1 vssd1 vccd1 vccd1 _06729_/X sky130_fd_sc_hd__and2_1
X_09517_ _09517_/A vssd1 vssd1 vccd1 vccd1 _09517_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06708__B _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_734 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11997__A1 _07126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout26_A _07099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09448_ _09610_/A _09448_/B vssd1 vssd1 vccd1 vccd1 _09450_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12726__A _12726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09379_ _09379_/A _09379_/B vssd1 vssd1 vccd1 vccd1 _09379_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_105_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12390_ _12568_/B _12391_/B vssd1 vssd1 vccd1 vccd1 _12401_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11410_ _11688_/A fanout15/X fanout6/X fanout70/X vssd1 vssd1 vccd1 vccd1 _11411_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09406__A3 _09281_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11341_ _11342_/A _11342_/B vssd1 vssd1 vccd1 vccd1 _11341_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_105_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08378__B1 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11272_ _11272_/A _11272_/B vssd1 vssd1 vccd1 vccd1 _11274_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12461__A _12620_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13011_ hold124/A _13013_/A2 _13020_/A2 hold92/X _13028_/A vssd1 vssd1 vccd1 vccd1
+ hold93/A sky130_fd_sc_hd__o221a_1
X_10223_ _10223_/A _10223_/B vssd1 vssd1 vccd1 vccd1 _10224_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_30_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10154_ _10155_/B _10155_/A vssd1 vssd1 vccd1 vccd1 _10154_/X sky130_fd_sc_hd__and2b_1
XANTENNA__07555__A _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06943__A4 _07086_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10085_ _10085_/A _10085_/B vssd1 vssd1 vccd1 vccd1 _10086_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_85_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10987_ _09842_/B _11198_/C hold295/A vssd1 vssd1 vccd1 vccd1 _10987_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06618__B _07153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ _12726_/A _12788_/B vssd1 vssd1 vccd1 vccd1 _12726_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07656__A2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12657_ _12657_/A _12657_/B _12657_/C _12657_/D vssd1 vssd1 vccd1 vccd1 _12660_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_108_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12937__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11608_ _11794_/A fanout15/X fanout6/X _11704_/A vssd1 vssd1 vccd1 vccd1 _11610_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10412__A1 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12588_ reg1_val[6] _12588_/B vssd1 vssd1 vccd1 vccd1 _12589_/B sky130_fd_sc_hd__and2_1
XFILLER_0_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10412__B2 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11539_ _11539_/A _11539_/B vssd1 vssd1 vccd1 vccd1 _11540_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_111_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13209_ _13305_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09581__A2 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08864_/A _08750_/B _08750_/C vssd1 vssd1 vccd1 vccd1 _08864_/B sky130_fd_sc_hd__nand3_2
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08681_ _08681_/A _08681_/B vssd1 vssd1 vccd1 vccd1 _08683_/B sky130_fd_sc_hd__or2_1
X_07701_ _08983_/B _08983_/A vssd1 vssd1 vccd1 vccd1 _07701_/Y sky130_fd_sc_hd__nand2b_1
X_07632_ _07632_/A _07632_/B vssd1 vssd1 vccd1 vccd1 _07651_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07895__A2 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09302_ _09302_/A _09302_/B _09302_/C _09302_/D vssd1 vssd1 vccd1 vccd1 _09303_/B
+ sky130_fd_sc_hd__or4_1
X_07563_ _07561_/X _07563_/B vssd1 vssd1 vccd1 vccd1 _07566_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_118_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07494_ _07590_/A _07494_/B vssd1 vssd1 vccd1 vccd1 _07495_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_61_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09233_ _08821_/B _10064_/B2 _09888_/B2 fanout36/X vssd1 vssd1 vccd1 vccd1 _09234_/B
+ sky130_fd_sc_hd__o22a_1
Xclkbuf_4_15_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13318_/CLK sky130_fd_sc_hd__clkbuf_8
XANTENNA__13141__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09164_ _09162_/X _09163_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09164_/X sky130_fd_sc_hd__mux2_1
X_08115_ _08118_/A _08118_/B vssd1 vssd1 vccd1 vccd1 _08115_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_44_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08072__A2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09095_ _08963_/A _08963_/B _09094_/X vssd1 vssd1 vccd1 vccd1 _09095_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08046_ _08821_/A _09752_/B vssd1 vssd1 vccd1 vccd1 _08109_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_102_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07280__B1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09997_ curr_PC[3] curr_PC[4] _09712_/B curr_PC[5] vssd1 vssd1 vccd1 vccd1 _09997_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11609__B _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ _08923_/A _08923_/B _08921_/X vssd1 vssd1 vccd1 vccd1 _08955_/A sky130_fd_sc_hd__a21o_1
X_08879_ _08880_/A _08880_/B vssd1 vssd1 vccd1 vccd1 _08879_/X sky130_fd_sc_hd__and2_1
X_10910_ _10910_/A _10910_/B vssd1 vssd1 vccd1 vccd1 _10921_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_67_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11419__B1 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ _11890_/A _11890_/B vssd1 vssd1 vccd1 vccd1 _11898_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_67_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10841_ _10842_/A _10842_/B vssd1 vssd1 vccd1 vccd1 _10841_/X sky130_fd_sc_hd__or2_1
XFILLER_0_94_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08835__A1 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__B2 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07638__A2 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10772_ _12556_/S _10772_/B vssd1 vssd1 vccd1 vccd1 _10772_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_109_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12511_ reg1_val[20] curr_PC[20] _12524_/S vssd1 vssd1 vccd1 vccd1 _12513_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_66_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12442_ _12443_/A _12443_/B _12443_/C vssd1 vssd1 vccd1 vccd1 _12450_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12373_ _12373_/A1 _09178_/X _09183_/Y _09215_/Y _12372_/X vssd1 vssd1 vccd1 vccd1
+ _12373_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_50_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07810__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11324_ _11325_/A _11325_/B vssd1 vssd1 vccd1 vccd1 _11434_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11255_ _11256_/A _11256_/B vssd1 vssd1 vccd1 vccd1 _11255_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__07285__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10206_ _10206_/A _10206_/B _10206_/C vssd1 vssd1 vccd1 vccd1 _10207_/B sky130_fd_sc_hd__nor3_1
X_11186_ _06814_/Y _11185_/Y _11738_/S vssd1 vssd1 vccd1 vccd1 _11187_/B sky130_fd_sc_hd__mux2_1
X_10137_ _10102_/Y _10105_/X _10136_/Y _12345_/A vssd1 vssd1 vccd1 vccd1 _10137_/X
+ sky130_fd_sc_hd__a31o_2
X_10068_ _10069_/A _10069_/B vssd1 vssd1 vccd1 vccd1 _10187_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07326__B2 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__A1 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11122__A2 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10330__B1 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12709_ _12707_/X _12709_/B vssd1 vssd1 vccd1 vccd1 _12711_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_73_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 hold215/A vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold259 hold259/A vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold248 hold297/A vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 hold237/A vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__A1 _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09920_ _09919_/B _09919_/C _09919_/A vssd1 vssd1 vccd1 vccd1 _09921_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12689__A2 _07086_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09851_ _12284_/A _09851_/B vssd1 vssd1 vccd1 vccd1 _09851_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09554__A2 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11429__B _11429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06672__A2_N _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08802_ _08801_/A _08801_/B _08801_/C vssd1 vssd1 vccd1 vccd1 _08804_/B sky130_fd_sc_hd__a21o_1
X_06994_ _07595_/A _06994_/B vssd1 vssd1 vccd1 vccd1 _07010_/A sky130_fd_sc_hd__or2_1
X_09782_ _09573_/A _09573_/B _09570_/A vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__o21ai_2
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _08733_/A _08733_/B vssd1 vssd1 vccd1 vccd1 _08741_/A sky130_fd_sc_hd__xnor2_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout180_A _12742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13136__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08514__B1 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout278_A _12658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11113__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08664_ _08664_/A _08664_/B vssd1 vssd1 vccd1 vccd1 _08667_/A sky130_fd_sc_hd__xor2_2
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08595_ _08595_/A _08595_/B _09514_/A vssd1 vssd1 vccd1 vccd1 _09034_/A sky130_fd_sc_hd__or3_1
X_07615_ _07615_/A _07615_/B vssd1 vssd1 vccd1 vccd1 _07617_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_119_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07546_ _10555_/A _07546_/B vssd1 vssd1 vccd1 vccd1 _07548_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09216_ _09178_/X _09183_/Y _09215_/Y _09158_/S _09204_/X vssd1 vssd1 vccd1 vccd1
+ _09217_/B sky130_fd_sc_hd__a221o_1
X_07477_ _07479_/B _07479_/A vssd1 vssd1 vccd1 vccd1 _07482_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__12377__A1 _12370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09147_ reg1_val[24] reg1_val[7] _09173_/S vssd1 vssd1 vccd1 vccd1 _09147_/X sky130_fd_sc_hd__mux2_1
X_09078_ _11820_/B _11820_/C _09076_/Y _11977_/A vssd1 vssd1 vccd1 vccd1 _09079_/B
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08029_ _08071_/A _08071_/B vssd1 vssd1 vccd1 vccd1 _08033_/A sky130_fd_sc_hd__or2_1
XANTENNA__12129__A1 _09198_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout93_A fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11040_ _11041_/A _11041_/B vssd1 vssd1 vccd1 vccd1 _11150_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_99_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10560__B1 _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12991_ _13265_/Q _12723_/A _13170_/B hold113/X _13013_/C1 vssd1 vssd1 vccd1 vccd1
+ hold114/A sky130_fd_sc_hd__o221a_1
XFILLER_0_99_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11942_ _12150_/B fanout15/X fanout6/X _12776_/A vssd1 vssd1 vccd1 vccd1 _11943_/B
+ sky130_fd_sc_hd__o22a_1
X_11873_ _11952_/A _11873_/B vssd1 vssd1 vccd1 vccd1 _11875_/B sky130_fd_sc_hd__nor2_1
X_10824_ _10824_/A _10824_/B _10824_/C vssd1 vssd1 vccd1 vccd1 _10825_/B sky130_fd_sc_hd__or3_1
XFILLER_0_82_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10615__A1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10755_ hold205/A _10755_/B vssd1 vssd1 vccd1 vccd1 _10874_/B sky130_fd_sc_hd__or2_1
XFILLER_0_109_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10686_ _10686_/A _10686_/B _10686_/C vssd1 vssd1 vccd1 vccd1 _10688_/A sky130_fd_sc_hd__and3_1
XANTENNA__08036__A2 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12425_ _12593_/B _12426_/B vssd1 vssd1 vccd1 vccd1 _12436_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09233__A1 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12356_ _12322_/S _06857_/X _12355_/X vssd1 vssd1 vccd1 vccd1 _12357_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__10918__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09233__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11307_ _09851_/B _11295_/X _11301_/X _11306_/Y vssd1 vssd1 vccd1 vccd1 _11307_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12287_ hold244/A _09842_/B _12337_/B _12286_/Y _12339_/B1 vssd1 vssd1 vccd1 vccd1
+ _12295_/A sky130_fd_sc_hd__a311o_2
XFILLER_0_77_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11238_ _11853_/A _11238_/B vssd1 vssd1 vccd1 vccd1 _11328_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11249__B _11250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11343__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ _11169_/A _11169_/B vssd1 vssd1 vccd1 vccd1 _11171_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_117_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08380_ _08383_/A _08383_/B vssd1 vssd1 vccd1 vccd1 _08380_/X sky130_fd_sc_hd__or2_1
X_07400_ _07401_/A _07400_/B _07400_/C vssd1 vssd1 vccd1 vccd1 _07678_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07331_ _08681_/A _10064_/B2 fanout33/X _09888_/B2 vssd1 vssd1 vccd1 vccd1 _07332_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07262_ _07261_/B _07260_/B _11429_/A vssd1 vssd1 vccd1 vccd1 _07262_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_115_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08027__A2 _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07193_ _08733_/A _10819_/A _07194_/C vssd1 vssd1 vccd1 vccd1 _07195_/A sky130_fd_sc_hd__nand3_1
X_09001_ _09660_/A _09001_/B vssd1 vssd1 vccd1 vccd1 _09559_/A sky130_fd_sc_hd__xor2_4
XANTENNA__09224__A1 _09559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07235__B1 _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11031__A1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11031__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10790__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire5 wire5/A vssd1 vssd1 vccd1 vccd1 wire5/X sky130_fd_sc_hd__buf_1
X_09903_ _07139_/A _07139_/B _10452_/B2 vssd1 vssd1 vccd1 vccd1 _09906_/B sky130_fd_sc_hd__a21o_1
X_09834_ _09690_/X _10865_/B _11089_/A vssd1 vssd1 vccd1 vccd1 _09834_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08749__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _07115_/X fanout9/X _09764_/Y _09898_/A vssd1 vssd1 vccd1 vccd1 _09767_/B
+ sky130_fd_sc_hd__o22ai_2
XANTENNA__06761__A2 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06977_ reg1_val[21] _06978_/B vssd1 vssd1 vccd1 vccd1 _09926_/A sky130_fd_sc_hd__xor2_4
X_08716_ _08717_/A _08717_/B vssd1 vssd1 vccd1 vccd1 _08722_/B sky130_fd_sc_hd__nand2b_1
X_09696_ _06770_/X _09695_/X _09192_/Y vssd1 vssd1 vccd1 vccd1 _09696_/Y sky130_fd_sc_hd__o21ai_1
X_08647_ _10156_/B2 _09925_/A1 _07179_/Y _08776_/B1 vssd1 vssd1 vccd1 vccd1 _08648_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07091__C _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12047__B1 _09079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08578_ _06864_/A _09478_/B2 _08758_/A2 _09476_/A vssd1 vssd1 vccd1 vccd1 _08579_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07529_ _09968_/A _07528_/X _12713_/A vssd1 vssd1 vccd1 vccd1 _07529_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09463__B2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09463__A1 _10553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_474 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10540_ _10662_/A _10540_/B vssd1 vssd1 vccd1 vccd1 _10544_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10471_ _10341_/A _10341_/B _10339_/Y vssd1 vssd1 vccd1 vccd1 _10476_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_17_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12734__A _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12210_ _12264_/A _12209_/C _12209_/A vssd1 vssd1 vccd1 vccd1 _12211_/B sky130_fd_sc_hd__o21a_1
X_13190_ _13310_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12141_ _12200_/A _12141_/B vssd1 vssd1 vccd1 vccd1 _12143_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12072_ _12072_/A _12072_/B vssd1 vssd1 vccd1 vccd1 _12221_/A sky130_fd_sc_hd__and2_1
XANTENNA__07529__A1 _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11023_ _11024_/A _11024_/B vssd1 vssd1 vccd1 vccd1 _11025_/A sky130_fd_sc_hd__and2_1
XANTENNA__09078__D_N _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12974_ _07080_/C _12744_/B hold135/X vssd1 vssd1 vccd1 vccd1 hold136/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_99_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11925_ _12373_/A1 _10386_/X _11913_/B _09183_/Y _11924_/Y vssd1 vssd1 vccd1 vccd1
+ _11926_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_59_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_0_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08394__A _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11856_ _12019_/A _11856_/B vssd1 vssd1 vccd1 vccd1 _11858_/B sky130_fd_sc_hd__xor2_1
XANTENNA__06626__B _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ _10807_/A _10807_/B vssd1 vssd1 vccd1 vccd1 _10815_/A sky130_fd_sc_hd__xnor2_1
X_11787_ _11701_/A _11701_/B _11691_/A vssd1 vssd1 vccd1 vccd1 _11800_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10738_ _10650_/X _10774_/B _10737_/Y vssd1 vssd1 vccd1 vccd1 _10738_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10064__A2 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12408_ _12408_/A _12408_/B _12408_/C vssd1 vssd1 vccd1 vccd1 _12409_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13002__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12644__A _12644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10669_ _10670_/A _10670_/B vssd1 vssd1 vccd1 vccd1 _10824_/A sky130_fd_sc_hd__and2_1
XFILLER_0_112_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07768__A1 _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07768__B2 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12339_ hold287/A _09842_/B _12337_/X _12339_/B1 vssd1 vssd1 vccd1 vccd1 _12339_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06900_ instruction[12] _06904_/B vssd1 vssd1 vccd1 vccd1 dest_idx[1] sky130_fd_sc_hd__and2_4
X_07880_ _07880_/A _07880_/B vssd1 vssd1 vccd1 vccd1 _07888_/B sky130_fd_sc_hd__xor2_4
X_06831_ _06829_/X _06830_/Y _11906_/A vssd1 vssd1 vccd1 vccd1 _06831_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06762_ reg1_val[4] _07001_/C vssd1 vssd1 vccd1 vccd1 _06762_/Y sky130_fd_sc_hd__nor2_1
X_09550_ reg1_val[2] _10377_/B _09549_/Y _09201_/X vssd1 vssd1 vccd1 vccd1 _09550_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12277__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08501_ _08524_/A _08524_/B _08490_/Y vssd1 vssd1 vccd1 vccd1 _08505_/A sky130_fd_sc_hd__a21oi_2
X_09481_ _09481_/A _09481_/B vssd1 vssd1 vccd1 vccd1 _09482_/B sky130_fd_sc_hd__xnor2_2
X_06693_ _06693_/A _06693_/B vssd1 vssd1 vccd1 vccd1 _11289_/A sky130_fd_sc_hd__nor2_2
X_08432_ _08432_/A _08432_/B vssd1 vssd1 vccd1 vccd1 _08435_/A sky130_fd_sc_hd__xor2_1
XANTENNA__08496__A2 _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12538__B _12538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08363_ _08390_/A _08363_/B vssd1 vssd1 vccd1 vccd1 _08406_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09445__B2 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09445__A1 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08294_ _08294_/A _08294_/B vssd1 vssd1 vccd1 vccd1 _08295_/C sky130_fd_sc_hd__xnor2_1
X_07314_ _10557_/B fanout83/X fanout13/X fanout81/X vssd1 vssd1 vccd1 vccd1 _07315_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_128_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07245_ _07434_/B _07245_/B vssd1 vssd1 vccd1 vccd1 _12786_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10058__B _10147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07759__A1 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ _07197_/A _07303_/A _07303_/C _07303_/B vssd1 vssd1 vccd1 vccd1 _07192_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_42_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07759__B2 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout300 _06540_/Y vssd1 vssd1 vccd1 vccd1 _07134_/A sky130_fd_sc_hd__buf_6
XANTENNA__07086__C _07086_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09817_ _09511_/B _09816_/X _09815_/X vssd1 vssd1 vccd1 vccd1 _09818_/B sky130_fd_sc_hd__o21a_2
X_09748_ _09748_/A _09748_/B vssd1 vssd1 vccd1 vccd1 _09749_/B sky130_fd_sc_hd__and2_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__A1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout56_A _07181_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09679_ _09356_/X _09366_/X _09679_/S vssd1 vssd1 vccd1 vccd1 _09679_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10818__B2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11710_ _11797_/B _11710_/B vssd1 vssd1 vccd1 vccd1 _11712_/B sky130_fd_sc_hd__or2_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11491__A1 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12690_ _12698_/A _12690_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[26] sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11812_/A _12216_/A vssd1 vssd1 vccd1 vccd1 _11730_/D sky130_fd_sc_hd__xnor2_1
X_11572_ hold280/A _12119_/B1 _11664_/B _11571_/Y _11400_/A vssd1 vssd1 vccd1 vccd1
+ _11572_/X sky130_fd_sc_hd__a311o_1
XANTENNA__09987__A2 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10046__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13311_ _13311_/CLK _13311_/D vssd1 vssd1 vccd1 vccd1 hold287/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10523_ _10523_/A _10523_/B _10523_/C _10524_/B vssd1 vssd1 vccd1 vccd1 _10523_/Y
+ sky130_fd_sc_hd__nor4b_1
XFILLER_0_9_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13242_ _13243_/CLK hold175/X vssd1 vssd1 vccd1 vccd1 hold209/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__09739__A2 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10454_ _10459_/A vssd1 vssd1 vccd1 vccd1 _10454_/Y sky130_fd_sc_hd__inv_2
X_13173_ hold171/X hold137/X _13179_/A _13172_/X vssd1 vssd1 vccd1 vccd1 hold172/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12743__A1 _10281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10385_ _09145_/X _09176_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _10385_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07277__B _07277_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12124_ hold183/A _12124_/B _12186_/B vssd1 vssd1 vccd1 vccd1 _12124_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08175__A1 _08774_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08389__A _10453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ _11197_/S _10111_/Y _12053_/X _12054_/Y vssd1 vssd1 vccd1 vccd1 _12055_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08175__B2 _08774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11006_ _11006_/A _11006_/B vssd1 vssd1 vccd1 vccd1 _11007_/B sky130_fd_sc_hd__nor2_1
X_12957_ hold41/X _13170_/B _12980_/A2 _07134_/A vssd1 vssd1 vccd1 vccd1 _12958_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12888_ _13157_/A _13158_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _13162_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_90_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07740__B _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11908_ reg1_val[23] curr_PC[23] vssd1 vssd1 vccd1 vccd1 _11910_/A sky130_fd_sc_hd__and2_1
XFILLER_0_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11839_ _07111_/B _11923_/A2 _10377_/B reg1_val[22] vssd1 vssd1 vccd1 vccd1 _11839_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07989__B2 _07055_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07989__A1 _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08571__B _08572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07030_ _08777_/A _07030_/B vssd1 vssd1 vccd1 vccd1 _07031_/B sky130_fd_sc_hd__or2_1
XFILLER_0_3_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08981_ _08970_/A _08970_/B _08971_/Y vssd1 vssd1 vccd1 vccd1 _08986_/A sky130_fd_sc_hd__a21bo_1
X_07932_ _07932_/A _07932_/B vssd1 vssd1 vccd1 vccd1 _07933_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07863_ _08477_/B fanout82/X _08672_/B _08776_/B1 vssd1 vssd1 vccd1 vccd1 _07864_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07913__A1 _08774_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07913__B2 _08774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06814_ _06705_/A _06812_/Y _06813_/Y vssd1 vssd1 vccd1 vccd1 _06814_/Y sky130_fd_sc_hd__o21ai_1
X_09602_ _12736_/A _07278_/B fanout7/X _09772_/A vssd1 vssd1 vccd1 vccd1 _09603_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07794_ _08821_/A _07322_/A _07322_/B _08748_/B1 fanout47/X vssd1 vssd1 vccd1 vccd1
+ _07795_/B sky130_fd_sc_hd__o32a_1
X_09533_ _09526_/X _09532_/X _11195_/A vssd1 vssd1 vccd1 vccd1 _09533_/X sky130_fd_sc_hd__mux2_1
X_06745_ reg2_val[6] _06778_/B vssd1 vssd1 vccd1 vccd1 _06745_/X sky130_fd_sc_hd__and2_1
XFILLER_0_64_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06676_ _06676_/A _06676_/B vssd1 vssd1 vccd1 vccd1 _06865_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09464_ _11125_/A _09464_/B vssd1 vssd1 vccd1 vccd1 _09465_/B sky130_fd_sc_hd__xnor2_1
X_08415_ _08415_/A _08415_/B vssd1 vssd1 vccd1 vccd1 _08436_/B sky130_fd_sc_hd__xor2_2
X_09395_ _11089_/A _09394_/A _09212_/Y vssd1 vssd1 vccd1 vccd1 _09395_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08346_ _08854_/B2 _08748_/B1 _12730_/A _08420_/B vssd1 vssd1 vccd1 vccd1 _08347_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07429__B1 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11225__A1 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11225__B2 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08277_ _08443_/A _08277_/B vssd1 vssd1 vccd1 vccd1 _08331_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12284__A _12284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07228_ _08532_/B _10557_/A fanout62/X _07058_/A vssd1 vssd1 vccd1 vccd1 _07229_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_104_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12725__A1 _11147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07159_ _08589_/A _07159_/B vssd1 vssd1 vccd1 vccd1 _07411_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07097__B _07097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10170_ _10171_/B _10170_/B vssd1 vssd1 vccd1 vccd1 _10320_/B sky130_fd_sc_hd__nand2b_1
Xfanout130 _09742_/A vssd1 vssd1 vccd1 vccd1 _08733_/A sky130_fd_sc_hd__buf_12
Xfanout163 _07150_/Y vssd1 vssd1 vccd1 vccd1 _08692_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout152 _12230_/A vssd1 vssd1 vccd1 vccd1 _12124_/B sky130_fd_sc_hd__buf_4
Xfanout141 _06996_/X vssd1 vssd1 vccd1 vccd1 _09888_/B2 sky130_fd_sc_hd__buf_8
Xfanout174 _06963_/Y vssd1 vssd1 vccd1 vccd1 _09478_/B2 sky130_fd_sc_hd__buf_6
XANTENNA__11347__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 _13151_/A2 vssd1 vssd1 vccd1 vccd1 _12721_/B sky130_fd_sc_hd__buf_6
Xfanout185 _08415_/A vssd1 vssd1 vccd1 vccd1 _08773_/A sky130_fd_sc_hd__clkbuf_16
X_12811_ hold295/A hold70/X vssd1 vssd1 vccd1 vccd1 _13087_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__13054__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12742_ hold73/X _12742_/B vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__or2_1
XFILLER_0_96_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10267__A2 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07668__B1 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ reg1_val[23] _12714_/A vssd1 vssd1 vccd1 vccd1 _12678_/D sky130_fd_sc_hd__xnor2_4
XANTENNA__09409__A1 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09409__B2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11624_ _11624_/A _11624_/B vssd1 vssd1 vccd1 vccd1 _11626_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_107_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08672__A _08672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12964__A1 _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08093__B1 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11555_ _11730_/A _11730_/B _11586_/A _12230_/A vssd1 vssd1 vccd1 vccd1 _11555_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11486_ _06674_/Y _11838_/A2 _10638_/B vssd1 vssd1 vccd1 vccd1 _11486_/Y sky130_fd_sc_hd__a21oi_1
X_10506_ _10110_/X _10505_/X _10752_/S vssd1 vssd1 vccd1 vccd1 _10507_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_122_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13225_ _13243_/CLK _13225_/D vssd1 vssd1 vccd1 vccd1 hold187/A sky130_fd_sc_hd__dfxtp_1
X_10437_ fanout32/X _11347_/A _11134_/B2 fanout29/X vssd1 vssd1 vccd1 vccd1 _10438_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11519__A2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12922__A _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12192__A2 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13156_ _13166_/A hold271/X vssd1 vssd1 vccd1 vccd1 _13309_/D sky130_fd_sc_hd__and2_1
XFILLER_0_103_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12641__B _12658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10368_ _10274_/X _10523_/C _10367_/Y vssd1 vssd1 vccd1 vccd1 _10368_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13087_ _13087_/A _13087_/B vssd1 vssd1 vccd1 vccd1 _13088_/B sky130_fd_sc_hd__nand2_1
X_12107_ _12107_/A _12221_/B vssd1 vssd1 vccd1 vccd1 _12107_/Y sky130_fd_sc_hd__nand2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _11853_/A _10299_/B vssd1 vssd1 vccd1 vccd1 _10303_/A sky130_fd_sc_hd__xor2_1
X_12038_ _11890_/A _12101_/A _12101_/B vssd1 vssd1 vccd1 vccd1 _12038_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08200_ _08201_/A _08201_/B vssd1 vssd1 vccd1 vccd1 _08202_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11207__A1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06882__A1 _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ _09180_/A curr_PC[0] vssd1 vssd1 vccd1 vccd1 _09180_/X sky130_fd_sc_hd__or2_1
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08084__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08131_ _08773_/A _08131_/B vssd1 vssd1 vccd1 vccd1 _08198_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08062_ _08062_/A _08062_/B vssd1 vssd1 vccd1 vccd1 _08066_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_71_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10966__B1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07013_ reg1_val[11] _07013_/B vssd1 vssd1 vccd1 vccd1 _08232_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout106_A _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12551__B _12551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07926__A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08964_ _08960_/A _08960_/B _08958_/X vssd1 vssd1 vccd1 vccd1 _08978_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08139__B2 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08139__A1 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07915_ _07919_/A _07919_/B vssd1 vssd1 vccd1 vccd1 _07915_/Y sky130_fd_sc_hd__nor2_1
X_08895_ _08861_/A _08861_/B _08860_/A vssd1 vssd1 vccd1 vccd1 _08902_/A sky130_fd_sc_hd__o21ai_1
X_07846_ _07812_/B _07846_/B vssd1 vssd1 vccd1 vccd1 _07847_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08757__A _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07777_ _09452_/A _07777_/B vssd1 vssd1 vccd1 vccd1 _07788_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12279__A _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11183__A _11379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06728_ _10638_/A _06728_/B vssd1 vssd1 vccd1 vccd1 _10621_/A sky130_fd_sc_hd__nand2_2
X_09516_ _10246_/S _09360_/X _09211_/B vssd1 vssd1 vccd1 vccd1 _09517_/A sky130_fd_sc_hd__o21ai_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11997__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09447_ _08532_/B _07132_/Y fanout22/X _07058_/A vssd1 vssd1 vccd1 vccd1 _09448_/B
+ sky130_fd_sc_hd__o22a_1
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06659_ reg1_val[21] _07052_/B vssd1 vssd1 vccd1 vccd1 _06660_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09378_ _13218_/Q hold211/A _11820_/A _12290_/C1 vssd1 vssd1 vccd1 vccd1 _09379_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_47_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08329_ _08329_/A _08329_/B vssd1 vssd1 vccd1 vccd1 _08330_/B sky130_fd_sc_hd__or2_1
XANTENNA__08075__B1 _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12726__B _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout19_A _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10527__A _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07822__B1 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11340_ _11340_/A _11340_/B vssd1 vssd1 vccd1 vccd1 _11342_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_22_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08378__A1 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13010_ _06965_/C _13020_/B2 hold125/X vssd1 vssd1 vccd1 vccd1 _13275_/D sky130_fd_sc_hd__o21a_1
X_11271_ _11272_/B _11272_/A vssd1 vssd1 vccd1 vccd1 _11369_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__08378__B2 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10222_ _10223_/A _10223_/B vssd1 vssd1 vccd1 vccd1 _10222_/X sky130_fd_sc_hd__or2_1
XFILLER_0_30_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13049__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11921__A2 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10153_ _10658_/A _10153_/B vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_100_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11134__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10084_ _10084_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10085_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07889__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10986_ hold274/A _10986_/B vssd1 vssd1 vccd1 vccd1 _11198_/C sky130_fd_sc_hd__or2_1
XFILLER_0_85_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10645__C1 _10644_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12725_ _11147_/B _12781_/A2 hold34/X _12946_/A vssd1 vssd1 vccd1 vccd1 hold35/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12656_ reg1_val[20] _12714_/A vssd1 vssd1 vccd1 vccd1 _12678_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_194 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12587_ reg1_val[6] _12588_/B vssd1 vssd1 vccd1 vccd1 _12589_/A sky130_fd_sc_hd__nor2_1
X_11607_ _11709_/A _11607_/B vssd1 vssd1 vccd1 vccd1 _11612_/A sky130_fd_sc_hd__or2_1
XANTENNA__06634__B _12598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10412__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11538_ _11539_/A _11539_/B vssd1 vssd1 vccd1 vccd1 _11538_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_20_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11469_ _06683_/X _11382_/X _06685_/B vssd1 vssd1 vccd1 vccd1 _11470_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_110_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13208_ _13305_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__07746__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__B1 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13139_ _13139_/A _13139_/B vssd1 vssd1 vccd1 vccd1 _13140_/B sky130_fd_sc_hd__nand2_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07700_ _07700_/A _07700_/B vssd1 vssd1 vccd1 vccd1 _08983_/B sky130_fd_sc_hd__xnor2_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08680_ _08821_/A _08680_/B vssd1 vssd1 vccd1 vccd1 _08685_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09333__A3 _10230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10900__A _12255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07631_ _07631_/A _07631_/B vssd1 vssd1 vccd1 vccd1 _07632_/B sky130_fd_sc_hd__nand2_1
X_07562_ _07562_/A _07562_/B _07562_/C _07562_/D vssd1 vssd1 vccd1 vccd1 _07563_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_76_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09301_ _09302_/A _09302_/B _09302_/C _09302_/D vssd1 vssd1 vccd1 vccd1 _09301_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07493_ _07494_/B _07590_/A vssd1 vssd1 vccd1 vccd1 _07495_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_29_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11731__A _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09232_ _09232_/A _09232_/B vssd1 vssd1 vccd1 vccd1 _09236_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09163_ reg1_val[17] reg1_val[14] _09173_/S vssd1 vssd1 vccd1 vccd1 _09163_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08114_ _08112_/A _08112_/B _08113_/Y vssd1 vssd1 vccd1 vccd1 _08118_/B sky130_fd_sc_hd__a21bo_2
X_09094_ _08932_/A _08932_/B _08963_/A _08963_/B vssd1 vssd1 vccd1 vccd1 _09094_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_44_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08045_ _08050_/A _08050_/B vssd1 vssd1 vccd1 vccd1 _08045_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_102_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07280__B2 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07280__A1 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13105__B2 _13146_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09996_ _11381_/A _09965_/Y _09966_/X _09995_/X _09964_/X vssd1 vssd1 vccd1 vccd1
+ _09996_/X sky130_fd_sc_hd__a311o_1
X_08947_ _08914_/A _08914_/C _08914_/B vssd1 vssd1 vccd1 vccd1 _08957_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08878_ _08878_/A _08878_/B vssd1 vssd1 vccd1 vccd1 _08880_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10810__A _10811_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07829_ _07829_/A _07829_/B _07829_/C vssd1 vssd1 vccd1 vccd1 _07844_/A sky130_fd_sc_hd__nand3_1
XANTENNA__07391__A _08544_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11419__A1 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10840_ _10842_/A _10842_/B vssd1 vssd1 vccd1 vccd1 _10840_/X sky130_fd_sc_hd__and2_1
XANTENNA__11419__B2 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08835__A2 _08672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10771_ curr_PC[11] _10887_/C vssd1 vssd1 vccd1 vccd1 _10772_/B sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_4_5_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12510_ _12515_/C _12510_/B vssd1 vssd1 vccd1 vccd1 new_PC[19] sky130_fd_sc_hd__xnor2_4
XFILLER_0_82_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12441_ _12450_/A _12441_/B vssd1 vssd1 vccd1 vccd1 _12443_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12372_ _12357_/A _09194_/Y _12370_/X _10638_/B _12371_/X vssd1 vssd1 vccd1 vccd1
+ _12372_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_50_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11323_ _11499_/A _11323_/B vssd1 vssd1 vccd1 vccd1 _11325_/B sky130_fd_sc_hd__xor2_1
X_11254_ _11356_/B _11254_/B vssd1 vssd1 vccd1 vccd1 _11256_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08220__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10205_ _10206_/A _10206_/B _10206_/C vssd1 vssd1 vccd1 vccd1 _10207_/A sky130_fd_sc_hd__o21a_1
X_11185_ _06705_/A _11080_/Y _06704_/B vssd1 vssd1 vccd1 vccd1 _11185_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08771__A1 _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10136_ _10108_/Y _10109_/X _10135_/Y vssd1 vssd1 vccd1 vccd1 _10136_/Y sky130_fd_sc_hd__a21oi_1
X_10067_ _10169_/A _10067_/B vssd1 vssd1 vccd1 vccd1 _10069_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10866__C1 _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_max_cap119_A _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07326__A2 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10330__B2 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10330__A1 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10881__A2 _09188_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10969_ _12131_/A _09059_/A _09059_/B _11381_/A vssd1 vssd1 vccd1 vccd1 _10969_/Y
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_85_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12708_ reg1_val[30] _12708_/B vssd1 vssd1 vccd1 vccd1 _12709_/B sky130_fd_sc_hd__or2_1
XFILLER_0_31_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12639_ _12639_/A _12639_/B _12639_/C vssd1 vssd1 vccd1 vccd1 _12640_/B sky130_fd_sc_hd__and3_2
XFILLER_0_26_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold205 hold205/A vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold249 hold249/A vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 hold238/A vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09850_ _09850_/A _09850_/B vssd1 vssd1 vccd1 vccd1 _09850_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__11429__C fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _08801_/A _08801_/B _08801_/C vssd1 vssd1 vccd1 vccd1 _08801_/X sky130_fd_sc_hd__and3_1
X_06993_ _06993_/A _06993_/B vssd1 vssd1 vccd1 vccd1 _06994_/B sky130_fd_sc_hd__nor2_1
X_09781_ _09781_/A _09781_/B vssd1 vssd1 vccd1 vccd1 _09795_/A sky130_fd_sc_hd__xnor2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _08348_/B _12752_/A fanout84/X _07181_/Y vssd1 vssd1 vccd1 vccd1 _08733_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08663_ _08664_/A _08664_/B vssd1 vssd1 vccd1 vccd1 _08663_/X sky130_fd_sc_hd__and2_1
XANTENNA__08514__A1 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08514__B2 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout173_A _08232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08594_ _08593_/X _08594_/B vssd1 vssd1 vccd1 vccd1 _09514_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_49_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07614_ _07615_/A _07615_/B vssd1 vssd1 vccd1 vccd1 _09226_/A sky130_fd_sc_hd__nand2b_1
X_07545_ _10144_/B2 _09295_/A _10433_/A _08681_/A vssd1 vssd1 vccd1 vccd1 _07546_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07476_ _07234_/B _07237_/B _07234_/A vssd1 vssd1 vccd1 vccd1 _07479_/B sky130_fd_sc_hd__o21ba_1
X_09215_ _12362_/A vssd1 vssd1 vccd1 vccd1 _09215_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13023__B1 _13151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09146_ _09130_/X _09145_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _09146_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12377__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09077_ _09077_/A _09077_/B vssd1 vssd1 vccd1 vccd1 _11977_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08450__B1 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08028_ _08443_/A _08028_/B vssd1 vssd1 vccd1 vccd1 _08071_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_102_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout86_A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ hold224/A _10119_/C _12124_/B vssd1 vssd1 vccd1 vccd1 _09980_/B sky130_fd_sc_hd__o21a_1
X_12990_ _07259_/B _12744_/B hold43/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__a21boi_1
X_11941_ _12206_/A _11941_/B vssd1 vssd1 vccd1 vccd1 _11950_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11872_ _11872_/A _11872_/B vssd1 vssd1 vccd1 vccd1 _11873_/B sky130_fd_sc_hd__and2_1
XFILLER_0_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10823_ _10824_/A _10824_/B _10824_/C vssd1 vssd1 vccd1 vccd1 _10825_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12467__A _12626_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10754_ _10752_/X _10753_/X _11831_/S vssd1 vssd1 vccd1 vccd1 _10754_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10685_ _11499_/A _10685_/B vssd1 vssd1 vccd1 vccd1 _10686_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08680__A _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12424_ reg1_val[7] curr_PC[7] _12556_/S vssd1 vssd1 vccd1 vccd1 _12426_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09233__A2 _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11576__B1 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ _06856_/A _12321_/X _09968_/A _06631_/A vssd1 vssd1 vccd1 vccd1 _12355_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11306_ _09115_/X _11196_/Y _11305_/X vssd1 vssd1 vccd1 vccd1 _11306_/Y sky130_fd_sc_hd__o21ai_1
X_12286_ _09842_/B _12337_/B hold244/A vssd1 vssd1 vccd1 vccd1 _12286_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11237_ _10553_/A _12150_/B _12776_/A fanout33/X vssd1 vssd1 vccd1 vccd1 _11238_/B
+ sky130_fd_sc_hd__o22a_1
X_11168_ _11169_/A _11169_/B vssd1 vssd1 vccd1 vccd1 _11274_/B sky130_fd_sc_hd__and2b_1
X_10119_ hold189/A hold224/A _10119_/C vssd1 vssd1 vccd1 vccd1 _10252_/B sky130_fd_sc_hd__or3_1
XFILLER_0_89_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11099_ reg1_val[14] _11099_/B vssd1 vssd1 vccd1 vccd1 _11099_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_117_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08855__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07330_ _07479_/A _07330_/B vssd1 vssd1 vccd1 vccd1 _07349_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_45_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09000_ _09000_/A _09000_/B vssd1 vssd1 vccd1 vccd1 _09001_/B sky130_fd_sc_hd__nand2_2
X_07261_ _11429_/A _07261_/B vssd1 vssd1 vccd1 vccd1 _07261_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_45_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07192_ _07192_/A _07192_/B vssd1 vssd1 vccd1 vccd1 _07192_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11031__A2 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07235__B2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07235__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10790__B2 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10790__A1 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09902_ _10894_/A _09902_/B vssd1 vssd1 vccd1 vccd1 _09911_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_1_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09833_ _09153_/X _09175_/X _10249_/S vssd1 vssd1 vccd1 vccd1 _10865_/B sky130_fd_sc_hd__mux2_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout290_A _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06761__A3 _12583_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09764_ _09764_/A fanout9/X vssd1 vssd1 vccd1 vccd1 _09764_/Y sky130_fd_sc_hd__nor2_1
X_06976_ reg1_val[20] _07087_/B _12658_/B _07105_/A vssd1 vssd1 vccd1 vccd1 _06978_/B
+ sky130_fd_sc_hd__o31a_4
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08715_ _08715_/A _08715_/B vssd1 vssd1 vccd1 vccd1 _08717_/B sky130_fd_sc_hd__xnor2_1
X_09695_ _06790_/Y _09694_/Y _12322_/S vssd1 vssd1 vccd1 vccd1 _09695_/X sky130_fd_sc_hd__mux2_1
X_08646_ _08775_/A _08646_/B vssd1 vssd1 vccd1 vccd1 _08650_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09360__S _09679_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _08577_/A _08602_/A _08577_/C vssd1 vssd1 vccd1 vccd1 _08577_/X sky130_fd_sc_hd__and3_1
XFILLER_0_49_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07528_ reg1_val[29] reg1_val[30] _07528_/C vssd1 vssd1 vccd1 vccd1 _07528_/X sky130_fd_sc_hd__or3_1
XANTENNA__09463__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07459_ _07459_/A _07459_/B vssd1 vssd1 vccd1 vccd1 _07462_/A sky130_fd_sc_hd__nor2_1
X_10470_ _10349_/A _10349_/B _10347_/X vssd1 vssd1 vccd1 vccd1 _10477_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_122_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12734__B _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11558__B1 _11559_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09129_ _09125_/X _09128_/X _09676_/S vssd1 vssd1 vccd1 vccd1 _09129_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_121_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10535__A _12255_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12140_ fanout19/X fanout15/X fanout6/X _12203_/A vssd1 vssd1 vccd1 vccd1 _12141_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_102_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12071_ _12005_/A _12069_/Y _12136_/B _12068_/X vssd1 vssd1 vccd1 vccd1 dest_val[25]
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11022_ _11853_/A _11022_/B vssd1 vssd1 vccd1 vccd1 _11024_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09923__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ _13256_/Q _12723_/A _13170_/B hold134/X _13066_/A vssd1 vssd1 vccd1 vccd1
+ hold135/A sky130_fd_sc_hd__o221a_1
XFILLER_0_99_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11924_ _06639_/B _11921_/X _11923_/X vssd1 vssd1 vccd1 vccd1 _11924_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06907__B _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11855_ fanout29/X _12301_/A fanout8/X fanout32/X vssd1 vssd1 vccd1 vccd1 _11856_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_55_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11786_ _11786_/A _11786_/B vssd1 vssd1 vccd1 vccd1 _11802_/A sky130_fd_sc_hd__xor2_1
X_10806_ _10807_/A _10807_/B vssd1 vssd1 vccd1 vccd1 _10943_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_27_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10737_ _10650_/X _10774_/B _12223_/B1 vssd1 vssd1 vccd1 vccd1 _10737_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__06671__A2_N _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12407_ _12408_/A _12408_/B _12408_/C vssd1 vssd1 vccd1 vccd1 _12415_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_70_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10668_ _11853_/A _10668_/B vssd1 vssd1 vccd1 vccd1 _10670_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07768__A2 _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08414__B1 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10599_ _10599_/A _10599_/B vssd1 vssd1 vccd1 vccd1 _10600_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_23_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12338_ _09842_/B _12337_/X hold287/A vssd1 vssd1 vccd1 vccd1 _12338_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_50_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12269_ _12312_/B _12270_/B vssd1 vssd1 vccd1 vccd1 _12269_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_37_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06830_ reg1_val[22] _07111_/B vssd1 vssd1 vccd1 vccd1 _06830_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10180__A _10180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06761_ _06783_/A _06649_/A _12583_/B _06759_/X vssd1 vssd1 vccd1 vccd1 _06761_/Y
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__11485__C1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06692_ _12641_/A _07167_/A vssd1 vssd1 vccd1 vccd1 _06693_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_78_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08500_ _08529_/A _08507_/B _08493_/X vssd1 vssd1 vccd1 vccd1 _08524_/B sky130_fd_sc_hd__a21o_1
X_09480_ _09481_/A _09481_/B vssd1 vssd1 vccd1 vccd1 _09480_/X sky130_fd_sc_hd__and2b_1
X_08431_ _09008_/A _09008_/B vssd1 vssd1 vccd1 vccd1 _08431_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08362_ _08362_/A _08362_/B vssd1 vssd1 vccd1 vccd1 _08406_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11788__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09445__A2 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08293_ _08296_/A _08296_/B vssd1 vssd1 vccd1 vccd1 _08295_/B sky130_fd_sc_hd__nand2_1
X_07313_ _07313_/A _07313_/B vssd1 vssd1 vccd1 vccd1 _10694_/A sky130_fd_sc_hd__nand2_8
XFILLER_0_34_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout136_A _07057_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07244_ _07434_/A _07434_/C _07434_/D _07303_/B vssd1 vssd1 vccd1 vccd1 _07245_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07175_ _07175_/A _07175_/B _07175_/C _07175_/D vssd1 vssd1 vccd1 vccd1 _07303_/C
+ sky130_fd_sc_hd__or4_4
XANTENNA_fanout303_A _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07759__A2 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06967__B1 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07664__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09905__B1 _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout301 reg1_val[1] vssd1 vssd1 vccd1 vccd1 _12563_/A sky130_fd_sc_hd__clkbuf_16
XANTENNA__09381__A1 _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07392__B1 _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ _09816_/A _10229_/A vssd1 vssd1 vccd1 vccd1 _09816_/X sky130_fd_sc_hd__or2_1
X_06959_ _06960_/A _12078_/A vssd1 vssd1 vccd1 vccd1 _06959_/Y sky130_fd_sc_hd__nor2_1
X_09747_ _09748_/A _09748_/B vssd1 vssd1 vccd1 vccd1 _09881_/B sky130_fd_sc_hd__nor2_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10818__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10279__B1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ _09363_/X _09365_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09678_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08495__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout49_A _07301_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ _08258_/Y _08628_/X _08210_/X vssd1 vssd1 vccd1 vccd1 _08629_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11640_ _10855_/B _11279_/Y _11637_/Y _11639_/X vssd1 vssd1 vccd1 vccd1 _12216_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11571_ _12119_/B1 _11664_/B hold280/A vssd1 vssd1 vccd1 vccd1 _11571_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11779__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13310_ _13310_/CLK _13310_/D vssd1 vssd1 vccd1 vccd1 hold244/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10522_ _12005_/A _10401_/X _10493_/X _10521_/X vssd1 vssd1 vccd1 vccd1 dest_val[9]
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_107_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13241_ _13241_/CLK _13241_/D vssd1 vssd1 vccd1 vccd1 hold173/A sky130_fd_sc_hd__dfxtp_1
X_10453_ _10453_/A _10453_/B vssd1 vssd1 vccd1 vccd1 _10459_/A sky130_fd_sc_hd__xnor2_2
X_13172_ hold171/X _12721_/B _12715_/Y _06537_/A vssd1 vssd1 vccd1 vccd1 _13172_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12743__A2 _12980_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ _10373_/A _11838_/A2 _10378_/X _10383_/Y vssd1 vssd1 vccd1 vccd1 _10384_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ _12124_/B _12186_/B hold183/A vssd1 vssd1 vccd1 vccd1 _12123_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_20_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12054_ _12053_/A _12053_/B _11197_/S vssd1 vssd1 vccd1 vccd1 _12054_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__08175__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ _11005_/A _11005_/B _11005_/C vssd1 vssd1 vccd1 vccd1 _11006_/B sky130_fd_sc_hd__and3_1
XFILLER_0_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12956_ _13169_/A hold150/X vssd1 vssd1 vccd1 vccd1 hold151/A sky130_fd_sc_hd__and2_1
X_12887_ hold21/X hold270/X vssd1 vssd1 vccd1 vccd1 _13157_/B sky130_fd_sc_hd__nand2b_1
X_11907_ _11906_/A _11906_/B _11906_/Y _12228_/B1 vssd1 vssd1 vccd1 vccd1 _11907_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11838_ _06645_/A _11838_/A2 _10638_/B vssd1 vssd1 vccd1 vccd1 _11838_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07989__A2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07749__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11769_ _07389_/B _12150_/B _12776_/A _12205_/A vssd1 vssd1 vccd1 vccd1 _11770_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11942__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12390__A _12568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08980_ _08975_/A _08975_/B _08973_/X vssd1 vssd1 vccd1 vccd1 _08989_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_11_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07931_ _07848_/A _07848_/B _07848_/C vssd1 vssd1 vccd1 vccd1 _07933_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07862_ _08773_/A _07862_/B vssd1 vssd1 vccd1 vccd1 _07904_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07913__A2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06813_ _07192_/A reg1_val[14] vssd1 vssd1 vccd1 vccd1 _06813_/Y sky130_fd_sc_hd__nand2b_1
X_09601_ _09472_/A _09472_/B _09468_/Y vssd1 vssd1 vccd1 vccd1 _09605_/A sky130_fd_sc_hd__a21oi_2
X_07793_ _08836_/A _07793_/B vssd1 vssd1 vccd1 vccd1 _07797_/A sky130_fd_sc_hd__xnor2_1
X_09532_ _09528_/X _09531_/X _11089_/A vssd1 vssd1 vccd1 vccd1 _09532_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06744_ _06742_/Y _06744_/B vssd1 vssd1 vccd1 vccd1 _06866_/D sky130_fd_sc_hd__nand2b_2
X_06675_ reg1_val[18] _07023_/A vssd1 vssd1 vccd1 vccd1 _06676_/B sky130_fd_sc_hd__nor2_1
XANTENNA_fanout253_A _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09463_ _10553_/B fanout95/X fanout54/X fanout69/X vssd1 vssd1 vccd1 vccd1 _09464_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_80_50 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08414_ _12734_/A _08532_/B _07058_/A _08819_/B2 vssd1 vssd1 vccd1 vccd1 _08415_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09394_ _09394_/A vssd1 vssd1 vccd1 vccd1 _09394_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_19_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08345_ _08345_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08365_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_58_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07429__A1 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07429__B2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11225__A2 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08276_ _08692_/A2 fanout82/X _08672_/B _08692_/B1 vssd1 vssd1 vccd1 vccd1 _08277_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07659__A _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07227_ _07225_/A _07225_/B _07226_/X vssd1 vssd1 vccd1 vccd1 _07354_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12725__A2 _12781_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07158_ _08588_/B _10677_/A _09273_/A1 fanout58/X vssd1 vssd1 vccd1 vccd1 _07159_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09051__B1 _10370_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07089_ reg1_val[29] _07165_/A _07528_/C vssd1 vssd1 vccd1 vccd1 _07090_/B sky130_fd_sc_hd__and3_1
Xfanout131 _09742_/A vssd1 vssd1 vccd1 vccd1 _08853_/A sky130_fd_sc_hd__buf_8
Xfanout120 _10169_/A vssd1 vssd1 vccd1 vccd1 _12022_/A sky130_fd_sc_hd__clkbuf_16
XFILLER_0_100_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout142 _10064_/B2 vssd1 vssd1 vccd1 vccd1 _08841_/B2 sky130_fd_sc_hd__buf_6
Xfanout153 _12230_/A vssd1 vssd1 vccd1 vccd1 _11820_/A sky130_fd_sc_hd__buf_2
Xfanout164 _07116_/X vssd1 vssd1 vccd1 vccd1 _09618_/A1 sky130_fd_sc_hd__buf_4
Xfanout197 _06891_/Y vssd1 vssd1 vccd1 vccd1 _13151_/A2 sky130_fd_sc_hd__buf_4
Xfanout175 _06963_/Y vssd1 vssd1 vccd1 vccd1 _08819_/B2 sky130_fd_sc_hd__clkbuf_8
XANTENNA__06707__A3 _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout186 _09452_/A vssd1 vssd1 vccd1 vccd1 _10458_/A sky130_fd_sc_hd__clkbuf_16
X_12810_ hold282/X hold65/X vssd1 vssd1 vccd1 vccd1 _13092_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12110__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12741_ _10149_/A _12980_/A2 hold57/X _13086_/A vssd1 vssd1 vccd1 vccd1 _13192_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09114__A _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07668__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07668__B2 _12768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12669_/B _12671_/B _12667_/X vssd1 vssd1 vccd1 vccd1 _12674_/A sky130_fd_sc_hd__a21o_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09409__A2 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11623_ _11624_/B _11624_/A vssd1 vssd1 vccd1 vccd1 _11623_/X sky130_fd_sc_hd__and2b_1
XANTENNA__12475__A _12632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08672__B _08672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10424__B1 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08093__A1 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08093__B2 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11554_ _11635_/B _11554_/B vssd1 vssd1 vccd1 vccd1 _11586_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07569__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11485_ hold289/A _12119_/B1 _11570_/B _11484_/Y _11400_/A vssd1 vssd1 vccd1 vccd1
+ _11490_/B sky130_fd_sc_hd__a311o_1
XFILLER_0_80_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10505_ _09354_/X _09368_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _10505_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_122_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13224_ _13243_/CLK hold230/X vssd1 vssd1 vccd1 vccd1 _13224_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__09784__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10436_ _10435_/B _10435_/C _10435_/A vssd1 vssd1 vccd1 vccd1 _10446_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13155_ hold270/X _13165_/A2 _13154_/X _13168_/A2 vssd1 vssd1 vccd1 vccd1 hold271/A
+ sky130_fd_sc_hd__a22o_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10367_ _10274_/X _10523_/C _09110_/X vssd1 vssd1 vccd1 vccd1 _10367_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13086_ _13086_/A _13086_/B vssd1 vssd1 vccd1 vccd1 _13294_/D sky130_fd_sc_hd__and2_1
X_12106_ _12107_/A _12221_/B vssd1 vssd1 vccd1 vccd1 _12106_/X sky130_fd_sc_hd__or2_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10553_/A _11431_/A _11347_/A fanout33/X vssd1 vssd1 vccd1 vccd1 _10299_/B
+ sky130_fd_sc_hd__o22a_1
X_12037_ _12102_/B _12102_/C vssd1 vssd1 vccd1 vccd1 _12163_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_18_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12939_ hold200/A _12947_/A2 _12947_/B1 hold192/X vssd1 vssd1 vccd1 vccd1 hold193/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08856__B1 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08130_ _08772_/B2 _08672_/B _08835_/B1 _08772_/A2 vssd1 vssd1 vccd1 vccd1 _08131_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_83_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_248 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08084__B2 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08084__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12955__A2 _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08061_ _08069_/B _08069_/A vssd1 vssd1 vccd1 vccd1 _08062_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07012_ reg1_val[10] _07027_/B _07105_/A vssd1 vssd1 vccd1 vccd1 _07013_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_70_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08963_ _08963_/A _08963_/B vssd1 vssd1 vccd1 vccd1 _09103_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__08139__A2 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07914_ _08775_/A _07914_/B vssd1 vssd1 vccd1 vccd1 _07919_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12340__B1 _12327_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08894_ _08894_/A _08894_/B vssd1 vssd1 vccd1 vccd1 _08914_/A sky130_fd_sc_hd__xnor2_1
X_07845_ _07844_/A _07844_/C _07844_/B vssd1 vssd1 vccd1 vccd1 _07848_/B sky130_fd_sc_hd__a21oi_2
X_07776_ _08477_/B _12752_/A fanout84/X _08776_/B1 vssd1 vssd1 vccd1 vccd1 _07777_/B
+ sky130_fd_sc_hd__o22a_1
X_06727_ reg1_val[10] _07319_/A vssd1 vssd1 vccd1 vccd1 _06728_/B sky130_fd_sc_hd__nand2_1
X_09515_ _08595_/B _09035_/B _09515_/S vssd1 vssd1 vccd1 vccd1 _09515_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10654__B1 fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09446_ _10658_/A _09446_/B vssd1 vssd1 vccd1 vccd1 _09450_/A sky130_fd_sc_hd__xnor2_1
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08773__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06658_ _07052_/B reg1_val[21] vssd1 vssd1 vccd1 vccd1 _11756_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09377_ hold211/A _11820_/A _13218_/Q vssd1 vssd1 vccd1 vccd1 _09379_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__12295__A _12295_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06589_ _12250_/A reg1_val[28] vssd1 vssd1 vccd1 vccd1 _06591_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_19_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08328_ _08328_/A _08328_/B vssd1 vssd1 vccd1 vccd1 _08329_/B sky130_fd_sc_hd__and2_1
XANTENNA__08075__B2 _08544_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08075__A1 _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07389__A _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10406__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08259_ _08259_/A _08259_/B vssd1 vssd1 vccd1 vccd1 _09070_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_104_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10527__B fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12742__B _12742_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08378__A2 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11270_ _11270_/A _11270_/B vssd1 vssd1 vccd1 vccd1 _11272_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06740__B _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ _10223_/A _10223_/B vssd1 vssd1 vccd1 vccd1 _10221_/X sky130_fd_sc_hd__and2_1
X_10152_ _10527_/A _12782_/A fanout20/X _10452_/B2 vssd1 vssd1 vccd1 vccd1 _10153_/B
+ sky130_fd_sc_hd__o22a_1
X_10083_ _10084_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10083_/Y sky130_fd_sc_hd__nor2_1
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07852__A _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__B2 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__A1 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__B2 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12724_ hold33/X _12778_/B vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__or2_1
X_10985_ hold215/A _12187_/A1 _11201_/C _12290_/C1 vssd1 vssd1 vccd1 vccd1 _10985_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08683__A _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06915__B _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12655_ _12655_/A _12657_/D vssd1 vssd1 vccd1 vccd1 loadstore_address[19] sky130_fd_sc_hd__xnor2_4
XFILLER_0_53_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12586_ _12585_/A _12582_/Y _12584_/B vssd1 vssd1 vccd1 vccd1 _12590_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11606_ _11605_/B _11606_/B vssd1 vssd1 vccd1 vccd1 _11607_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_123_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11537_ _11446_/A _11445_/B _11443_/X vssd1 vssd1 vccd1 vccd1 _11539_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11468_ _11468_/A _11468_/B vssd1 vssd1 vccd1 vccd1 _11468_/Y sky130_fd_sc_hd__xnor2_1
Xmax_cap128 _07894_/A vssd1 vssd1 vccd1 vccd1 _10184_/A sky130_fd_sc_hd__buf_4
XFILLER_0_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11399_ _11398_/B _11483_/B hold260/A vssd1 vssd1 vccd1 vccd1 _11400_/C sky130_fd_sc_hd__a21oi_1
X_13207_ _13303_/CLK _13207_/D vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09566__B2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09566__A1 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10419_ _10420_/A _10420_/B _10420_/C vssd1 vssd1 vccd1 vccd1 _10421_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__10453__A _10453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13138_ _13147_/A hold263/X vssd1 vssd1 vccd1 vccd1 _13305_/D sky130_fd_sc_hd__and2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13069_ hold272/X _13068_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13069_/X sky130_fd_sc_hd__mux2_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07630_ _08941_/A _08941_/B _07627_/X vssd1 vssd1 vccd1 vccd1 _07690_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_45_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07561_ _07562_/A _07562_/B _07562_/C _07562_/D vssd1 vssd1 vccd1 vccd1 _07561_/X
+ sky130_fd_sc_hd__o22a_1
X_09300_ _10559_/A _09300_/B vssd1 vssd1 vccd1 vccd1 _09302_/D sky130_fd_sc_hd__nor2_1
XFILLER_0_118_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07492_ _07459_/B _07462_/B _07459_/A vssd1 vssd1 vccd1 vccd1 _07494_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09231_ _10306_/A _09231_/B vssd1 vssd1 vccd1 vccd1 _09232_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_90_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09162_ reg1_val[16] reg1_val[15] _09172_/S vssd1 vssd1 vccd1 vccd1 _09162_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09254__B1 _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08113_ _08121_/B _08121_/A vssd1 vssd1 vccd1 vccd1 _08113_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_114_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13050__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09093_ _09092_/A _09092_/B _12230_/B vssd1 vssd1 vccd1 vccd1 _12278_/B sky130_fd_sc_hd__o21bai_2
XFILLER_0_44_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08044_ _08107_/A _08107_/B _08040_/X vssd1 vssd1 vccd1 vccd1 _08050_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_114_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07280__A2 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12562__B _12563_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09557__A1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07568__B1 fanout26/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13105__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09995_ _09192_/Y _09970_/Y _09972_/Y _12373_/A1 _09994_/X vssd1 vssd1 vccd1 vccd1
+ _09995_/X sky130_fd_sc_hd__a221o_1
X_08946_ _08946_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _08959_/A sky130_fd_sc_hd__xor2_4
X_08877_ _08878_/A _08878_/B vssd1 vssd1 vccd1 vccd1 _08886_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10810__B _12255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07828_ _07825_/B _07825_/C _07825_/A vssd1 vssd1 vccd1 vccd1 _07829_/C sky130_fd_sc_hd__a21o_1
XANTENNA__07391__B _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11419__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ _08841_/B2 _08217_/B fanout55/X _08837_/B2 vssd1 vssd1 vccd1 vccd1 _07760_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10770_ curr_PC[11] _10887_/C vssd1 vssd1 vccd1 vccd1 _10770_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout31_A fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09429_ _07553_/A fanout46/X fanout12/X _10927_/A vssd1 vssd1 vccd1 vccd1 _09430_/B
+ sky130_fd_sc_hd__o22a_1
X_12440_ _12603_/B _12440_/B vssd1 vssd1 vccd1 vccd1 _12441_/B sky130_fd_sc_hd__or2_1
XANTENNA__06735__B _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13041__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12371_ reg1_val[31] _12370_/B wire201/X _12369_/Y vssd1 vssd1 vccd1 vccd1 _12371_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11322_ _12301_/A fanout13/X fanout8/X _10557_/B vssd1 vssd1 vccd1 vccd1 _11323_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11253_ _11252_/B _11253_/B vssd1 vssd1 vccd1 vccd1 _11254_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08220__A1 _08774_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10204_ _10204_/A _10204_/B vssd1 vssd1 vccd1 vccd1 _10206_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__08220__B2 _08774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11184_ _11184_/A _11184_/B _11183_/X vssd1 vssd1 vccd1 vccd1 _11184_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_100_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10135_ _09115_/X _10111_/Y _10134_/X vssd1 vssd1 vccd1 vccd1 _10135_/Y sky130_fd_sc_hd__o21ai_2
X_10066_ _08821_/B fanout83/X fanout81/X fanout36/X vssd1 vssd1 vccd1 vccd1 _10067_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09720__B2 _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__A1 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10330__A2 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10968_ _12131_/A _09059_/A _09059_/B vssd1 vssd1 vccd1 vccd1 _10968_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_85_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12707_ reg1_val[30] _12708_/B vssd1 vssd1 vccd1 vccd1 _12707_/X sky130_fd_sc_hd__and2_1
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12638_ _12639_/A _12639_/B _12639_/C vssd1 vssd1 vccd1 vccd1 _12640_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10899_ _11347_/A fanout27/X _12205_/A _11134_/B2 vssd1 vssd1 vccd1 vccd1 _10900_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13032__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12569_ _12567_/Y _12569_/B vssd1 vssd1 vccd1 vccd1 _12570_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_26_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold206 hold206/A vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 hold237/X vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold239 hold239/A vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold228 hold228/A vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _08800_/A _08800_/B vssd1 vssd1 vccd1 vccd1 _08801_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08588__A _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06992_ _06993_/A _06993_/B vssd1 vssd1 vccd1 vccd1 _07595_/A sky130_fd_sc_hd__and2_1
X_09780_ _09780_/A _09780_/B vssd1 vssd1 vccd1 vccd1 _09781_/B sky130_fd_sc_hd__xnor2_2
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08731_ _08731_/A _08731_/B vssd1 vssd1 vccd1 vccd1 _08754_/A sky130_fd_sc_hd__xor2_1
XANTENNA__07970__B1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08662_ _10565_/A _08662_/B vssd1 vssd1 vccd1 vccd1 _08664_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__08514__A2 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07613_ _07354_/A _07354_/B _07352_/X vssd1 vssd1 vccd1 vccd1 _07615_/B sky130_fd_sc_hd__a21bo_2
XANTENNA_fanout166_A _07110_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08593_ reg1_val[0] _09283_/A _08544_/C _09362_/S vssd1 vssd1 vccd1 vccd1 _08593_/X
+ sky130_fd_sc_hd__a22o_1
X_07544_ _10169_/A _07544_/B vssd1 vssd1 vccd1 vccd1 _07548_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12557__B _12557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11282__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07475_ _07475_/A _07475_/B vssd1 vssd1 vccd1 vccd1 _07482_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06555__B _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09214_ _09214_/A _11195_/B _11195_/C vssd1 vssd1 vccd1 vccd1 _12362_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_8_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13023__A1 _06537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11585__A1 _12382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09145_ _09137_/X _09144_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09145_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09076_ _09076_/A _09076_/B vssd1 vssd1 vccd1 vccd1 _09076_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__08450__B2 _08477_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08450__A1 _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08027_ _07149_/Y _07179_/A _11012_/A _07155_/X vssd1 vssd1 vccd1 vccd1 _08028_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09978_ _09975_/X _09977_/X _10251_/S vssd1 vssd1 vccd1 vccd1 _09978_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07961__B1 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ _08929_/A _08929_/B vssd1 vssd1 vccd1 vccd1 _08930_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_99_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11940_ fanout27/X _12203_/A _12150_/A _12205_/A vssd1 vssd1 vccd1 vccd1 _11941_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09106__B _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11871_ _11872_/A _11872_/B vssd1 vssd1 vccd1 vccd1 _11952_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09466__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10822_ _10925_/A _10925_/B vssd1 vssd1 vccd1 vccd1 _10824_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10753_ _10753_/A _10753_/B vssd1 vssd1 vccd1 vccd1 _10753_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_109_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13014__A1 _07097_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10684_ fanout58/X _10557_/B fanout13/X _11935_/A vssd1 vssd1 vccd1 vccd1 _10685_/B
+ sky130_fd_sc_hd__o22a_1
X_12423_ _12429_/B _12423_/B vssd1 vssd1 vccd1 vccd1 new_PC[6] sky130_fd_sc_hd__and2_4
XANTENNA__08680__B _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12354_ _12353_/A _12353_/B _09109_/Y vssd1 vssd1 vccd1 vccd1 _12354_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_35_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11305_ _09183_/Y _11208_/X _11303_/Y _11304_/X vssd1 vssd1 vccd1 vccd1 _11305_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12285_ hold270/A _12285_/B vssd1 vssd1 vccd1 vccd1 _12337_/B sky130_fd_sc_hd__or2_1
XANTENNA__10000__A1 _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11236_ _11354_/B _11236_/B vssd1 vssd1 vccd1 vccd1 _11256_/A sky130_fd_sc_hd__or2_1
X_11167_ _11167_/A _11167_/B vssd1 vssd1 vccd1 vccd1 _11169_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07952__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10118_ _10752_/S _10116_/X _10117_/X vssd1 vssd1 vccd1 vccd1 _10118_/Y sky130_fd_sc_hd__o21ai_1
X_11098_ hold282/A _11096_/X _11097_/Y vssd1 vssd1 vccd1 vccd1 _11098_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10049_ _10049_/A _10049_/B vssd1 vssd1 vccd1 vccd1 _10050_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12658__A _12658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06656__A _06687_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10178__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07260_ _07261_/B _07260_/B vssd1 vssd1 vccd1 vccd1 _07260_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07191_ _07192_/A _07192_/B vssd1 vssd1 vccd1 vccd1 _11012_/A sky130_fd_sc_hd__xor2_4
XANTENNA__10906__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07235__A2 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09901_ fanout58/X fanout98/X fanout56/X _10557_/A vssd1 vssd1 vccd1 vccd1 _09902_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10790__A2 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09832_ _09830_/X _09831_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _09832_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _10155_/A _09763_/B vssd1 vssd1 vccd1 vccd1 _09766_/B sky130_fd_sc_hd__xnor2_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _08715_/B _08715_/A vssd1 vssd1 vccd1 vccd1 _08722_/A sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout283_A _06898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06975_ _07015_/B _06975_/B vssd1 vssd1 vccd1 vccd1 _10281_/A sky130_fd_sc_hd__xnor2_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09694_ _09694_/A _09694_/B vssd1 vssd1 vccd1 vccd1 _09694_/Y sky130_fd_sc_hd__nor2_1
X_08645_ _12766_/A _08774_/A2 _08774_/B1 fanout70/X vssd1 vssd1 vccd1 vccd1 _08646_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12047__A2 _09079_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08576_ _08577_/A _08577_/C _08602_/A vssd1 vssd1 vccd1 vccd1 _08576_/X sky130_fd_sc_hd__a21o_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07527_ _07527_/A _07527_/B vssd1 vssd1 vccd1 vccd1 _07541_/A sky130_fd_sc_hd__xor2_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07458_ _07458_/A _07458_/B vssd1 vssd1 vccd1 vccd1 _07459_/B sky130_fd_sc_hd__and2_1
XFILLER_0_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07389_ _08588_/A _07389_/B vssd1 vssd1 vccd1 vccd1 _07629_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_45_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09128_ _09126_/X _09127_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09128_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_114_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09059_ _09059_/A _09059_/B _09059_/C vssd1 vssd1 vccd1 vccd1 _11183_/B sky130_fd_sc_hd__and3_1
XFILLER_0_60_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12750__B _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12070_ curr_PC[24] curr_PC[25] _12070_/C vssd1 vssd1 vccd1 vccd1 _12136_/B sky130_fd_sc_hd__and3_1
X_11021_ _10553_/A _11935_/A _12772_/A fanout33/X vssd1 vssd1 vccd1 vccd1 _11022_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10551__A _10551_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__B2 _10553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09923__A1 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12972_ _08773_/A _12742_/B hold122/X vssd1 vssd1 vccd1 vccd1 hold123/A sky130_fd_sc_hd__a21boi_1
XANTENNA__09687__B1 _12361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11923_ _07119_/A _11923_/A2 _10377_/B reg1_val[23] _11922_/Y vssd1 vssd1 vccd1 vccd1
+ _11923_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_59_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11494__B1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11854_ _11938_/A _11854_/B vssd1 vssd1 vccd1 vccd1 _11858_/A sky130_fd_sc_hd__or2_1
X_10805_ _10805_/A _10805_/B vssd1 vssd1 vccd1 vccd1 _10807_/B sky130_fd_sc_hd__xor2_1
X_11785_ _11861_/A _11785_/B vssd1 vssd1 vccd1 vccd1 _11786_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_125_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10736_ _10736_/A _10736_/B vssd1 vssd1 vccd1 vccd1 _10774_/B sky130_fd_sc_hd__or2_1
XFILLER_0_70_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10667_ _10553_/A _11704_/A _11688_/A fanout33/X vssd1 vssd1 vccd1 vccd1 _10668_/B
+ sky130_fd_sc_hd__o22a_1
X_12406_ _12415_/A _12406_/B vssd1 vssd1 vccd1 vccd1 _12408_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08414__A1 _12734_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08414__B2 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10598_ _10599_/A _10599_/B vssd1 vssd1 vccd1 vccd1 _10598_/Y sky130_fd_sc_hd__nor2_1
X_12337_ hold244/A _12337_/B vssd1 vssd1 vccd1 vccd1 _12337_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12268_ _12215_/B _12165_/B _12214_/A _12214_/B _12267_/Y vssd1 vssd1 vccd1 vccd1
+ _12270_/B sky130_fd_sc_hd__a41o_1
XFILLER_0_10_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11219_ _11431_/A fanout15/X fanout6/X _11347_/A vssd1 vssd1 vccd1 vccd1 _11220_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07925__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09390__A2 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12199_ _12301_/A fanout15/X fanout6/X fanout19/X vssd1 vssd1 vccd1 vccd1 _12200_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06760_ _06783_/A _06649_/A _12583_/B _06759_/X vssd1 vssd1 vccd1 vccd1 _06760_/X
+ sky130_fd_sc_hd__a31o_1
X_06691_ _12641_/A _07167_/A vssd1 vssd1 vccd1 vccd1 _06691_/Y sky130_fd_sc_hd__nand2_1
X_08430_ _08430_/A _08430_/B vssd1 vssd1 vccd1 vccd1 _09008_/B sky130_fd_sc_hd__xor2_2
XANTENNA__10400__S _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11237__B1 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08361_ _08390_/A _08363_/B vssd1 vssd1 vccd1 vccd1 _08361_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11788__A1 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08292_ _08290_/A _08290_/B _08291_/X vssd1 vssd1 vccd1 vccd1 _08296_/B sky130_fd_sc_hd__o21bai_2
X_07312_ _07313_/A _07313_/B vssd1 vssd1 vccd1 vccd1 _07312_/X sky130_fd_sc_hd__and2_2
XANTENNA__11788__B2 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06664__B1 _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07243_ _07243_/A _12250_/A vssd1 vssd1 vccd1 vccd1 _07434_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout129_A _09742_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07174_ _07180_/B _07174_/B vssd1 vssd1 vccd1 vccd1 _08348_/B sky130_fd_sc_hd__or2_4
XANTENNA__09602__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06967__A1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10763__A2 wire201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06967__B2 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 reg1_val[0] vssd1 vssd1 vccd1 vccd1 _09180_/A sky130_fd_sc_hd__buf_6
XANTENNA__07916__B1 _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _09504_/X _09657_/X _09658_/X vssd1 vssd1 vccd1 vccd1 _09815_/X sky130_fd_sc_hd__a21o_1
XANTENNA__09381__A2 _12726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06958_ _11780_/A _06965_/C vssd1 vssd1 vccd1 vccd1 _12078_/A sky130_fd_sc_hd__nor2_1
X_09746_ _09746_/A _09746_/B vssd1 vssd1 vccd1 vccd1 _09748_/B sky130_fd_sc_hd__xnor2_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07680__A _08415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09677_ _09211_/A _09676_/X _10249_/S vssd1 vssd1 vccd1 vccd1 _09677_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10279__B2 _07099_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10279__A1 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _08630_/A _08630_/B vssd1 vssd1 vccd1 vccd1 _08628_/X sky130_fd_sc_hd__or2_1
X_06889_ _06752_/A _06572_/X _09199_/B instruction[4] _06888_/Y vssd1 vssd1 vccd1
+ vccd1 _12723_/B sky130_fd_sc_hd__a221oi_2
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08559_ _08559_/A _08559_/B _08559_/C vssd1 vssd1 vccd1 vccd1 _08568_/B sky130_fd_sc_hd__and3_1
XFILLER_0_49_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11779__A1 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11570_ hold289/A _11570_/B vssd1 vssd1 vccd1 vccd1 _11664_/B sky130_fd_sc_hd__or2_1
XFILLER_0_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11779__B2 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10521_ _10494_/Y _10495_/X _10520_/X vssd1 vssd1 vccd1 vccd1 _10521_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13240_ _13241_/CLK hold194/X vssd1 vssd1 vccd1 vccd1 hold226/A sky130_fd_sc_hd__dfxtp_1
X_10452_ _10527_/A fanout18/X fanout9/X _10452_/B2 vssd1 vssd1 vccd1 vccd1 _10453_/B
+ sky130_fd_sc_hd__o22a_1
X_13171_ hold137/X _06537_/A _13179_/A hold138/X vssd1 vssd1 vccd1 vccd1 hold139/A
+ sky130_fd_sc_hd__o211a_1
X_10383_ _10383_/A vssd1 vssd1 vccd1 vccd1 _10383_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12122_ hold209/A _12122_/B vssd1 vssd1 vccd1 vccd1 _12186_/B sky130_fd_sc_hd__or2_1
XFILLER_0_32_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12053_ _12053_/A _12053_/B vssd1 vssd1 vccd1 vccd1 _12053_/X sky130_fd_sc_hd__or2_1
XFILLER_0_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10281__A _10281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ _11005_/A _11005_/B _11005_/C vssd1 vssd1 vccd1 vccd1 _11006_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08580__B1 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__B1 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12955_ hold231/A _12955_/A2 _13168_/B1 hold149/X vssd1 vssd1 vccd1 vccd1 hold150/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11906_ _11906_/A _11906_/B vssd1 vssd1 vccd1 vccd1 _11906_/Y sky130_fd_sc_hd__nand2_1
X_12886_ _13153_/A _12885_/B _12885_/A vssd1 vssd1 vccd1 vccd1 _13158_/A sky130_fd_sc_hd__o21bai_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11837_ hold200/A _11559_/A _11918_/B _11920_/C1 vssd1 vssd1 vccd1 vccd1 _11837_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11219__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11768_ _11972_/A _11972_/B _11973_/A vssd1 vssd1 vccd1 vccd1 _11768_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_83_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10719_ _10719_/A _10719_/B vssd1 vssd1 vccd1 vccd1 _10720_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06653__B _06653_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11699_ _11698_/B _11699_/B vssd1 vssd1 vccd1 vccd1 _11700_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10456__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12195__A1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07765__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11942__A1 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11942__B2 _12776_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07930_ _07939_/A _07939_/B vssd1 vssd1 vccd1 vccd1 _07941_/A sky130_fd_sc_hd__and2b_1
X_07861_ _08772_/B2 _12752_/A fanout84/X _08772_/A2 vssd1 vssd1 vccd1 vccd1 _07862_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_48_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07792_ _07969_/A _08134_/B fanout51/X _12734_/A vssd1 vssd1 vccd1 vccd1 _07793_/B
+ sky130_fd_sc_hd__o22a_1
X_06812_ _10972_/A _06810_/X _06811_/X vssd1 vssd1 vccd1 vccd1 _06812_/Y sky130_fd_sc_hd__a21oi_1
X_09600_ _09600_/A _09775_/A vssd1 vssd1 vccd1 vccd1 _09606_/A sky130_fd_sc_hd__nand2_1
X_06743_ reg1_val[7] _06986_/A vssd1 vssd1 vccd1 vccd1 _06744_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09531_ _09529_/X _09530_/X _10246_/S vssd1 vssd1 vccd1 vccd1 _09531_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08323__B1 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06674_ reg1_val[18] _07023_/A vssd1 vssd1 vccd1 vccd1 _06674_/Y sky130_fd_sc_hd__nand2_1
X_09462_ _09462_/A _09462_/B vssd1 vssd1 vccd1 vccd1 _09465_/A sky130_fd_sc_hd__nand2_1
X_08413_ _08413_/A _08413_/B vssd1 vssd1 vccd1 vccd1 _08436_/A sky130_fd_sc_hd__xnor2_2
X_09393_ _10246_/S _09392_/X _09211_/B vssd1 vssd1 vccd1 vccd1 _09394_/A sky130_fd_sc_hd__o21ai_1
X_08344_ _08344_/A _08344_/B vssd1 vssd1 vccd1 vccd1 _08367_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_86_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07429__A2 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06563__B _06915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08275_ _08278_/A _08278_/B vssd1 vssd1 vccd1 vccd1 _08275_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_6_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07226_ _07423_/B _07423_/A vssd1 vssd1 vccd1 vccd1 _07226_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_1_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13241_/CLK sky130_fd_sc_hd__clkbuf_8
X_07157_ _07157_/A _07157_/B vssd1 vssd1 vccd1 vccd1 _07157_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_42_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10197__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09366__S _12726_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07088_ _07165_/A _07528_/C reg1_val[29] vssd1 vssd1 vccd1 vccd1 _07090_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout121 _06944_/X vssd1 vssd1 vccd1 vccd1 _10169_/A sky130_fd_sc_hd__clkbuf_16
Xfanout165 _07116_/X vssd1 vssd1 vccd1 vccd1 _08774_/B1 sky130_fd_sc_hd__buf_4
Xfanout154 _11559_/A vssd1 vssd1 vccd1 vccd1 _12187_/A1 sky130_fd_sc_hd__buf_4
Xfanout143 _06985_/X vssd1 vssd1 vccd1 vccd1 _10064_/B2 sky130_fd_sc_hd__buf_6
Xfanout132 _10156_/A1 vssd1 vssd1 vccd1 vccd1 _08776_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout176 _12781_/A2 vssd1 vssd1 vccd1 vccd1 _13020_/B2 sky130_fd_sc_hd__buf_4
Xfanout198 _09199_/X vssd1 vssd1 vccd1 vccd1 _12290_/C1 sky130_fd_sc_hd__buf_4
Xfanout187 _09452_/A vssd1 vssd1 vccd1 vccd1 _08777_/A sky130_fd_sc_hd__buf_8
XANTENNA__08562__B1 _09600_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout61_A _07153_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09729_ _09729_/A _09729_/B vssd1 vssd1 vccd1 vccd1 _09731_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07117__A1 _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12740_ hold56/X _12788_/B vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__or2_1
XANTENNA__10121__B1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07668__A2 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12671_ _12678_/C _12671_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[22] sky130_fd_sc_hd__xnor2_4
XANTENNA__12949__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11622_ _11622_/A _11622_/B vssd1 vssd1 vccd1 vccd1 _11624_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06628__B1 _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10424__A1 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08093__A2 _08420_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10424__B2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11553_ _11179_/B _11552_/X _11551_/X vssd1 vssd1 vccd1 vccd1 _11554_/B sky130_fd_sc_hd__a21o_1
X_11484_ _12119_/B1 _11570_/B hold289/A vssd1 vssd1 vccd1 vccd1 _11484_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10504_ _10504_/A _10504_/B vssd1 vssd1 vccd1 vccd1 _10504_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13223_ _13248_/CLK hold191/X vssd1 vssd1 vccd1 vccd1 hold228/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10435_ _10435_/A _10435_/B _10435_/C vssd1 vssd1 vccd1 vccd1 _10446_/A sky130_fd_sc_hd__and3_1
X_13154_ hold254/X _13153_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13154_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _12215_/A _12105_/B vssd1 vssd1 vccd1 vccd1 _12221_/B sky130_fd_sc_hd__xnor2_2
X_10366_ _10607_/A _10366_/B vssd1 vssd1 vccd1 vccd1 _10523_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13085_ hold295/X _13165_/A2 _13084_/X _12722_/A vssd1 vssd1 vccd1 vccd1 _13086_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ _10297_/A _10297_/B vssd1 vssd1 vccd1 vccd1 _10311_/A sky130_fd_sc_hd__xor2_1
X_12036_ _12036_/A _12036_/B _12036_/C vssd1 vssd1 vccd1 vccd1 _12102_/C sky130_fd_sc_hd__and3_1
XFILLER_0_18_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06564__C1 _06633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09305__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12938_ _12946_/A hold201/X vssd1 vssd1 vccd1 vccd1 hold202/A sky130_fd_sc_hd__and2_1
XANTENNA__08856__B2 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08856__A1 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12869_ hold5/X hold277/X vssd1 vssd1 vccd1 vccd1 _13121_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_56_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08084__A2 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08060_ _08060_/A _08060_/B vssd1 vssd1 vccd1 vccd1 _08069_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_114_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09033__A1 _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07011_ _07595_/B _07011_/B vssd1 vssd1 vccd1 vccd1 _07225_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10179__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10914__A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08962_ _08963_/A _08963_/B vssd1 vssd1 vccd1 vccd1 _08962_/X sky130_fd_sc_hd__or2_1
X_07913_ _08774_/A2 fanout94/X _12752_/A _08774_/B1 vssd1 vssd1 vccd1 vccd1 _07914_/B
+ sky130_fd_sc_hd__o22a_1
X_08893_ _08894_/A _08894_/B vssd1 vssd1 vccd1 vccd1 _08949_/B sky130_fd_sc_hd__nand2b_1
XANTENNA_fanout196_A _13151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07844_ _07844_/A _07844_/B _07844_/C vssd1 vssd1 vccd1 vccd1 _07848_/A sky130_fd_sc_hd__and3_1
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07775_ _07775_/A _07775_/B vssd1 vssd1 vccd1 vccd1 _07778_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11183__C _11183_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06726_ reg1_val[10] _07319_/A vssd1 vssd1 vccd1 vccd1 _10638_/A sky130_fd_sc_hd__or2_1
XFILLER_0_78_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09514_ _09514_/A _12230_/A vssd1 vssd1 vccd1 vccd1 _09515_/S sky130_fd_sc_hd__nand2_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06657_ reg2_val[21] _06752_/A _06688_/B1 _06656_/Y vssd1 vssd1 vccd1 vccd1 _07052_/B
+ sky130_fd_sc_hd__o2bb2a_2
X_09445_ _10452_/B2 _10557_/A fanout62/X _10527_/A vssd1 vssd1 vccd1 vccd1 _09446_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10654__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10654__B2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06588_ reg2_val[28] _06752_/A _06688_/B1 _06587_/Y vssd1 vssd1 vccd1 vccd1 _12250_/A
+ sky130_fd_sc_hd__o2bb2a_4
X_09376_ _12361_/B _09370_/X _09375_/X _09851_/B vssd1 vssd1 vccd1 vccd1 _09376_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10406__A1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08075__A2 _07168_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08327_ _08359_/A _08359_/B vssd1 vssd1 vccd1 vccd1 _08360_/A sky130_fd_sc_hd__or2_2
XANTENNA__07389__B _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10406__B2 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08258_ _08259_/A _08259_/B vssd1 vssd1 vccd1 vccd1 _08258_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_117_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09885__A _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07209_ _07209_/A _07209_/B vssd1 vssd1 vccd1 vccd1 _07223_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08189_ _08773_/A _08189_/B vssd1 vssd1 vccd1 vccd1 _08190_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10220_ _10220_/A _10220_/B vssd1 vssd1 vccd1 vccd1 _10223_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09109__B _09199_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10151_ _10050_/A _10050_/B _10048_/X vssd1 vssd1 vccd1 vccd1 _10160_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ _09936_/A _09936_/B _09934_/Y vssd1 vssd1 vccd1 vccd1 _10084_/B sky130_fd_sc_hd__a21boi_2
XANTENNA__11655__A _11746_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08535__A0 _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11134__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07889__A2 _08854_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07852__B _07852_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10984_ _12187_/A1 _11201_/C hold215/A vssd1 vssd1 vccd1 vccd1 _10984_/Y sky130_fd_sc_hd__a21oi_1
X_12723_ _12723_/A _12723_/B vssd1 vssd1 vccd1 vccd1 _12723_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_85_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10645__B2 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12654_ reg1_val[19] _12714_/A vssd1 vssd1 vccd1 vccd1 _12657_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12585_ _12585_/A _12585_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[5] sky130_fd_sc_hd__xor2_4
X_11605_ _11606_/B _11605_/B vssd1 vssd1 vccd1 vccd1 _11709_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_108_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11536_ _11536_/A _11536_/B vssd1 vssd1 vccd1 vccd1 _11539_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13206_ _13303_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
X_11467_ _11379_/B _11379_/C _12131_/A vssd1 vssd1 vccd1 vccd1 _11468_/B sky130_fd_sc_hd__a21o_1
XANTENNA__06931__B _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11398_ hold260/A _11398_/B _11483_/B vssd1 vssd1 vccd1 vccd1 _11400_/B sky130_fd_sc_hd__and3_1
XANTENNA__09566__A2 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10418_ _10418_/A _10418_/B vssd1 vssd1 vccd1 vccd1 _10420_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_110_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13137_ hold262/X _13165_/A2 _13136_/X _13146_/B2 vssd1 vssd1 vccd1 vccd1 hold263/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__08774__B1 _08774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10349_ _10349_/A _10349_/B vssd1 vssd1 vccd1 vccd1 _10351_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ _13068_/A _13068_/B vssd1 vssd1 vccd1 vccd1 _13068_/Y sky130_fd_sc_hd__xnor2_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12019_ _12019_/A _12019_/B vssd1 vssd1 vccd1 vccd1 _12020_/B sky130_fd_sc_hd__and2_1
XFILLER_0_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12086__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07560_ _07559_/B _07559_/C _10555_/A vssd1 vssd1 vccd1 vccd1 _07562_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09230_ _10144_/B2 fanout30/X _10433_/A _08680_/B vssd1 vssd1 vccd1 vccd1 _09231_/B
+ sky130_fd_sc_hd__o22a_1
X_07491_ _07589_/A _07589_/B vssd1 vssd1 vccd1 vccd1 _07590_/A sky130_fd_sc_hd__and2_1
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13050__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09161_ _09153_/X _09160_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09161_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08112_ _08112_/A _08112_/B vssd1 vssd1 vccd1 vccd1 _08121_/B sky130_fd_sc_hd__xnor2_2
X_09092_ _09092_/A _09092_/B vssd1 vssd1 vccd1 vccd1 _09092_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08043_ _08043_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08107_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout209_A _06918_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout111_A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07568__A1 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09994_ _09837_/A _09978_/X _09980_/Y _09981_/X _09993_/X vssd1 vssd1 vccd1 vccd1
+ _09994_/X sky130_fd_sc_hd__a221o_1
XANTENNA__07568__B2 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07953__A _10578_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08945_ _08945_/A _08945_/B vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__nand2_2
XANTENNA__08517__B1 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08876_ _08876_/A _08876_/B vssd1 vssd1 vccd1 vccd1 _08878_/B sky130_fd_sc_hd__xnor2_2
X_07827_ _08443_/A _07827_/B vssd1 vssd1 vccd1 vccd1 _07829_/B sky130_fd_sc_hd__xor2_2
X_07758_ _08853_/A _07758_/B vssd1 vssd1 vccd1 vccd1 _07783_/A sky130_fd_sc_hd__xor2_2
X_06709_ reg1_val[13] _07197_/A vssd1 vssd1 vccd1 vccd1 _06710_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_94_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11922__B wire201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07689_ _08940_/A _07688_/B _07688_/A vssd1 vssd1 vccd1 vccd1 _08969_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_39_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10819__A _10819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09428_ _09428_/A _09428_/B vssd1 vssd1 vccd1 vccd1 _09432_/A sky130_fd_sc_hd__xor2_1
XANTENNA_fanout24_A _07132_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09359_ _09155_/X _09157_/X _09359_/S vssd1 vssd1 vccd1 vccd1 _09359_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13041__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08493__A_N _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12370_ reg1_val[31] _12370_/B vssd1 vssd1 vccd1 vccd1 _12370_/X sky130_fd_sc_hd__or2_1
X_11321_ _11429_/A _11321_/B vssd1 vssd1 vccd1 vccd1 _11325_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11252_ _11253_/B _11252_/B vssd1 vssd1 vccd1 vccd1 _11356_/B sky130_fd_sc_hd__and2b_1
X_11183_ _11379_/A _11183_/B _11183_/C vssd1 vssd1 vccd1 vccd1 _11183_/X sky130_fd_sc_hd__or3_1
XANTENNA__08756__B1 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ _11695_/A _10203_/B vssd1 vssd1 vccd1 vccd1 _10204_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08220__A2 _08672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10134_ _09837_/Y _10118_/Y _10120_/Y _10121_/X _10133_/Y vssd1 vssd1 vccd1 vccd1
+ _10134_/X sky130_fd_sc_hd__o221a_1
X_10065_ _10551_/B _10065_/B vssd1 vssd1 vccd1 vccd1 _10069_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09181__B1 _11197_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09720__A2 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07731__B2 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__A1 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12068__B1 _12345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10967_ _10890_/X _11215_/B _10966_/Y vssd1 vssd1 vccd1 vccd1 _10967_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12706_ _12706_/A _12706_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[29] sky130_fd_sc_hd__xnor2_4
X_10898_ _10898_/A _10898_/B vssd1 vssd1 vccd1 vccd1 _10910_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_128_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12637_ reg1_val[15] _12637_/B vssd1 vssd1 vccd1 vccd1 _12639_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13032__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12568_ reg1_val[2] _12568_/B vssd1 vssd1 vccd1 vccd1 _12569_/B sky130_fd_sc_hd__nand2_1
X_12499_ _12516_/A _12499_/B vssd1 vssd1 vccd1 vccd1 _12515_/A sky130_fd_sc_hd__nand2_1
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
X_11519_ fanout32/X _12150_/A _12150_/B fanout29/X vssd1 vssd1 vccd1 vccd1 _11520_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_123_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold229 hold229/A vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 hold218/A vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10554__B1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07970__A1 _07308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06773__A2 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08588__B _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06991_ _10555_/A _06991_/B vssd1 vssd1 vccd1 vccd1 _06993_/B sky130_fd_sc_hd__xnor2_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08730_ _09580_/A _08730_/B vssd1 vssd1 vccd1 vccd1 _08731_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08661_ _08819_/B2 _07322_/A _07322_/B fanout47/X _06952_/Y vssd1 vssd1 vccd1 vccd1
+ _08662_/B sky130_fd_sc_hd__o32a_1
X_07612_ _07612_/A _07612_/B vssd1 vssd1 vccd1 vccd1 _07615_/A sky130_fd_sc_hd__xnor2_4
X_08592_ _08592_/A _08598_/S vssd1 vssd1 vccd1 vccd1 _08595_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_76_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06836__B _12250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07543_ _09772_/A fanout36/X _12736_/A _08821_/B vssd1 vssd1 vccd1 vccd1 _07544_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout159_A _08681_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ _10301_/A _07474_/B vssd1 vssd1 vccd1 vccd1 _07475_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09213_ _11089_/A _09213_/B vssd1 vssd1 vccd1 vccd1 _11195_/C sky130_fd_sc_hd__or2_2
XFILLER_0_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09144_ _09140_/X _09143_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09144_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07238__B1 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12231__B1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12573__B _12573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09075_ _11820_/B _11820_/C vssd1 vssd1 vccd1 vccd1 _09075_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08450__A2 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08026_ _09621_/A _08026_/B vssd1 vssd1 vccd1 vccd1 _08071_/A sky130_fd_sc_hd__xnor2_2
Xfanout1 hold243/A vssd1 vssd1 vccd1 vccd1 fanout1/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07961__A1 _07034_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ _09517_/Y _10979_/B _11089_/A vssd1 vssd1 vccd1 vccd1 _09977_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07961__B2 _09925_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ _08929_/A _08929_/B vssd1 vssd1 vccd1 vccd1 _08928_/X sky130_fd_sc_hd__and2_1
XFILLER_0_99_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08859_ _08859_/A _08859_/B vssd1 vssd1 vccd1 vccd1 _08860_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12748__B _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11870_ _12206_/A _11870_/B vssd1 vssd1 vccd1 vccd1 _11872_/B sky130_fd_sc_hd__xnor2_1
X_10821_ _08733_/A _07174_/B _07435_/Y _10820_/Y vssd1 vssd1 vccd1 vccd1 _10925_/B
+ sky130_fd_sc_hd__a31o_2
XANTENNA__09466__A1 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09466__B2 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10752_ _09828_/Y _10751_/Y _10752_/S vssd1 vssd1 vccd1 vccd1 _10752_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13014__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12422_ _12422_/A _12422_/B _12422_/C vssd1 vssd1 vccd1 vccd1 _12423_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_82_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10683_ _10683_/A _10683_/B _10683_/C vssd1 vssd1 vccd1 vccd1 _10686_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07858__A _09580_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11576__A2 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12353_ _12353_/A _12353_/B vssd1 vssd1 vccd1 vccd1 _12353_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_105_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11304_ hold207/A _12332_/B _11480_/C _11920_/C1 vssd1 vssd1 vccd1 vccd1 _11304_/X
+ sky130_fd_sc_hd__a31o_1
X_12284_ _12284_/A _12284_/B vssd1 vssd1 vccd1 vccd1 _12284_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__10784__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08729__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11235_ _11234_/B _11235_/B vssd1 vssd1 vccd1 vccd1 _11236_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10536__B1 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10000__A2 _09996_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ _11166_/A _11166_/B vssd1 vssd1 vccd1 vccd1 _11169_/A sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_14_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13289_/CLK sky130_fd_sc_hd__clkbuf_8
X_11097_ hold282/A _11096_/X _09200_/X vssd1 vssd1 vccd1 vccd1 _11097_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__07952__A1 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07952__B2 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10117_ _11194_/S _10114_/X _10113_/X _10251_/S vssd1 vssd1 vccd1 vccd1 _10117_/X
+ sky130_fd_sc_hd__a211o_1
X_10048_ _10049_/A _10049_/B vssd1 vssd1 vccd1 vccd1 _10048_/X sky130_fd_sc_hd__or2_1
XFILLER_0_26_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06656__B _12588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11999_ _09183_/Y _10245_/X _10251_/X _09173_/S _11998_/Y vssd1 vssd1 vccd1 vccd1
+ _12000_/A sky130_fd_sc_hd__a221o_1
XFILLER_0_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07468__B1 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07190_ _08733_/A _07194_/C vssd1 vssd1 vccd1 vccd1 _08672_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_14_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_453 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10775__B1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09900_ _09900_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _09900_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09831_ _09144_/X _09168_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09831_/X sky130_fd_sc_hd__mux2_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06974_ _07015_/B _06975_/B vssd1 vssd1 vccd1 vccd1 _06974_/X sky130_fd_sc_hd__xor2_1
XANTENNA__06746__A2 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09762_ _07058_/A _12784_/A fanout18/X _08532_/B vssd1 vssd1 vccd1 vccd1 _09763_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _08713_/A _08713_/B vssd1 vssd1 vccd1 vccd1 _08715_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07008__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09693_ _09544_/A _09544_/B _06777_/B vssd1 vssd1 vccd1 vccd1 _09694_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08644_ _09068_/A _08636_/X _08642_/X _08643_/X _08065_/Y vssd1 vssd1 vccd1 vccd1
+ _09077_/A sky130_fd_sc_hd__a311oi_4
XFILLER_0_83_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08575_ _08577_/A _08577_/C vssd1 vssd1 vccd1 vccd1 _08602_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12568__B _12568_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06566__B _06567_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07526_ _07526_/A _07526_/B vssd1 vssd1 vccd1 vccd1 _07527_/B sky130_fd_sc_hd__xnor2_1
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07457_ _07458_/A _07458_/B vssd1 vssd1 vccd1 vccd1 _07459_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_106_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07388_ _07388_/A _07388_/B vssd1 vssd1 vccd1 vccd1 _07414_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12755__A1 _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09127_ reg1_val[7] reg1_val[24] _09172_/S vssd1 vssd1 vccd1 vccd1 _09127_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09058_ _09058_/A _09058_/B vssd1 vssd1 vccd1 vccd1 _09059_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08009_ _08009_/A _08009_/B vssd1 vssd1 vccd1 vccd1 _08011_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_4_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout91_A _07197_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13180__B2 _06537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ _11499_/A _11020_/B vssd1 vssd1 vccd1 vccd1 _11024_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09923__A2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10551__B _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12971_ hold121/X _12723_/A _13170_/B _13256_/Q _13066_/A vssd1 vssd1 vccd1 vccd1
+ hold122/A sky130_fd_sc_hd__o221a_1
XFILLER_0_99_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11922_ _11922_/A wire201/X vssd1 vssd1 vccd1 vccd1 _11922_/Y sky130_fd_sc_hd__nand2_1
X_11853_ _11853_/A _11853_/B vssd1 vssd1 vccd1 vccd1 _11854_/B sky130_fd_sc_hd__and2_1
XFILLER_0_95_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10804_ _12019_/A _10804_/B vssd1 vssd1 vccd1 vccd1 _10805_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12994__A1 _11429_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11784_ _11783_/B _11783_/C _11783_/A vssd1 vssd1 vccd1 vccd1 _11785_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_103_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10735_ _10734_/B _10734_/C _10959_/A vssd1 vssd1 vccd1 vccd1 _10736_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07870__B1 _08695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10666_ _12022_/A _10666_/B vssd1 vssd1 vccd1 vccd1 _10670_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12405_ _12578_/B _12405_/B vssd1 vssd1 vccd1 vccd1 _12406_/B sky130_fd_sc_hd__or2_1
XFILLER_0_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08414__A2 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10597_ _10476_/A _10476_/B _10474_/Y vssd1 vssd1 vccd1 vccd1 _10599_/B sky130_fd_sc_hd__a21oi_4
X_12336_ _12373_/A1 _09370_/X _09396_/X _09183_/Y _12335_/Y vssd1 vssd1 vccd1 vccd1
+ _12336_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12267_ _12159_/A _12214_/A _12214_/B vssd1 vssd1 vccd1 vccd1 _12267_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_120_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11218_ _11129_/A _11129_/B _11126_/A vssd1 vssd1 vccd1 vccd1 _11221_/A sky130_fd_sc_hd__a21o_1
X_12198_ _12145_/Y _12148_/B _12144_/A vssd1 vssd1 vccd1 vccd1 _12202_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__07925__A1 _08748_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07925__B2 _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11182__B1 _11183_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11149_ _11150_/A _11150_/B vssd1 vssd1 vccd1 vccd1 _11151_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_128_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06690_ reg1_val[16] _07168_/A vssd1 vssd1 vccd1 vccd1 _06693_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_77_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07262__S _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08360_ _08360_/A _08360_/B vssd1 vssd1 vccd1 vccd1 _08363_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11237__A1 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07311_ _07319_/A _06946_/X _07319_/B _06807_/B vssd1 vssd1 vccd1 vccd1 _07313_/B
+ sky130_fd_sc_hd__a211o_2
XANTENNA__11237__B2 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08291_ _08299_/B _08299_/A vssd1 vssd1 vccd1 vccd1 _08291_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_73_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10996__B1 _12345_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11788__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07861__B1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07242_ _09467_/A _07242_/B vssd1 vssd1 vccd1 vccd1 _07249_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_6_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07498__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07173_ _07180_/B _07174_/B vssd1 vssd1 vccd1 vccd1 _07173_/Y sky130_fd_sc_hd__nor2_4
XFILLER_0_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09602__A1 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09602__B2 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06967__A2 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout303 _11823_/S vssd1 vssd1 vccd1 vccd1 _09968_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09814_ _09814_/A _09814_/B vssd1 vssd1 vccd1 vccd1 _10229_/B sky130_fd_sc_hd__xnor2_4
X_06957_ _11780_/A _06965_/C vssd1 vssd1 vccd1 vccd1 _06960_/A sky130_fd_sc_hd__and2_1
X_09745_ _09746_/A _09746_/B vssd1 vssd1 vccd1 vccd1 _09881_/A sky130_fd_sc_hd__nor2_1
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06888_ instruction[6] instruction[5] instruction[4] vssd1 vssd1 vccd1 vccd1 _06888_/Y
+ sky130_fd_sc_hd__a21oi_1
X_09676_ _09357_/X _09359_/X _09676_/S vssd1 vssd1 vccd1 vccd1 _09676_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10279__A2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _09061_/A _09061_/B _09070_/B _08624_/Y vssd1 vssd1 vccd1 vccd1 _09064_/B
+ sky130_fd_sc_hd__a31o_2
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ _09898_/A _08558_/B vssd1 vssd1 vccd1 vccd1 _08559_/C sky130_fd_sc_hd__xor2_1
XANTENNA__12976__A1 _08777_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08489_ _08489_/A _08489_/B vssd1 vssd1 vccd1 vccd1 _08491_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11779__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07509_ _11134_/B2 fanout52/X _10677_/B fanout57/X vssd1 vssd1 vccd1 vccd1 _07510_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_119_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10520_ _09205_/B _10508_/X _10519_/X _10499_/X vssd1 vssd1 vccd1 vccd1 _10520_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10451_ _10337_/A _10337_/B _10334_/A vssd1 vssd1 vccd1 vccd1 _10463_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13170_ hold137/X _13170_/B vssd1 vssd1 vccd1 vccd1 hold138/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10382_ _09201_/X _10380_/Y _10381_/X _12243_/B1 _06739_/B vssd1 vssd1 vccd1 vccd1
+ _10383_/A sky130_fd_sc_hd__o32a_1
XFILLER_0_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07855__B _07855_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12121_ hold264/A _12119_/X _12120_/Y vssd1 vssd1 vccd1 vccd1 _12121_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12052_ _12050_/Y _12052_/B vssd1 vssd1 vccd1 vccd1 _12053_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10281__B _10551_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ _11003_/A _11003_/B vssd1 vssd1 vccd1 vccd1 _11005_/C sky130_fd_sc_hd__nor2_1
XANTENNA__08580__A1 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10911__B1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07871__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08580__B2 _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13084__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ _13169_/A hold232/X vssd1 vssd1 vccd1 vccd1 hold233/A sky130_fd_sc_hd__and2_1
X_11905_ _11738_/S _11904_/X _11903_/X vssd1 vssd1 vccd1 vccd1 _11906_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_59_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12885_ _12885_/A _12885_/B vssd1 vssd1 vccd1 vccd1 _13153_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11219__A1 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _11559_/A _11918_/B hold200/A vssd1 vssd1 vccd1 vccd1 _11836_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11219__B2 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11767_ _11730_/D _11767_/B vssd1 vssd1 vccd1 vccd1 _11972_/B sky130_fd_sc_hd__and2b_1
X_10718_ _10718_/A _10718_/B vssd1 vssd1 vccd1 vccd1 _10719_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_83_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11698_ _11699_/B _11698_/B vssd1 vssd1 vccd1 vccd1 _11791_/B sky130_fd_sc_hd__and2b_1
X_10649_ _10400_/S _10645_/X _10648_/X vssd1 vssd1 vccd1 vccd1 dest_val[10] sky130_fd_sc_hd__o21ai_4
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12319_ _12319_/A _12319_/B vssd1 vssd1 vccd1 vccd1 _12319_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11942__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13299_ _13309_/CLK _13299_/D vssd1 vssd1 vccd1 vccd1 hold289/A sky130_fd_sc_hd__dfxtp_1
X_07860_ _07880_/A _07880_/B vssd1 vssd1 vccd1 vccd1 _07860_/Y sky130_fd_sc_hd__nor2_1
X_07791_ _07790_/A _07790_/B _07790_/C vssd1 vssd1 vccd1 vccd1 _07802_/B sky130_fd_sc_hd__o21ai_1
X_06811_ _07197_/A reg1_val[13] vssd1 vssd1 vccd1 vccd1 _06811_/X sky130_fd_sc_hd__and2b_1
X_06742_ reg1_val[7] _06986_/A vssd1 vssd1 vccd1 vccd1 _06742_/Y sky130_fd_sc_hd__nor2_1
X_09530_ _09149_/X _09174_/X _09679_/S vssd1 vssd1 vccd1 vccd1 _09530_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08323__A1 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08323__B2 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _09461_/A _09461_/B vssd1 vssd1 vccd1 vccd1 _09462_/B sky130_fd_sc_hd__nand2_1
X_06673_ reg1_val[18] _07023_/A vssd1 vssd1 vccd1 vccd1 _06676_/A sky130_fd_sc_hd__and2_1
XFILLER_0_78_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08412_ _08413_/A _08413_/B vssd1 vssd1 vccd1 vccd1 _08412_/X sky130_fd_sc_hd__or2_1
XFILLER_0_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09392_ _09159_/X _09213_/B _09392_/S vssd1 vssd1 vccd1 vccd1 _09392_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07005__B _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__B1 _08672_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08343_ _08343_/A _08343_/B vssd1 vssd1 vccd1 vccd1 _08367_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout239_A _09201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08274_ _09621_/A _08274_/B vssd1 vssd1 vccd1 vccd1 _08278_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10969__B1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09220__B _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07225_ _07225_/A _07225_/B vssd1 vssd1 vccd1 vccd1 _07423_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07156_ _07126_/B _07128_/B _07128_/C _07135_/B vssd1 vssd1 vccd1 vccd1 _07157_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__10197__A1 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07087_ reg1_val[28] _07087_/B _07087_/C _12697_/B vssd1 vssd1 vccd1 vccd1 _07528_/C
+ sky130_fd_sc_hd__or4_2
XANTENNA__10197__B2 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout122 _07324_/Y vssd1 vssd1 vccd1 vccd1 _10433_/A sky130_fd_sc_hd__buf_8
Xfanout111 _11604_/A vssd1 vssd1 vccd1 vccd1 _10565_/A sky130_fd_sc_hd__buf_12
Xfanout100 _09925_/A1 vssd1 vssd1 vccd1 vccd1 _11134_/B2 sky130_fd_sc_hd__buf_8
XFILLER_0_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout155 _11559_/A vssd1 vssd1 vccd1 vccd1 _12332_/B sky130_fd_sc_hd__buf_4
Xfanout144 _10144_/B2 vssd1 vssd1 vccd1 vccd1 _08841_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout133 _07081_/Y vssd1 vssd1 vccd1 vccd1 _10156_/A1 sky130_fd_sc_hd__buf_8
Xfanout177 _12781_/A2 vssd1 vssd1 vccd1 vccd1 _12980_/A2 sky130_fd_sc_hd__clkbuf_4
Xfanout199 _09199_/X vssd1 vssd1 vccd1 vccd1 _11920_/C1 sky130_fd_sc_hd__buf_2
Xfanout188 _07026_/Y vssd1 vssd1 vccd1 vccd1 _09452_/A sky130_fd_sc_hd__clkbuf_16
Xfanout166 _07110_/Y vssd1 vssd1 vccd1 vccd1 _09618_/B2 sky130_fd_sc_hd__buf_4
XANTENNA__08562__B2 _08544_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07989_ _07134_/A fanout62/X _07869_/B _07055_/Y vssd1 vssd1 vccd1 vccd1 _07990_/B
+ sky130_fd_sc_hd__o22a_2
X_09728_ _10301_/A _09728_/B vssd1 vssd1 vccd1 vccd1 _09729_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout54_A fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09659_ _09659_/A _09659_/B vssd1 vssd1 vccd1 vccd1 _10229_/A sky130_fd_sc_hd__xnor2_4
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12662_/Y _12666_/B _12664_/B vssd1 vssd1 vccd1 vccd1 _12671_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__11941__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11621_ _11536_/A _11536_/B _11534_/Y vssd1 vssd1 vccd1 vccd1 _11622_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10557__A _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10424__A2 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11552_ _11552_/A _11552_/B vssd1 vssd1 vccd1 vccd1 _11552_/X sky130_fd_sc_hd__and2_1
X_11483_ hold260/A _11483_/B vssd1 vssd1 vccd1 vccd1 _11570_/B sky130_fd_sc_hd__or2_1
XFILLER_0_107_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12772__A _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10503_ _10501_/Y _10503_/B vssd1 vssd1 vccd1 vccd1 _10504_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_52_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13222_ _13243_/CLK _13222_/D vssd1 vssd1 vccd1 vccd1 hold189/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10434_ _10433_/C _10433_/D _07325_/Y _10551_/B vssd1 vssd1 vccd1 vccd1 _10435_/C
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13079__S fanout1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13153_ _13153_/A _13153_/B vssd1 vssd1 vccd1 vccd1 _13153_/Y sky130_fd_sc_hd__xnor2_1
X_10365_ _09818_/B _10362_/Y _10851_/B vssd1 vssd1 vccd1 vccd1 _10366_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_103_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06800__A1 _06866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _11967_/A _11816_/B _11967_/B _12101_/X _12103_/X vssd1 vssd1 vccd1 vccd1
+ _12105_/B sky130_fd_sc_hd__a41o_1
X_13084_ hold274/X _13083_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13084_/X sky130_fd_sc_hd__mux2_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10297_/A _10297_/B vssd1 vssd1 vccd1 vccd1 _10420_/B sky130_fd_sc_hd__and2_1
XFILLER_0_109_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12035_ _12035_/A vssd1 vssd1 vccd1 vccd1 _12102_/B sky130_fd_sc_hd__inv_2
XANTENNA__09750__B1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_46 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12937_ hold221/A _12947_/A2 _13168_/B1 hold200/X vssd1 vssd1 vccd1 vccd1 hold201/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08856__A2 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12868_ _13117_/A _12867_/B _12804_/X vssd1 vssd1 vccd1 vccd1 _13122_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11851__A _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11819_ _11820_/A _11820_/B _11820_/C vssd1 vssd1 vccd1 vccd1 _11819_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12799_ hold262/X hold17/X vssd1 vssd1 vccd1 vccd1 _13139_/A sky130_fd_sc_hd__nand2b_1
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07816__B1 fanout55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07010_ _07010_/A _07010_/B vssd1 vssd1 vccd1 vccd1 _07011_/B sky130_fd_sc_hd__and2_1
XANTENNA__10179__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10179__B2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_4_14_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08961_ _08930_/A _08930_/B _08928_/X vssd1 vssd1 vccd1 vccd1 _08963_/B sky130_fd_sc_hd__a21oi_4
X_07912_ _09621_/A _07912_/B vssd1 vssd1 vccd1 vccd1 _07919_/A sky130_fd_sc_hd__xnor2_2
X_08892_ _08949_/A _08892_/B vssd1 vssd1 vccd1 vccd1 _08894_/B sky130_fd_sc_hd__and2_1
X_07843_ _07829_/A _07829_/C _07829_/B vssd1 vssd1 vccd1 vccd1 _07844_/C sky130_fd_sc_hd__a21o_1
XANTENNA__09741__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06839__B _07157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07774_ _08415_/A _07774_/B vssd1 vssd1 vccd1 vccd1 _07775_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_79_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06725_ _07319_/A vssd1 vssd1 vccd1 vccd1 _07318_/A sky130_fd_sc_hd__inv_2
X_09513_ _09403_/X _09559_/D _09512_/Y vssd1 vssd1 vccd1 vccd1 _09513_/Y sky130_fd_sc_hd__a21oi_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06656_ _06687_/A _12588_/B vssd1 vssd1 vccd1 vccd1 _06656_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09444_ _09444_/A _09444_/B vssd1 vssd1 vccd1 vccd1 _09485_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10654__A2 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09231__A _10306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06587_ _06687_/A _12626_/B vssd1 vssd1 vccd1 vccd1 _06587_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_93_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09375_ _11197_/S _09375_/B vssd1 vssd1 vccd1 vccd1 _09375_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07807__B1 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08326_ _08777_/A _08326_/B vssd1 vssd1 vccd1 vccd1 _08359_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10406__A2 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08257_ _08259_/A _08259_/B vssd1 vssd1 vccd1 vccd1 _08257_/X sky130_fd_sc_hd__and2_1
XFILLER_0_105_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09885__B _12349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08188_ _08841_/A1 _08772_/A2 _08835_/B1 _08772_/B2 vssd1 vssd1 vccd1 vccd1 _08189_/B
+ sky130_fd_sc_hd__o22a_1
X_07208_ _07209_/B _07209_/A vssd1 vssd1 vccd1 vccd1 _07208_/Y sky130_fd_sc_hd__nand2b_1
X_07139_ _07139_/A _07139_/B vssd1 vssd1 vccd1 vccd1 _09252_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_30_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10150_ _10150_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _10175_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10081_ _09919_/A _09919_/C _09919_/B vssd1 vssd1 vccd1 vccd1 _10084_/A sky130_fd_sc_hd__a21boi_2
XFILLER_0_97_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10983_ hold195/A _10983_/B vssd1 vssd1 vccd1 vccd1 _11201_/C sky130_fd_sc_hd__or2_1
XFILLER_0_69_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12722_ _12722_/A _12722_/B vssd1 vssd1 vccd1 vccd1 _12742_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_85_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12653_ _12650_/B _12652_/B _12648_/X vssd1 vssd1 vccd1 vccd1 _12655_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_108_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11604_ _11604_/A _11604_/B vssd1 vssd1 vccd1 vccd1 _11605_/B sky130_fd_sc_hd__xnor2_1
X_12584_ _12582_/Y _12584_/B vssd1 vssd1 vccd1 vccd1 _12585_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_53_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11535_ _11535_/A _11535_/B vssd1 vssd1 vccd1 vccd1 _11536_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13205_ _13303_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xmax_cap119 _12143_/A vssd1 vssd1 vccd1 vccd1 _10301_/A sky130_fd_sc_hd__clkbuf_8
X_11466_ _11406_/X _11586_/A _11465_/Y vssd1 vssd1 vccd1 vccd1 _11466_/X sky130_fd_sc_hd__a21o_1
X_11397_ hold294/A _11397_/B vssd1 vssd1 vccd1 vccd1 _11483_/B sky130_fd_sc_hd__or2_1
XFILLER_0_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10417_ _10284_/A _10284_/B _10283_/A vssd1 vssd1 vccd1 vccd1 _10418_/B sky130_fd_sc_hd__a21o_1
X_13136_ hold256/X _13135_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13136_/X sky130_fd_sc_hd__mux2_1
XANTENNA__08774__B2 _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08774__A1 _12768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__B1 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _10348_/A _10348_/B vssd1 vssd1 vccd1 vccd1 _10349_/B sky130_fd_sc_hd__xnor2_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13067_/A _13067_/B vssd1 vssd1 vccd1 vccd1 _13068_/B sky130_fd_sc_hd__nand2_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _07389_/B fanout83/X fanout81/X _07099_/X vssd1 vssd1 vccd1 vccd1 _10280_/B
+ sky130_fd_sc_hd__o22a_1
X_12018_ _12019_/A _12019_/B vssd1 vssd1 vccd1 vccd1 _12020_/A sky130_fd_sc_hd__nor2_1
XANTENNA__06659__B _07052_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12086__A1 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12086__B2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07490_ _10565_/A _07490_/B vssd1 vssd1 vccd1 vccd1 _07589_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09160_ _09156_/X _09159_/X _09392_/S vssd1 vssd1 vccd1 vccd1 _09160_/X sky130_fd_sc_hd__mux2_1
X_08111_ _08108_/A _08108_/B _08166_/A vssd1 vssd1 vccd1 vccd1 _08121_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_114_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09091_ _09090_/A _09090_/B _09103_/B vssd1 vssd1 vccd1 vccd1 _09092_/B sky130_fd_sc_hd__a21oi_2
X_08042_ _08853_/A _08042_/B vssd1 vssd1 vccd1 vccd1 _08107_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_44_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout104_A _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09993_ _12361_/B _09851_/B _09992_/Y _09987_/X vssd1 vssd1 vccd1 vccd1 _09993_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__07568__A2 _07389_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08944_ _08944_/A _08944_/B vssd1 vssd1 vccd1 vccd1 _08945_/B sky130_fd_sc_hd__or2_1
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08517__B2 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08517__A1 _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ _08876_/A _08876_/B vssd1 vssd1 vccd1 vccd1 _08886_/A sky130_fd_sc_hd__nand2b_1
X_07826_ _12762_/A _08692_/A2 _08692_/B1 _12760_/A vssd1 vssd1 vccd1 vccd1 _07827_/B
+ sky130_fd_sc_hd__o22a_1
X_07757_ _10281_/A _07182_/X _07325_/Y _07173_/Y vssd1 vssd1 vccd1 vccd1 _07758_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06708_ reg1_val[13] _07197_/A vssd1 vssd1 vccd1 vccd1 _06708_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07688_ _07688_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _08940_/B sky130_fd_sc_hd__and2_1
X_06639_ _11922_/A _06639_/B vssd1 vssd1 vccd1 vccd1 _11906_/A sky130_fd_sc_hd__nor2_1
X_09427_ _09428_/A _09428_/B vssd1 vssd1 vccd1 vccd1 _09596_/A sky130_fd_sc_hd__and2_1
XFILLER_0_19_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09358_ _09356_/X _09357_/X _09676_/S vssd1 vssd1 vccd1 vccd1 _09358_/X sky130_fd_sc_hd__mux2_1
XANTENNA__09896__A _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08309_ _08309_/A _08309_/B _08309_/C vssd1 vssd1 vccd1 vccd1 _08309_/X sky130_fd_sc_hd__and3_1
XANTENNA_fanout17_A _12786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_123 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11320_ _11429_/A _11321_/B vssd1 vssd1 vccd1 vccd1 _11434_/A sky130_fd_sc_hd__nor2_1
X_09289_ _09289_/A _09289_/B vssd1 vssd1 vccd1 vccd1 _09291_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08305__A _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12001__A1 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11251_ _11327_/A _11251_/B vssd1 vssd1 vccd1 vccd1 _11253_/B sky130_fd_sc_hd__nor2_1
X_11182_ _11379_/A _11183_/B _11183_/C vssd1 vssd1 vccd1 vccd1 _11184_/B sky130_fd_sc_hd__o21a_1
XANTENNA__08756__B2 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08756__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ fanout69/X fanout46/X _11603_/A _11431_/A vssd1 vssd1 vccd1 vccd1 _10203_/B
+ sky130_fd_sc_hd__o22a_1
X_10133_ _11831_/S _09851_/B _10132_/Y _10127_/X vssd1 vssd1 vccd1 vccd1 _10133_/Y
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_30_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09705__B1 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ _10144_/B2 _07278_/B fanout7/X _10064_/B2 vssd1 vssd1 vccd1 vccd1 _10065_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07731__A2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10966_ _10890_/X _11215_/B _12223_/B1 vssd1 vssd1 vccd1 vccd1 _10966_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13017__B1 _13151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08692__B1 _08692_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12705_ _12705_/A _12705_/B vssd1 vssd1 vccd1 vccd1 _12706_/B sky130_fd_sc_hd__or2_2
X_10897_ _10898_/B _10898_/A vssd1 vssd1 vccd1 vccd1 _11005_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12636_ _12639_/B _12636_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[14] sky130_fd_sc_hd__and2_4
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12567_ reg1_val[2] _12568_/B vssd1 vssd1 vccd1 vccd1 _12567_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12498_ _12551_/A _12498_/B vssd1 vssd1 vccd1 vccd1 _12499_/B sky130_fd_sc_hd__or2_1
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11518_ _12206_/A _11518_/B vssd1 vssd1 vccd1 vccd1 _11522_/A sky130_fd_sc_hd__xnor2_1
Xhold219 hold219/A vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11449_ _11449_/A _11449_/B vssd1 vssd1 vccd1 vccd1 _11451_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13119_ hold277/X _13165_/A2 _13118_/X _13146_/B2 vssd1 vssd1 vccd1 vccd1 hold278/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10554__A1 _06989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _10144_/B2 _08681_/A _10064_/B2 fanout33/X vssd1 vssd1 vccd1 vccd1 _06991_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07970__A2 _07308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06773__A3 _12573_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08660_ _08836_/A _08660_/B vssd1 vssd1 vccd1 vccd1 _08664_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07183__B1 _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ _07611_/A _07611_/B vssd1 vssd1 vccd1 vccd1 _07612_/B sky130_fd_sc_hd__xor2_4
XANTENNA__06930__B1 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08591_ _08592_/A _08591_/B vssd1 vssd1 vccd1 vccd1 _08591_/X sky130_fd_sc_hd__and2_1
XFILLER_0_88_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07542_ _07542_/A _07542_/B vssd1 vssd1 vccd1 vccd1 _07579_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12200__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07473_ _08821_/B _09888_/B2 _12736_/A fanout36/X vssd1 vssd1 vccd1 vccd1 _07474_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09212_ _11089_/A _09213_/B vssd1 vssd1 vccd1 vccd1 _09212_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_57_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09143_ _09141_/X _09142_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09143_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07238__A1 _12782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10242__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout221_A _07279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07238__B2 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10655__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09074_ _09074_/A _09074_/B vssd1 vssd1 vccd1 vccd1 _11820_/C sky130_fd_sc_hd__xnor2_4
XANTENNA__08125__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10255__A2_N _06928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08025_ _07134_/A _12760_/A _07869_/B _09925_/A1 vssd1 vssd1 vccd1 vccd1 _08026_/B
+ sky130_fd_sc_hd__o22a_1
Xfanout2 hold243/A vssd1 vssd1 vccd1 vccd1 fanout2/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_4_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09976_ _09358_/X _09367_/X _10249_/S vssd1 vssd1 vccd1 vccd1 _10979_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07961__A2 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08927_ _08927_/A _08927_/B vssd1 vssd1 vccd1 vccd1 _08929_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12298__A1 _07243_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08858_ _08859_/A _08859_/B vssd1 vssd1 vccd1 vccd1 _08860_/A sky130_fd_sc_hd__or2_1
X_07809_ _07809_/A _07809_/B vssd1 vssd1 vccd1 vccd1 _07812_/B sky130_fd_sc_hd__xor2_1
XANTENNA__11933__B _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06921__B1 _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08789_ _08700_/A _08700_/B _08698_/X vssd1 vssd1 vccd1 vccd1 _08791_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10820_ _07180_/B _07435_/Y _08733_/A vssd1 vssd1 vccd1 vccd1 _10820_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__09466__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10751_ _10751_/A vssd1 vssd1 vccd1 vccd1 _10751_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07204__A _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12421_ _12422_/A _12422_/B _12422_/C vssd1 vssd1 vccd1 vccd1 _12429_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10682_ _10683_/A _10683_/B _10683_/C vssd1 vssd1 vccd1 vccd1 _10686_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06762__B _07001_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10565__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12352_ _12352_/A _12352_/B vssd1 vssd1 vccd1 vccd1 _12353_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10784__A1 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11303_ _12332_/B _11480_/C hold207/A vssd1 vssd1 vccd1 vccd1 _11303_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11981__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12283_ _12361_/C _12282_/Y _12361_/B vssd1 vssd1 vccd1 vccd1 _12283_/X sky130_fd_sc_hd__o21a_1
XANTENNA__10784__B2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__A _08443_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08729__A1 _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08729__B2 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ _11235_/B _11234_/B vssd1 vssd1 vccd1 vccd1 _11354_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_120_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10536__B2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10536__A1 fanout32/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11165_ _11166_/A _11166_/B vssd1 vssd1 vccd1 vccd1 _11274_/A sky130_fd_sc_hd__and2_1
X_11096_ hold295/A _11198_/C _09842_/B vssd1 vssd1 vccd1 vccd1 _11096_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07952__A2 _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ _09394_/Y _11089_/B _11089_/A vssd1 vssd1 vccd1 vccd1 _10116_/X sky130_fd_sc_hd__mux2_1
X_10047_ _11125_/A _10047_/B vssd1 vssd1 vccd1 vccd1 _10049_/B sky130_fd_sc_hd__xnor2_1
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13116__A _13116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11998_ _06602_/Y _12243_/B1 _11996_/Y _06603_/X _11997_/X vssd1 vssd1 vccd1 vccd1
+ _11998_/Y sky130_fd_sc_hd__o221ai_4
XFILLER_0_128_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08665__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07114__A _07126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07468__B2 _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07468__A1 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10949_ _10949_/A _10949_/B vssd1 vssd1 vccd1 vccd1 _10951_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12619_ reg1_val[12] _12620_/B vssd1 vssd1 vccd1 vccd1 _12629_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09830_ _09129_/X _09137_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09830_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _07175_/A _07175_/B _07303_/B vssd1 vssd1 vccd1 vccd1 _06975_/B sky130_fd_sc_hd__o21ai_4
XANTENNA__06746__A3 _12593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09761_ _09761_/A _09761_/B vssd1 vssd1 vccd1 vccd1 _09770_/A sky130_fd_sc_hd__xor2_2
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _08712_/A _08712_/B vssd1 vssd1 vccd1 vccd1 _08713_/B sky130_fd_sc_hd__xor2_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09692_ _11195_/A _09691_/X _09214_/A vssd1 vssd1 vccd1 vccd1 _12235_/B sky130_fd_sc_hd__o21a_1
X_08643_ _08643_/A _08643_/B _09076_/A _09074_/B vssd1 vssd1 vccd1 vccd1 _08643_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA_fanout171_A _07047_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08574_ _08568_/B _08567_/C _08567_/B vssd1 vssd1 vccd1 vccd1 _08577_/C sky130_fd_sc_hd__o21ai_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07525_ _07525_/A _07525_/B vssd1 vssd1 vccd1 vccd1 _07526_/B sky130_fd_sc_hd__xor2_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06863__A _09180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07456_ _10658_/A _07456_/B vssd1 vssd1 vccd1 vccd1 _07458_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08408__B1 _09618_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ _07387_/A _07387_/B vssd1 vssd1 vccd1 vccd1 _07388_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12755__A2 _12781_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09126_ reg1_val[6] reg1_val[25] _09172_/S vssd1 vssd1 vccd1 vccd1 _09126_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09057_ _09057_/A _09057_/B vssd1 vssd1 vccd1 vccd1 _09059_/B sky130_fd_sc_hd__xnor2_2
X_08008_ _08008_/A _08008_/B vssd1 vssd1 vccd1 vccd1 _08009_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_4_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13180__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout84_A _07305_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _09657_/X _09812_/X _09813_/X vssd1 vssd1 vccd1 vccd1 _09959_/Y sky130_fd_sc_hd__a21oi_1
X_12970_ _07046_/B _12788_/B hold153/X vssd1 vssd1 vccd1 vccd1 _13255_/D sky130_fd_sc_hd__a21boi_1
XANTENNA__12140__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11921_ _11922_/A _09383_/B _09191_/X vssd1 vssd1 vccd1 vccd1 _11921_/X sky130_fd_sc_hd__o21a_1
X_11852_ _11853_/A _11853_/B vssd1 vssd1 vccd1 vccd1 _11938_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08647__B1 _07179_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10803_ fanout32/X _11688_/A fanout70/X fanout29/X vssd1 vssd1 vccd1 vccd1 _10804_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_28_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07869__A _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11783_ _11783_/A _11783_/B _11783_/C vssd1 vssd1 vccd1 vccd1 _11861_/A sky130_fd_sc_hd__nor3_2
XANTENNA__12994__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10734_ _10959_/A _10734_/B _10734_/C vssd1 vssd1 vccd1 vccd1 _10736_/A sky130_fd_sc_hd__and3_1
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10665_ fanout37/X _11347_/A _11134_/B2 fanout35/X vssd1 vssd1 vccd1 vccd1 _10666_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_106_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12404_ _12578_/B _12405_/B vssd1 vssd1 vccd1 vccd1 _12415_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_51_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12335_ _06631_/B _12333_/X _12334_/X vssd1 vssd1 vccd1 vccd1 _12335_/Y sky130_fd_sc_hd__o21ai_1
X_10596_ _10596_/A _10596_/B vssd1 vssd1 vccd1 vccd1 _10599_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12266_ _12266_/A _12266_/B vssd1 vssd1 vccd1 vccd1 _12312_/B sky130_fd_sc_hd__or2_1
XFILLER_0_10_118 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13171__A2 _06537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12197_ _12152_/A _12152_/B _12151_/C vssd1 vssd1 vccd1 vccd1 _12209_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__09308__B _09309_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11217_ _11217_/A _11217_/B vssd1 vssd1 vccd1 vccd1 _11272_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07925__A2 _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11182__A1 _11379_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11148_ _11148_/A _11148_/B vssd1 vssd1 vccd1 vccd1 _11150_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11079_ _09059_/C _11077_/X _11078_/Y vssd1 vssd1 vccd1 vccd1 _11079_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__06948__A _06964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11237__A2 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07310_ _07318_/A _07050_/A _07075_/B _07018_/A vssd1 vssd1 vccd1 vccd1 _07313_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08290_ _08290_/A _08290_/B vssd1 vssd1 vccd1 vccd1 _08299_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07861__B2 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07861__A1 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07241_ _09618_/B2 _10677_/A fanout58/X _09618_/A1 vssd1 vssd1 vccd1 vccd1 _07242_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__12737__A2 _12788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07172_ _08855_/A _07172_/B vssd1 vssd1 vccd1 vccd1 _07174_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09602__A2 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout304 instruction[7] vssd1 vssd1 vccd1 vccd1 _11823_/S sky130_fd_sc_hd__buf_6
XANTENNA__07916__A2 _07168_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07019__A _07178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09813_ _09814_/A _09814_/B vssd1 vssd1 vccd1 vccd1 _09813_/X sky130_fd_sc_hd__and2_1
X_06956_ _06956_/A _06956_/B vssd1 vssd1 vccd1 vccd1 _06965_/C sky130_fd_sc_hd__xnor2_4
X_09744_ _10458_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _09746_/B sky130_fd_sc_hd__xnor2_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09675_ _09671_/X _09674_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _09675_/X sky130_fd_sc_hd__mux2_1
X_06887_ _09200_/A instruction[5] vssd1 vssd1 vccd1 vccd1 _09202_/B sky130_fd_sc_hd__nand2_2
XANTENNA__09234__A _10301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _08295_/X _08626_/B vssd1 vssd1 vccd1 vccd1 _09063_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__10684__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08557_ _08825_/A2 _09618_/B2 _09618_/A1 _08588_/A vssd1 vssd1 vccd1 vccd1 _08558_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08488_ _08488_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08491_/A sky130_fd_sc_hd__or2_1
X_07508_ _10894_/A _07508_/B vssd1 vssd1 vccd1 vccd1 _07512_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07439_ _07440_/A _07440_/B vssd1 vssd1 vccd1 vccd1 _07439_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_107_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11430__A2_N fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10450_ _10592_/A _10448_/C _10448_/A vssd1 vssd1 vccd1 vccd1 _10464_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09109_ _09188_/C _09199_/B vssd1 vssd1 vccd1 vccd1 _09109_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10381_ hold268/A _10381_/B vssd1 vssd1 vccd1 vccd1 _10381_/X sky130_fd_sc_hd__and2_1
XFILLER_0_103_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12120_ hold264/A _12119_/X _09200_/X vssd1 vssd1 vccd1 vccd1 _12120_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12051_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _12052_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07368__B1 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11002_ _10920_/A _10920_/B _10917_/A vssd1 vssd1 vccd1 vccd1 _11007_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10911__B2 _10553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10911__A1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08580__A2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11467__A2 _11379_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ _13246_/Q _12955_/A2 _13168_/B1 hold231/X vssd1 vssd1 vccd1 vccd1 hold232/A
+ sky130_fd_sc_hd__a22o_1
X_11904_ _11824_/A _11821_/X _06647_/A vssd1 vssd1 vccd1 vccd1 _11904_/X sky130_fd_sc_hd__a21o_1
X_12884_ hold254/X hold7/X vssd1 vssd1 vccd1 vccd1 _12885_/B sky130_fd_sc_hd__and2b_1
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11835_ hold221/A _11835_/B vssd1 vssd1 vccd1 vccd1 _11918_/B sky130_fd_sc_hd__or2_1
XFILLER_0_83_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11219__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11766_ _10400_/S _11762_/X _11765_/X vssd1 vssd1 vccd1 vccd1 dest_val[21] sky130_fd_sc_hd__o21ai_4
XFILLER_0_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10717_ _10718_/A _10718_/B vssd1 vssd1 vccd1 vccd1 _10717_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_126_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11697_ _11853_/A _11697_/B vssd1 vssd1 vccd1 vccd1 _11698_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11927__B1 _12382_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10648_ _12005_/A _10887_/C _10648_/C vssd1 vssd1 vccd1 vccd1 _10648_/X sky130_fd_sc_hd__or3_1
XFILLER_0_2_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10579_ _10580_/A _10580_/B vssd1 vssd1 vccd1 vccd1 _10581_/A sky130_fd_sc_hd__or2_1
XFILLER_0_121_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13298_ _13309_/CLK _13298_/D vssd1 vssd1 vccd1 vccd1 hold260/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__08223__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12318_ _11973_/B _12317_/A _12221_/X _12317_/B _11973_/A vssd1 vssd1 vccd1 vccd1
+ _12319_/B sky130_fd_sc_hd__a41o_1
XFILLER_0_121_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12249_ _12224_/X _12229_/X _12232_/Y _12248_/X _06930_/Y vssd1 vssd1 vccd1 vccd1
+ _12249_/X sky130_fd_sc_hd__a41o_1
XANTENNA__07359__B1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07790_ _07790_/A _07790_/B _07790_/C vssd1 vssd1 vccd1 vccd1 _07802_/A sky130_fd_sc_hd__or3_1
X_06810_ _10863_/A _06808_/Y _06809_/X vssd1 vssd1 vccd1 vccd1 _06810_/X sky130_fd_sc_hd__a21o_1
X_06741_ _06783_/A _06649_/A _12598_/B _06740_/X vssd1 vssd1 vccd1 vccd1 _06986_/A
+ sky130_fd_sc_hd__a31o_4
XANTENNA__08323__A2 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09460_ _09461_/A _09461_/B vssd1 vssd1 vccd1 vccd1 _09462_/A sky130_fd_sc_hd__or2_1
X_06672_ _06670_/Y _06680_/B1 _06752_/A reg2_val[18] vssd1 vssd1 vccd1 vccd1 _07023_/A
+ sky130_fd_sc_hd__a2bb2o_2
X_08411_ _09452_/A _08411_/B vssd1 vssd1 vccd1 vccd1 _08413_/B sky130_fd_sc_hd__xnor2_2
X_09391_ _09192_/Y _09381_/Y _09382_/X _09390_/X _09379_/Y vssd1 vssd1 vccd1 vccd1
+ _09391_/X sky130_fd_sc_hd__a311o_1
XANTENNA__07005__C _07005_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__A1 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08087__B2 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08342_ _08342_/A _08342_/B vssd1 vssd1 vccd1 vccd1 _08343_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_86_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13080__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08273_ _07134_/A _12752_/A fanout84/X _08758_/A2 vssd1 vssd1 vccd1 vccd1 _08274_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10969__A1 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout134_A _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ _07379_/A _07379_/B _07210_/Y vssd1 vssd1 vccd1 vccd1 _07423_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07155_ _07149_/A _07149_/B _08443_/A vssd1 vssd1 vccd1 vccd1 _07155_/X sky130_fd_sc_hd__mux2_2
XANTENNA__10197__A2 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ reg1_val[26] reg1_val[27] _07086_/C vssd1 vssd1 vccd1 vccd1 _12697_/B sky130_fd_sc_hd__or3_2
XANTENNA__09229__A _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout101 _07167_/Y vssd1 vssd1 vccd1 vccd1 _09925_/A1 sky130_fd_sc_hd__clkbuf_8
Xfanout112 _09926_/A vssd1 vssd1 vccd1 vccd1 _11604_/A sky130_fd_sc_hd__buf_12
XFILLER_0_1_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout156 _12230_/A vssd1 vssd1 vccd1 vccd1 _11559_/A sky130_fd_sc_hd__clkbuf_4
Xfanout123 _07324_/Y vssd1 vssd1 vccd1 vccd1 _08835_/B1 sky130_fd_sc_hd__clkbuf_8
Xfanout145 _06974_/X vssd1 vssd1 vccd1 vccd1 _10144_/B2 sky130_fd_sc_hd__buf_6
Xfanout134 _10156_/B2 vssd1 vssd1 vccd1 vccd1 _08477_/B sky130_fd_sc_hd__clkbuf_8
Xfanout178 _12723_/Y vssd1 vssd1 vccd1 vccd1 _12781_/A2 sky130_fd_sc_hd__buf_4
X_07988_ _07995_/A vssd1 vssd1 vccd1 vccd1 _07988_/Y sky130_fd_sc_hd__inv_2
Xfanout167 _07110_/Y vssd1 vssd1 vccd1 vccd1 _08774_/A2 sky130_fd_sc_hd__buf_4
Xfanout189 _07075_/B vssd1 vssd1 vccd1 vccd1 _07135_/B sky130_fd_sc_hd__buf_4
X_06939_ reg1_val[18] reg1_val[19] _06939_/C vssd1 vssd1 vccd1 vccd1 _12658_/B sky130_fd_sc_hd__or3_4
X_09727_ _08821_/B _09295_/B _10433_/A fanout36/X vssd1 vssd1 vccd1 vccd1 _09728_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout47_A _07852_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07522__B1 _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ _09659_/A _09659_/B vssd1 vssd1 vccd1 vccd1 _09658_/X sky130_fd_sc_hd__and2_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08609_ _08609_/A _08609_/B vssd1 vssd1 vccd1 vccd1 _09047_/B sky130_fd_sc_hd__xnor2_1
X_09589_ _09736_/B _09589_/B vssd1 vssd1 vccd1 vccd1 _09592_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12949__A2 _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10409__B1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11620_ _11620_/A _11620_/B vssd1 vssd1 vccd1 vccd1 _11622_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08308__A _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11082__B1 _12228_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07212__A _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10557__B _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11551_ _11371_/X _11552_/B _11549_/X vssd1 vssd1 vccd1 vccd1 _11551_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10502_ reg1_val[9] curr_PC[9] vssd1 vssd1 vccd1 vccd1 _10503_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_65_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11482_ hold168/A _12187_/A1 _11573_/B _11481_/Y _11920_/C1 vssd1 vssd1 vccd1 vccd1
+ _11490_/A sky130_fd_sc_hd__a311o_1
XFILLER_0_18_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13221_ _13248_/CLK _13221_/D vssd1 vssd1 vccd1 vccd1 hold224/A sky130_fd_sc_hd__dfxtp_1
X_10433_ _10433_/A _12349_/B _10433_/C _10433_/D vssd1 vssd1 vccd1 vccd1 _10435_/B
+ sky130_fd_sc_hd__or4_1
X_13152_ _13166_/A hold255/X vssd1 vssd1 vccd1 vccd1 _13308_/D sky130_fd_sc_hd__and2_1
XFILLER_0_20_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_747 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10364_ _10097_/Y _10609_/C _10363_/Y vssd1 vssd1 vccd1 vccd1 _10851_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_103_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ _11966_/Y _12101_/X _12100_/Y vssd1 vssd1 vccd1 vccd1 _12103_/X sky130_fd_sc_hd__a21o_1
X_13083_ _13083_/A _13083_/B vssd1 vssd1 vccd1 vccd1 _13083_/Y sky130_fd_sc_hd__xnor2_1
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10295_ _10295_/A _10295_/B vssd1 vssd1 vccd1 vccd1 _10297_/B sky130_fd_sc_hd__xnor2_1
X_12034_ _12036_/A _12036_/B _12036_/C vssd1 vssd1 vccd1 vccd1 _12035_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_18_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09750__B2 fanout75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09750__A1 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12936_ _12946_/A hold222/X vssd1 vssd1 vccd1 vccd1 hold223/A sky130_fd_sc_hd__and2_1
XANTENNA__07513__B1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12867_ _12804_/X _12867_/B vssd1 vssd1 vccd1 vccd1 _13117_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11818_ _11768_/X _11972_/C _11817_/Y vssd1 vssd1 vccd1 vccd1 _11818_/X sky130_fd_sc_hd__a21o_1
XANTENNA__08218__A _08857_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12798_ _12796_/X _12798_/B vssd1 vssd1 vccd1 vccd1 _13144_/A sky130_fd_sc_hd__nand2b_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07816__A1 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11749_ _12119_/B1 _11832_/B hold252/A vssd1 vssd1 vccd1 vccd1 _11749_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__07816__B2 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10820__B1 _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10179__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08960_ _08960_/A _08960_/B vssd1 vssd1 vccd1 vccd1 _08963_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__12325__B1 _12278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07911_ _07134_/A _12762_/A _12760_/A _07869_/B vssd1 vssd1 vccd1 vccd1 _07912_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08891_ _08891_/A _08891_/B _08891_/C vssd1 vssd1 vccd1 vccd1 _08892_/B sky130_fd_sc_hd__or3_1
X_07842_ _07842_/A _07842_/B vssd1 vssd1 vccd1 vccd1 _07844_/B sky130_fd_sc_hd__xor2_2
XANTENNA__09741__B2 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__A1 _10557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12203__A _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07773_ _09252_/A _07179_/A _11012_/A _09253_/A vssd1 vssd1 vccd1 vccd1 _07774_/B
+ sky130_fd_sc_hd__a22o_1
X_09512_ _09403_/X _09559_/D _12223_/B1 vssd1 vssd1 vccd1 vccd1 _09512_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06724_ _06783_/A _06641_/A _12614_/B _06723_/X vssd1 vssd1 vccd1 vccd1 _07319_/A
+ sky130_fd_sc_hd__a31o_4
X_06655_ instruction[0] instruction[1] instruction[2] instruction[31] pred_val vssd1
+ vssd1 vccd1 vccd1 _12588_/B sky130_fd_sc_hd__o311a_4
XFILLER_0_78_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09443_ _09444_/A _09444_/B vssd1 vssd1 vccd1 vccd1 _09575_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__10658__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09374_ _09374_/A _09374_/B vssd1 vssd1 vccd1 vccd1 _09375_/B sky130_fd_sc_hd__xnor2_1
X_06586_ instruction[38] _06633_/B vssd1 vssd1 vccd1 vccd1 _12626_/B sky130_fd_sc_hd__and2_4
X_08325_ _12734_/A _08477_/B _08776_/B1 _08819_/B2 vssd1 vssd1 vccd1 vccd1 _08326_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10377__B _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07807__B2 _08772_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07807__A1 _08772_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08256_ _08259_/A _08259_/B vssd1 vssd1 vccd1 vccd1 _08256_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12592__B _12593_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08187_ _08855_/A _08187_/B vssd1 vssd1 vccd1 vccd1 _08190_/A sky130_fd_sc_hd__xnor2_2
X_07207_ _09452_/A _07207_/B vssd1 vssd1 vccd1 vccd1 _07209_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06590__B _12250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07138_ _07139_/A _07139_/B vssd1 vssd1 vccd1 vccd1 _07138_/X sky130_fd_sc_hd__and2_2
XFILLER_0_15_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07069_ _07821_/B _07821_/C vssd1 vssd1 vccd1 vccd1 _07069_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07991__B1 _08774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10080_ _09876_/A _09876_/B _09874_/Y vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__07743__B1 _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07207__A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10982_ _10978_/Y _10981_/Y _11197_/S vssd1 vssd1 vccd1 vccd1 _10982_/X sky130_fd_sc_hd__mux2_1
X_12721_ rst _12721_/B _12721_/C vssd1 vssd1 vccd1 vccd1 _13183_/D sky130_fd_sc_hd__nor3_1
XFILLER_0_97_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06765__B _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12652_ _12657_/C _12652_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[18] sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11603_ _11603_/A fanout8/X vssd1 vssd1 vccd1 vccd1 _11604_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_80_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ reg1_val[5] _12583_/B vssd1 vssd1 vccd1 vccd1 _12584_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07877__A _07974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06781__A _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11534_ _11532_/A _11532_/B _11535_/B vssd1 vssd1 vccd1 vccd1 _11534_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11465_ _11406_/X _11586_/A _12223_/B1 vssd1 vssd1 vccd1 vccd1 _11465_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13204_ _13303_/CLK _13204_/D vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_111_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10416_ _10416_/A _10416_/B vssd1 vssd1 vccd1 vccd1 _10418_/A sky130_fd_sc_hd__and2_1
XFILLER_0_110_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11396_ _12373_/A1 _11092_/Y _11391_/B _09183_/Y _11395_/X vssd1 vssd1 vccd1 vccd1
+ _11404_/C sky130_fd_sc_hd__a221o_1
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13135_ _13135_/A _13135_/B vssd1 vssd1 vccd1 vccd1 _13135_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__08774__A2 _08774_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10347_ _10346_/A _10346_/B _10348_/A vssd1 vssd1 vccd1 vccd1 _10347_/X sky130_fd_sc_hd__o21a_1
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ _13066_/A hold273/X vssd1 vssd1 vccd1 vccd1 _13290_/D sky130_fd_sc_hd__and2_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10278_ _10551_/B _10278_/B vssd1 vssd1 vccd1 vccd1 _10284_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12017_ _12206_/A _12017_/B vssd1 vssd1 vccd1 vccd1 _12019_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12086__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12919_ hold195/X _12947_/A2 _12947_/B1 hold215/X vssd1 vssd1 vccd1 vccd1 hold216/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08110_ _08165_/A _08165_/B vssd1 vssd1 vccd1 vccd1 _08166_/A sky130_fd_sc_hd__or2_1
XANTENNA__06691__A _12641_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09090_ _09090_/A _09090_/B _09103_/B vssd1 vssd1 vccd1 vccd1 _09092_/A sky130_fd_sc_hd__and3_1
XFILLER_0_28_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08041_ _08837_/B2 _08348_/B _07181_/Y _07969_/A vssd1 vssd1 vccd1 vccd1 _08042_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10925__B _10925_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09992_ _09992_/A _09992_/B vssd1 vssd1 vccd1 vccd1 _09992_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07973__B1 fanout47/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__B wire201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08943_ _08944_/A _08944_/B vssd1 vssd1 vccd1 vccd1 _08945_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08411__A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout299_A _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08517__A2 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__A1 _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08874_ _08792_/A _08792_/B _08790_/Y vssd1 vssd1 vccd1 vccd1 _08876_/B sky130_fd_sc_hd__a21o_1
X_07825_ _07825_/A _07825_/B _07825_/C vssd1 vssd1 vccd1 vccd1 _07829_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_79_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07756_ _07756_/A _07756_/B vssd1 vssd1 vccd1 vccd1 _07782_/A sky130_fd_sc_hd__nor2_2
XANTENNA__11772__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09478__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06707_ _06898_/A _06641_/A _12632_/B _06706_/X vssd1 vssd1 vccd1 vccd1 _07197_/A
+ sky130_fd_sc_hd__a31o_4
XFILLER_0_67_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12587__B _12588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07687_ _07687_/A _07687_/B _08904_/A vssd1 vssd1 vccd1 vccd1 _07688_/B sky130_fd_sc_hd__or3_1
X_09426_ _10555_/A _09426_/B vssd1 vssd1 vccd1 vccd1 _09428_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__06700__A1 _06898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06638_ reg1_val[23] _07112_/A vssd1 vssd1 vccd1 vccd1 _06639_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06569_ instruction[0] instruction[2] instruction[1] pred_val vssd1 vssd1 vccd1 vccd1
+ _06569_/X sky130_fd_sc_hd__or4bb_4
XFILLER_0_81_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09357_ _09151_/X _09154_/X _09359_/S vssd1 vssd1 vccd1 vccd1 _09357_/X sky130_fd_sc_hd__mux2_1
X_08308_ _08394_/A _08308_/B _08308_/C vssd1 vssd1 vccd1 vccd1 _08309_/C sky130_fd_sc_hd__or3_1
XFILLER_0_35_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09288_ _09288_/A _09288_/B vssd1 vssd1 vccd1 vccd1 _09289_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_105_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08239_ _08235_/A _08235_/B _08238_/Y vssd1 vssd1 vccd1 vccd1 _08264_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11012__A _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11250_ _11250_/A _11250_/B vssd1 vssd1 vccd1 vccd1 _11251_/B sky130_fd_sc_hd__and2_1
XFILLER_0_113_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08756__A2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10201_ _10201_/A _10201_/B vssd1 vssd1 vccd1 vccd1 _10204_/A sky130_fd_sc_hd__nor2_1
X_11181_ _11110_/X _11215_/D _11180_/Y vssd1 vssd1 vccd1 vccd1 _11181_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10132_ _10132_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _10132_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__09705__A1 _06964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10063_ _10280_/A _10063_/B vssd1 vssd1 vccd1 vccd1 _10071_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_89_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12704_ _12704_/A _12704_/B vssd1 vssd1 vccd1 vccd1 _12706_/A sky130_fd_sc_hd__nand2_2
X_10965_ _11173_/A _10965_/B vssd1 vssd1 vccd1 vccd1 _11215_/B sky130_fd_sc_hd__xor2_2
XANTENNA__08692__A1 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08692__B2 _12768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10896_ _11125_/A _10896_/B vssd1 vssd1 vccd1 vccd1 _10898_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12635_ _12635_/A _12635_/B _12635_/C vssd1 vssd1 vccd1 vccd1 _12636_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12566_ _12565_/A _12565_/B _12564_/B vssd1 vssd1 vccd1 vccd1 _12570_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11517_ _11794_/A _12205_/A _12772_/A fanout27/X vssd1 vssd1 vccd1 vccd1 _11518_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12497_ _12551_/A _12498_/B vssd1 vssd1 vccd1 vccd1 _12516_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12018__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold209 hold209/A vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11448_ _11449_/A _11449_/B vssd1 vssd1 vccd1 vccd1 _11544_/A sky130_fd_sc_hd__and2b_1
X_11379_ _11379_/A _11379_/B _11379_/C vssd1 vssd1 vccd1 vccd1 _11381_/B sky130_fd_sc_hd__or3_1
XFILLER_0_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13118_ hold280/A _13117_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13118_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10554__A2 _11782_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ hold284/A _13048_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13049_/X sky130_fd_sc_hd__mux2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07183__A1 _11222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07183__B2 _07182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08590_ _08592_/A _08591_/B vssd1 vssd1 vccd1 vccd1 _08597_/A sky130_fd_sc_hd__nor2_1
X_07610_ _07611_/A _07611_/B vssd1 vssd1 vccd1 vccd1 _07610_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_88_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07541_ _07541_/A _07541_/B vssd1 vssd1 vccd1 vccd1 _07542_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_49_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13008__A1 _11780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07472_ _07472_/A _07472_/B vssd1 vssd1 vccd1 vccd1 _07475_/A sky130_fd_sc_hd__nand2_1
X_09211_ _09211_/A _09211_/B vssd1 vssd1 vccd1 vccd1 _11195_/B sky130_fd_sc_hd__and2_1
XFILLER_0_8_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11019__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09142_ reg1_val[15] reg1_val[16] _09172_/S vssd1 vssd1 vccd1 vccd1 _09142_/X sky130_fd_sc_hd__mux2_1
XANTENNA__07238__A2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09227__A3 _07526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10242__A1 _06866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09073_ _11559_/B _11559_/C _09073_/C _09073_/D vssd1 vssd1 vccd1 vccd1 _11820_/B
+ sky130_fd_sc_hd__or4_2
XANTENNA_fanout214_A _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08024_ _08024_/A _08024_/B vssd1 vssd1 vccd1 vccd1 _08060_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_114_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09975_ _09973_/X _09974_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _09975_/X sky130_fd_sc_hd__mux2_1
X_08926_ _08927_/B _08927_/A vssd1 vssd1 vccd1 vccd1 _08926_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__09699__B1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12298__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08857_ _08857_/A _08857_/B vssd1 vssd1 vccd1 vccd1 _08859_/B sky130_fd_sc_hd__xnor2_1
X_07808_ _08773_/A _07808_/B vssd1 vssd1 vccd1 vccd1 _07809_/B sky130_fd_sc_hd__xnor2_2
X_08788_ _08689_/A _08689_/C _08689_/B vssd1 vssd1 vccd1 vccd1 _08791_/A sky130_fd_sc_hd__a21boi_2
X_07739_ _07738_/A _07738_/B _07738_/C vssd1 vssd1 vccd1 vccd1 _07754_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10750_ _09674_/X _09680_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _10751_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09871__B1 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12537__S _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10681_ _11695_/A _10681_/B vssd1 vssd1 vccd1 vccd1 _10683_/C sky130_fd_sc_hd__xnor2_1
X_09409_ _08680_/B _09295_/B _10433_/A fanout30/X vssd1 vssd1 vccd1 vccd1 _09410_/B
+ sky130_fd_sc_hd__o22a_1
X_12420_ _12429_/A _12420_/B vssd1 vssd1 vccd1 vccd1 _12422_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08316__A _10453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09623__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12351_ _12266_/B _12269_/X _12309_/X _12311_/A vssd1 vssd1 vccd1 vccd1 _12352_/B
+ sky130_fd_sc_hd__o31a_1
X_11302_ hold239/A _11302_/B vssd1 vssd1 vccd1 vccd1 _11480_/C sky130_fd_sc_hd__or2_1
X_12282_ reg1_val[28] _12281_/C reg1_val[29] vssd1 vssd1 vccd1 vccd1 _12282_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__10784__A2 fanout52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08729__A2 _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11233_ _12022_/A _11233_/B vssd1 vssd1 vccd1 vccd1 _11234_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__10536__A2 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11164_ _11164_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11166_/B sky130_fd_sc_hd__xnor2_1
X_11095_ hold180/A _11095_/B vssd1 vssd1 vccd1 vccd1 _11095_/Y sky130_fd_sc_hd__xnor2_1
X_10115_ _09527_/X _09530_/X _10249_/S vssd1 vssd1 vccd1 vccd1 _11089_/B sky130_fd_sc_hd__mux2_1
XANTENNA__07890__A _08855_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10046_ _10557_/A fanout95/X fanout54/X fanout62/X vssd1 vssd1 vccd1 vccd1 _10047_/B
+ sky130_fd_sc_hd__o22a_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12301__A _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11997_ _07126_/B _12250_/B _10377_/B reg1_val[24] vssd1 vssd1 vccd1 vccd1 _11997_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_58_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08665__B2 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08665__A1 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07468__A2 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10948_ _10949_/B _10949_/A vssd1 vssd1 vccd1 vccd1 _10948_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_45_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09610__A _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10879_ hold274/A _09842_/B _10986_/B _12339_/B1 vssd1 vssd1 vccd1 vccd1 _10879_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08226__A _08311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12618_ _12623_/B _12618_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[11] sky130_fd_sc_hd__and2_4
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12549_ reg1_val[26] curr_PC[26] _12556_/S vssd1 vssd1 vccd1 vccd1 _12551_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _07073_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ _06986_/A _06996_/A _06972_/C _07001_/C vssd1 vssd1 vccd1 vccd1 _07175_/B
+ sky130_fd_sc_hd__or4_4
X_09760_ _10578_/A _09760_/B vssd1 vssd1 vccd1 vccd1 _09761_/B sky130_fd_sc_hd__xnor2_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _08712_/A _08712_/B vssd1 vssd1 vccd1 vccd1 _08711_/Y sky130_fd_sc_hd__nor2_1
X_09691_ _11194_/S _09690_/X _11195_/C vssd1 vssd1 vccd1 vccd1 _09691_/X sky130_fd_sc_hd__o21a_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08642_ _09076_/A _09074_/B vssd1 vssd1 vccd1 vccd1 _08642_/X sky130_fd_sc_hd__and2_1
XANTENNA__06636__A2_N _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07156__A1 _07126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout164_A _07116_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08573_ _09898_/A _08583_/B _08572_/X vssd1 vssd1 vccd1 vccd1 _08602_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07524_ _07524_/A _07524_/B vssd1 vssd1 vccd1 vccd1 _07525_/B sky130_fd_sc_hd__xor2_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11660__B1 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07455_ _10452_/B2 fanout75/X _10553_/B _10527_/A vssd1 vssd1 vccd1 vccd1 _07456_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_107_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06863__B _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10666__A _12022_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08408__A1 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08408__B2 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07386_ _07694_/A _07694_/B _07382_/X vssd1 vssd1 vccd1 vccd1 _07417_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09125_ _09123_/X _09124_/X _09365_/S vssd1 vssd1 vccd1 vccd1 _09125_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11412__B1 _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09056_ _10740_/B _10740_/C _10859_/A vssd1 vssd1 vccd1 vccd1 _09059_/A sky130_fd_sc_hd__and3_1
XFILLER_0_115_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08007_ _08007_/A _08007_/B vssd1 vssd1 vccd1 vccd1 _08008_/B sky130_fd_sc_hd__xor2_4
XANTENNA__11497__A _11853_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09958_ _09958_/A _09958_/B vssd1 vssd1 vccd1 vccd1 _10229_/C sky130_fd_sc_hd__xnor2_4
X_08909_ _08908_/A _08908_/B _08908_/C vssd1 vssd1 vccd1 vccd1 _08910_/C sky130_fd_sc_hd__a21o_1
XANTENNA_fanout77_A _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09889_ _10551_/B _09889_/B vssd1 vssd1 vccd1 vccd1 _09891_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12140__A1 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12140__B2 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11920_ hold226/A _12187_/A1 _11992_/B _11919_/Y _11920_/C1 vssd1 vssd1 vccd1 vccd1
+ _11920_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_87_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11851_ _12143_/A _11851_/B vssd1 vssd1 vccd1 vccd1 _11853_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__08647__A1 _10156_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11782_ _11782_/A fanout8/X vssd1 vssd1 vccd1 vccd1 _11783_/C sky130_fd_sc_hd__nor2_1
X_10802_ _10802_/A _10802_/B vssd1 vssd1 vccd1 vccd1 _10805_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08647__B2 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10733_ _10230_/X _10231_/X _10233_/Y _10732_/Y vssd1 vssd1 vccd1 vccd1 _10734_/C
+ sky130_fd_sc_hd__a31o_2
XANTENNA__09430__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07869__B _07869_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10576__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08046__A _08821_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10664_ _10664_/A _10664_/B vssd1 vssd1 vccd1 vccd1 _10710_/A sky130_fd_sc_hd__xnor2_1
X_12403_ reg1_val[4] curr_PC[4] _12524_/S vssd1 vssd1 vccd1 vccd1 _12405_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_63_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10595_ _10595_/A _10595_/B vssd1 vssd1 vccd1 vccd1 _10596_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_121_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12334_ _06631_/A wire201/X _09202_/B reg1_val[30] vssd1 vssd1 vccd1 vccd1 _12334_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_51_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12265_ _12264_/A _12264_/B _12264_/C vssd1 vssd1 vccd1 vccd1 _12266_/B sky130_fd_sc_hd__o21a_1
X_12196_ _12168_/X _12172_/X _12195_/X _12139_/Y _12382_/S vssd1 vssd1 vccd1 vccd1
+ dest_val[27] sky130_fd_sc_hd__o32a_4
X_11216_ _11000_/A _11316_/A _11316_/C _12278_/A vssd1 vssd1 vccd1 vccd1 _11216_/X
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_128_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11147_ _11147_/A _11147_/B vssd1 vssd1 vccd1 vccd1 _11148_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_37_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11078_ _09059_/C _11077_/X _11184_/A vssd1 vssd1 vccd1 vccd1 _11078_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__06948__B _10249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10029_ _10030_/A _10030_/B _10030_/C vssd1 vssd1 vccd1 vccd1 _10212_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__07125__A _07157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11870__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06964__A _06964_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11081__S _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10996__A2 _10995_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11642__B1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07861__A2 _12752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07240_ _07240_/A vssd1 vssd1 vccd1 vccd1 _07250_/A sky130_fd_sc_hd__inv_2
XFILLER_0_27_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07171_ _08855_/A _07172_/B vssd1 vssd1 vccd1 vccd1 _07180_/B sky130_fd_sc_hd__and2_1
XANTENNA__07795__A _11604_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12206__A _12206_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout305 _09198_/C vssd1 vssd1 vccd1 vccd1 _09200_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__07019__B _07192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09812_ _09814_/A _09814_/B vssd1 vssd1 vccd1 vccd1 _09812_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout281_A _06569_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06955_ reg1_val[25] _06955_/B vssd1 vssd1 vccd1 vccd1 _07364_/A sky130_fd_sc_hd__xor2_4
X_09743_ _10156_/B2 _07132_/Y fanout22/X _10156_/A1 vssd1 vssd1 vccd1 vccd1 _09744_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09674_ _09672_/X _09673_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09674_/X sky130_fd_sc_hd__mux2_1
X_06886_ _09200_/A _09200_/B vssd1 vssd1 vccd1 vccd1 _09199_/B sky130_fd_sc_hd__nand2_8
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _08295_/X _08626_/B vssd1 vssd1 vccd1 vccd1 _09070_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10684__B2 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10684__A1 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _08549_/A _08549_/B _08549_/C vssd1 vssd1 vccd1 vccd1 _08559_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__11780__A _11780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09826__B1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07507_ _10553_/B fanout98/X fanout56/X fanout69/X vssd1 vssd1 vccd1 vccd1 _07508_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__06593__B _06633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08487_ _08487_/A _08487_/B vssd1 vssd1 vccd1 vccd1 _08488_/B sky130_fd_sc_hd__and2_1
XFILLER_0_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07438_ _08595_/A _07438_/B vssd1 vssd1 vccd1 vccd1 _07440_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07369_ _10565_/A _07369_/B vssd1 vssd1 vccd1 vccd1 _07371_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09108_ _09559_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09108_/Y sky130_fd_sc_hd__nand2_1
X_10380_ hold268/A _10381_/B vssd1 vssd1 vccd1 vccd1 _10380_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_102_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ _09039_/A _09039_/B vssd1 vssd1 vccd1 vccd1 _09040_/B sky130_fd_sc_hd__xor2_2
X_12050_ reg1_val[25] curr_PC[25] vssd1 vssd1 vccd1 vccd1 _12050_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11020__A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07368__B2 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07368__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ _10947_/A _10947_/B _10948_/Y vssd1 vssd1 vccd1 vccd1 _11064_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__10911__A2 _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06768__B _11194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12952_ _13169_/A hold166/X vssd1 vssd1 vccd1 vccd1 hold167/A sky130_fd_sc_hd__and2_1
XFILLER_0_87_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11903_ _11824_/A _11822_/X _06830_/Y _11823_/S vssd1 vssd1 vccd1 vccd1 _11903_/X
+ sky130_fd_sc_hd__o211a_1
X_12883_ _13148_/A _13149_/A _13148_/B vssd1 vssd1 vccd1 vccd1 _13153_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__12786__A _12786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ hold293/A _12119_/B1 _11989_/C _11833_/Y _11400_/A vssd1 vssd1 vccd1 vccd1
+ _11834_/X sky130_fd_sc_hd__a311o_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11765_ _12556_/S _11765_/B _11929_/C vssd1 vssd1 vccd1 vccd1 _11765_/X sky130_fd_sc_hd__or3_2
XFILLER_0_28_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11696_ fanout33/X _12301_/A fanout8/X _10553_/A vssd1 vssd1 vccd1 vccd1 _11697_/B
+ sky130_fd_sc_hd__o22a_1
X_10716_ _10571_/A _10571_/B _10569_/Y vssd1 vssd1 vccd1 vccd1 _10718_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_126_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10647_ curr_PC[9] _10646_/C curr_PC[10] vssd1 vssd1 vccd1 vccd1 _10648_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10578_ _10578_/A _10578_/B vssd1 vssd1 vccd1 vccd1 _10580_/B sky130_fd_sc_hd__xnor2_2
X_13297_ _13309_/CLK _13297_/D vssd1 vssd1 vccd1 vccd1 hold294/A sky130_fd_sc_hd__dfxtp_1
X_12317_ _12317_/A _12317_/B vssd1 vssd1 vccd1 vccd1 _12317_/X sky130_fd_sc_hd__and2_1
XFILLER_0_121_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12248_ _12238_/Y _12239_/X _12247_/X _12236_/X vssd1 vssd1 vccd1 vccd1 _12248_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__07359__B2 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07359__A1 fanout36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ _12179_/A _12179_/B vssd1 vssd1 vccd1 vccd1 _12179_/Y sky130_fd_sc_hd__nor2_1
X_06740_ reg2_val[7] _06778_/B vssd1 vssd1 vccd1 vccd1 _06740_/X sky130_fd_sc_hd__and2_1
XFILLER_0_64_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06671_ reg2_val[18] _06752_/A _06680_/B1 _06670_/Y vssd1 vssd1 vccd1 vccd1 _07075_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_08410_ _08776_/B1 _08748_/B1 _12730_/A _08477_/B vssd1 vssd1 vccd1 vccd1 _08411_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09390_ _09544_/A _10638_/B _09383_/Y _09389_/X vssd1 vssd1 vccd1 vccd1 _09390_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13080__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08341_ _08341_/A _08341_/B vssd1 vssd1 vccd1 vccd1 _08619_/A sky130_fd_sc_hd__xor2_4
XANTENNA__08087__A2 fanout82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08272_ _08775_/A _08272_/B vssd1 vssd1 vccd1 vccd1 _08278_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07223_ _07632_/A _07223_/B vssd1 vssd1 vccd1 vccd1 _07379_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__09036__A1 _08589_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout127_A _07894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07154_ _07150_/A _07150_/B _08443_/A vssd1 vssd1 vccd1 vccd1 _07154_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_42_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11394__A2 _06928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07085_ _07409_/A _07409_/B _07065_/Y vssd1 vssd1 vccd1 vccd1 _07162_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09339__A2 _12131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout102 _10527_/A vssd1 vssd1 vccd1 vccd1 _08854_/B2 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08547__B1 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout113 _06999_/A vssd1 vssd1 vccd1 vccd1 _11853_/A sky130_fd_sc_hd__clkbuf_16
Xfanout124 _07319_/Y vssd1 vssd1 vccd1 vccd1 _09295_/B sky130_fd_sc_hd__buf_8
Xfanout146 _09772_/A vssd1 vssd1 vccd1 vccd1 _12734_/A sky130_fd_sc_hd__buf_6
Xfanout135 _07073_/X vssd1 vssd1 vccd1 vccd1 _10156_/B2 sky130_fd_sc_hd__buf_6
Xfanout179 _12742_/B vssd1 vssd1 vccd1 vccd1 _12778_/B sky130_fd_sc_hd__buf_4
X_07987_ _08443_/A _07987_/B vssd1 vssd1 vccd1 vccd1 _07995_/A sky130_fd_sc_hd__xnor2_4
Xfanout168 _08748_/B1 vssd1 vssd1 vccd1 vccd1 _08825_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout157 _09002_/X vssd1 vssd1 vccd1 vccd1 _12230_/A sky130_fd_sc_hd__buf_4
X_06938_ reg1_val[16] reg1_val[17] vssd1 vssd1 vccd1 vccd1 _06939_/C sky130_fd_sc_hd__or2_2
X_09726_ _09726_/A _09726_/B vssd1 vssd1 vccd1 vccd1 _09729_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_96_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06869_ _08594_/B _06864_/Y _10373_/A vssd1 vssd1 vccd1 vccd1 _06870_/D sky130_fd_sc_hd__a21oi_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07522__A1 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ _09659_/A _09659_/B vssd1 vssd1 vccd1 vccd1 _09657_/X sky130_fd_sc_hd__or2_1
XFILLER_0_96_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ _08553_/X _08608_/B vssd1 vssd1 vccd1 vccd1 _09045_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_49_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09588_ _09588_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09589_/B sky130_fd_sc_hd__and2_1
XFILLER_0_65_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08539_ _08609_/A _08609_/B vssd1 vssd1 vccd1 vccd1 _09049_/A sky130_fd_sc_hd__or2_1
XFILLER_0_49_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10409__A1 fanout22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10409__B2 _12150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07286__B1 _07553_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11550_ _11550_/A _11635_/A vssd1 vssd1 vccd1 vccd1 _11552_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10501_ reg1_val[9] curr_PC[9] vssd1 vssd1 vccd1 vccd1 _10501_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout6_A fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11481_ _12187_/A1 _11573_/B hold168/A vssd1 vssd1 vccd1 vccd1 _11481_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13220_ _13248_/CLK _13220_/D vssd1 vssd1 vccd1 vccd1 hold237/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08324__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10432_ _10432_/A _10432_/B vssd1 vssd1 vccd1 vccd1 _10448_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13151_ hold254/X _13151_/A2 _13150_/X _13168_/A2 vssd1 vssd1 vccd1 vccd1 hold255/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10363_ _10092_/X _10225_/X _10226_/X vssd1 vssd1 vccd1 vccd1 _10363_/Y sky130_fd_sc_hd__a21oi_1
X_13082_ _13082_/A _13082_/B vssd1 vssd1 vccd1 vccd1 _13083_/B sky130_fd_sc_hd__nand2_1
X_12102_ _12102_/A _12102_/B _12102_/C vssd1 vssd1 vccd1 vccd1 _12216_/C sky130_fd_sc_hd__or3_1
XFILLER_0_21_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12033_ _12098_/B _12033_/B vssd1 vssd1 vccd1 vccd1 _12036_/C sky130_fd_sc_hd__nand2_1
X_10294_ _10295_/A _10295_/B vssd1 vssd1 vccd1 vccd1 _10420_/A sky130_fd_sc_hd__and2b_1
XANTENNA__09750__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12935_ hold234/A _12947_/A2 _13168_/B1 hold221/X vssd1 vssd1 vccd1 vccd1 hold222/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11845__B1 _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07513__B2 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07513__A1 _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12866_ hold280/A hold23/X vssd1 vssd1 vccd1 vccd1 _12867_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_87_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11817_ _11768_/X _11972_/C _12223_/B1 vssd1 vssd1 vccd1 vccd1 _11817_/Y sky130_fd_sc_hd__o21ai_1
X_12797_ hold286/A hold79/X vssd1 vssd1 vccd1 vccd1 _12798_/B sky130_fd_sc_hd__nand2b_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11748_ hold277/A _11748_/B vssd1 vssd1 vccd1 vccd1 _11832_/B sky130_fd_sc_hd__or2_1
XANTENNA__07816__A2 _08217_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11679_ _11680_/A _11680_/B vssd1 vssd1 vccd1 vccd1 _11777_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08234__A _08773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_247 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07910_ _07928_/A _07928_/B vssd1 vssd1 vccd1 vccd1 _07910_/Y sky130_fd_sc_hd__nand2b_1
X_08890_ _08891_/A _08891_/B _08891_/C vssd1 vssd1 vccd1 vccd1 _08949_/A sky130_fd_sc_hd__o21ai_1
X_07841_ _07841_/A _07841_/B vssd1 vssd1 vccd1 vccd1 _07883_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__07201__B1 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09741__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ _08855_/A _07772_/B vssd1 vssd1 vccd1 vccd1 _07775_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12203__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06723_ reg2_val[10] _06729_/B vssd1 vssd1 vccd1 vccd1 _06723_/X sky130_fd_sc_hd__and2_1
X_09511_ _09816_/A _09511_/B vssd1 vssd1 vccd1 vccd1 _09559_/D sky130_fd_sc_hd__xnor2_2
XANTENNA__11300__A2 wire201/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08409__A _08775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06654_ _06654_/A _06654_/B vssd1 vssd1 vccd1 vccd1 _06661_/C sky130_fd_sc_hd__and2_1
X_09442_ _09442_/A _09442_/B vssd1 vssd1 vccd1 vccd1 _09444_/B sky130_fd_sc_hd__xnor2_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09373_ _09373_/A _09373_/B vssd1 vssd1 vccd1 vccd1 _09374_/B sky130_fd_sc_hd__nor2_1
X_06585_ _06583_/X _06585_/B vssd1 vssd1 vccd1 vccd1 _12276_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_47_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08324_ _08773_/A _08324_/B vssd1 vssd1 vccd1 vccd1 _08359_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout244_A _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07268__B1 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07807__A2 fanout94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08255_ _08255_/A _08255_/B vssd1 vssd1 vccd1 vccd1 _08259_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08186_ _07969_/A _08420_/B _08854_/B2 _12734_/A vssd1 vssd1 vccd1 vccd1 _08187_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_61_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07206_ _11704_/A _10156_/B2 _10156_/A1 _11688_/A vssd1 vssd1 vccd1 vccd1 _07207_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07137_ _07127_/X _07130_/Y _07136_/X _07135_/B vssd1 vssd1 vccd1 vccd1 _07139_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_42_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10575__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07991__A1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ _07068_/A _07135_/B _07128_/B vssd1 vssd1 vccd1 vccd1 _07821_/C sky130_fd_sc_hd__or3_1
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07991__B2 _12762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10981_ _11195_/A _09518_/Y _10980_/X vssd1 vssd1 vccd1 vccd1 _10981_/Y sky130_fd_sc_hd__a21oi_2
X_09709_ _11381_/A _09667_/Y _09668_/X _09708_/X vssd1 vssd1 vccd1 vccd1 _09709_/X
+ sky130_fd_sc_hd__a31o_1
X_12720_ _12723_/A hold177/X vssd1 vssd1 vccd1 vccd1 _12721_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_69_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08319__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12651_ _12657_/A _12657_/B _12714_/A _06939_/C vssd1 vssd1 vccd1 vccd1 _12652_/B
+ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_108_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11602_ _11853_/A _11602_/B vssd1 vssd1 vccd1 vccd1 _11606_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12252__B1 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12582_ reg1_val[5] _12583_/B vssd1 vssd1 vccd1 vccd1 _12582_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06781__B _09392_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11533_ _11431_/A _12304_/B _11509_/A _11435_/A vssd1 vssd1 vccd1 vccd1 _11535_/B
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_20_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11464_ _11635_/A _11464_/B vssd1 vssd1 vccd1 vccd1 _11586_/A sky130_fd_sc_hd__xnor2_2
X_13203_ _13309_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_33_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _10415_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10416_/B sky130_fd_sc_hd__or2_1
XFILLER_0_21_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11395_ _06685_/B wire201/X _11838_/A2 _06865_/C _11394_/X vssd1 vssd1 vccd1 vccd1
+ _11395_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_0_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13134_ _13147_/A hold257/X vssd1 vssd1 vccd1 vccd1 _13304_/D sky130_fd_sc_hd__and2_1
XANTENNA__06785__A2 _06778_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10346_ _10346_/A _10346_/B vssd1 vssd1 vccd1 vccd1 _10348_/B sky130_fd_sc_hd__nor2_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ hold272/X _13151_/A2 _13064_/X _12722_/A vssd1 vssd1 vccd1 vccd1 hold273/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12304__A _12786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10277_ _07277_/Y _09295_/B _10433_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _10278_/B
+ sky130_fd_sc_hd__o22a_1
X_12016_ _12205_/A _12203_/A fanout19/X fanout27/X vssd1 vssd1 vccd1 vccd1 _12017_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_0_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13243_/CLK sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12918_ _12946_/A hold196/X vssd1 vssd1 vccd1 vccd1 hold197/A sky130_fd_sc_hd__and2_1
XFILLER_0_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07133__A _07134_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ hold81/X hold276/X vssd1 vssd1 vccd1 vccd1 _13072_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_68_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12243__B1 _12243_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08040_ _08043_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08040_/X sky130_fd_sc_hd__or2_1
XFILLER_0_114_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07670__B1 _07157_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09991_ _09989_/Y _09991_/B vssd1 vssd1 vccd1 vccd1 _09992_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_3_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07973__A1 _12730_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07973__B2 _08819_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08942_ _08942_/A _08942_/B vssd1 vssd1 vccd1 vccd1 _08944_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07308__A _07308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09714__A2 _09710_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_A _13151_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08873_ _08873_/A _08873_/B vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07824_ _08394_/A _07824_/B _07824_/C vssd1 vssd1 vccd1 vccd1 _07825_/C sky130_fd_sc_hd__or3_1
X_07755_ _07754_/A _07754_/B _07754_/C vssd1 vssd1 vccd1 vccd1 _07756_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09478__B2 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09478__A1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06706_ reg2_val[13] _06729_/B vssd1 vssd1 vccd1 vccd1 _06706_/X sky130_fd_sc_hd__and2_1
X_07686_ _07686_/A _08908_/A vssd1 vssd1 vccd1 vccd1 _08940_/A sky130_fd_sc_hd__nand2_2
XANTENNA__07489__B1 _09295_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06637_ reg1_val[23] _07112_/A vssd1 vssd1 vccd1 vccd1 _11922_/A sky130_fd_sc_hd__and2_1
X_09425_ _08681_/A fanout83/X fanout81/X _09295_/A vssd1 vssd1 vccd1 vccd1 _09426_/B
+ sky130_fd_sc_hd__o22a_1
X_06568_ instruction[0] instruction[2] instruction[1] pred_val vssd1 vssd1 vccd1 vccd1
+ _06568_/X sky130_fd_sc_hd__and4bb_1
X_09356_ _09148_/X _09150_/X _09359_/S vssd1 vssd1 vccd1 vccd1 _09356_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08307_ _08308_/B _08308_/C _08394_/A vssd1 vssd1 vccd1 vccd1 _08309_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09287_ _09288_/B _09288_/A vssd1 vssd1 vccd1 vccd1 _09287_/X sky130_fd_sc_hd__and2b_1
X_08238_ _08285_/B _08285_/A vssd1 vssd1 vccd1 vccd1 _08238_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__10260__A2 _09191_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10796__B1 _11347_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11012__B _11147_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08169_ _08169_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _08205_/A sky130_fd_sc_hd__xnor2_2
X_10200_ _10200_/A _10200_/B vssd1 vssd1 vccd1 vccd1 _10201_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_30_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11180_ _11110_/X _11215_/D _12223_/B1 vssd1 vssd1 vccd1 vccd1 _11180_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10131_ _10129_/Y _10131_/B vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__and2b_1
XANTENNA__06767__A2 _06649_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09705__A2 _12250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10062_ _07098_/Y _09295_/B _10433_/A fanout26/X vssd1 vssd1 vccd1 vccd1 _10063_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__06776__B _07279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12703_ reg1_val[29] _12708_/B vssd1 vssd1 vccd1 vccd1 _12704_/B sky130_fd_sc_hd__nand2_1
X_10964_ _09962_/B _10487_/Y _10960_/Y _10961_/Y _10963_/Y vssd1 vssd1 vccd1 vccd1
+ _10965_/B sky130_fd_sc_hd__o311a_2
XFILLER_0_128_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13017__A2 _06537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08692__A2 _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10895_ fanout54/X fanout18/X fanout9/X fanout95/X vssd1 vssd1 vccd1 vccd1 _10896_/B
+ sky130_fd_sc_hd__o22a_1
X_12634_ _12635_/A _12635_/B _12635_/C vssd1 vssd1 vccd1 vccd1 _12639_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_26_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12565_ _12565_/A _12565_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[1] sky130_fd_sc_hd__xor2_4
XFILLER_0_81_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07099__S _10280_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11516_ _11516_/A _11516_/B vssd1 vssd1 vccd1 vccd1 _11529_/A sky130_fd_sc_hd__xnor2_1
X_12496_ reg1_val[18] curr_PC[18] _12524_/S vssd1 vssd1 vccd1 vccd1 _12498_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_80_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11447_ _11358_/A _11357_/B _11355_/X vssd1 vssd1 vccd1 vccd1 _11449_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07404__B1 _12766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ _11317_/X _11730_/B _11377_/Y vssd1 vssd1 vccd1 vccd1 _11378_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09608__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13117_ _13117_/A _13117_/B vssd1 vssd1 vccd1 vccd1 _13117_/Y sky130_fd_sc_hd__xnor2_1
X_10329_ _11429_/A _10329_/B vssd1 vssd1 vccd1 vccd1 _10333_/A sky130_fd_sc_hd__xnor2_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _13048_/A _13048_/B vssd1 vssd1 vccd1 vccd1 _13048_/Y sky130_fd_sc_hd__xnor2_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07183__A2 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09062__B _11183_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07540_ _07541_/A _07541_/B vssd1 vssd1 vccd1 vccd1 _07540_/X sky130_fd_sc_hd__and2_1
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13008__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07471_ _07471_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07472_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_91_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09210_ _10249_/S _09213_/B vssd1 vssd1 vccd1 vccd1 _09211_/B sky130_fd_sc_hd__or2_1
XFILLER_0_8_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11019__A1 _12203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11019__B2 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ reg1_val[14] reg1_val[17] _09172_/S vssd1 vssd1 vccd1 vccd1 _09141_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_16_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09072_ _09072_/A _09072_/B vssd1 vssd1 vccd1 vccd1 _09073_/D sky130_fd_sc_hd__xnor2_4
XFILLER_0_112_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10778__B1 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08023_ _08023_/A _08023_/B vssd1 vssd1 vccd1 vccd1 _08066_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_112_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout207_A _07763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09974_ _09353_/X _09364_/X _10246_/S vssd1 vssd1 vccd1 vccd1 _09974_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08925_ _08925_/A _08925_/B vssd1 vssd1 vccd1 vccd1 _08927_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_99_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08856_ _08217_/B fanout84/X fanout82/X fanout55/X vssd1 vssd1 vccd1 vccd1 _08857_/B
+ sky130_fd_sc_hd__o22a_1
X_07807_ _08772_/B2 fanout94/X _12752_/A _08772_/A2 vssd1 vssd1 vccd1 vccd1 _07808_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12598__B _12598_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06921__A2 _09205_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08787_ _07976_/Y _08658_/B _08656_/X vssd1 vssd1 vccd1 vccd1 _08792_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_79_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07738_ _07738_/A _07738_/B _07738_/C vssd1 vssd1 vccd1 vccd1 _07754_/A sky130_fd_sc_hd__or3_1
XFILLER_0_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07669_ _09467_/A _07669_/B vssd1 vssd1 vccd1 vccd1 _07676_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__09871__A1 _08680_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout22_A _07138_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10680_ fanout77/X _07322_/A _07322_/B fanout62/X fanout46/X vssd1 vssd1 vccd1 vccd1
+ _10681_/B sky130_fd_sc_hd__o32a_1
X_09408_ _10280_/A _09408_/B vssd1 vssd1 vccd1 vccd1 _09412_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__09871__B2 fanout30/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09339_ _08594_/B _12131_/A _09338_/X vssd1 vssd1 vccd1 vccd1 _09339_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09623__B2 fanout77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09623__A1 fanout62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12350_ _12350_/A _12350_/B vssd1 vssd1 vccd1 vccd1 _12352_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11430__B2 _10559_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11301_ _11289_/A _11838_/A2 _11297_/X _11298_/Y _11300_/X vssd1 vssd1 vccd1 vccd1
+ _11301_/X sky130_fd_sc_hd__a221o_1
X_12281_ reg1_val[28] reg1_val[29] _12281_/C vssd1 vssd1 vccd1 vccd1 _12361_/C sky130_fd_sc_hd__and3_1
XFILLER_0_50_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11232_ fanout37/X _11794_/A _11704_/A fanout35/X vssd1 vssd1 vccd1 vccd1 _11233_/B
+ sky130_fd_sc_hd__o22a_1
X_11163_ _11164_/A _11164_/B vssd1 vssd1 vccd1 vccd1 _11217_/B sky130_fd_sc_hd__nand2b_1
X_10114_ _09524_/X _09529_/X _10246_/S vssd1 vssd1 vccd1 vccd1 _10114_/X sky130_fd_sc_hd__mux2_1
X_11094_ hold215/A _11201_/C _11559_/A vssd1 vssd1 vccd1 vccd1 _11095_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__06787__A _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11693__A _12019_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10045_ _10658_/A _10045_/B vssd1 vssd1 vccd1 vccd1 _10049_/A sky130_fd_sc_hd__xnor2_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12301__B fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11996_ _06602_/Y _09194_/Y _10638_/B vssd1 vssd1 vccd1 vccd1 _11996_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08665__A2 _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10947_ _10947_/A _10947_/B vssd1 vssd1 vccd1 vccd1 _10949_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07873__B1 _08692_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12749__A1 _10694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10878_ _09842_/B _10986_/B hold274/A vssd1 vssd1 vccd1 vccd1 _10878_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ _12617_/A _12617_/B _12617_/C vssd1 vssd1 vccd1 vccd1 _12618_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12548_ _12548_/A _12548_/B vssd1 vssd1 vccd1 vccd1 new_PC[25] sky130_fd_sc_hd__xnor2_4
XANTENNA__07130__B _07153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12479_ _12485_/B _12479_/B vssd1 vssd1 vccd1 vccd1 new_PC[14] sky130_fd_sc_hd__and2_4
XANTENNA_2 _07157_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10772__A _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11868__A _12772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13174__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09378__B1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ reg1_val[23] _06971_/B vssd1 vssd1 vccd1 vccd1 _06999_/A sky130_fd_sc_hd__xor2_4
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _07980_/A _07980_/C _07980_/B vssd1 vssd1 vccd1 vccd1 _08712_/B sky130_fd_sc_hd__o21ba_1
X_09690_ _10246_/S _09160_/X _09211_/B vssd1 vssd1 vccd1 vccd1 _09690_/X sky130_fd_sc_hd__o21a_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08641_ _08641_/A _08641_/B vssd1 vssd1 vccd1 vccd1 _08641_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08572_ _09362_/S _08572_/B _08583_/A vssd1 vssd1 vccd1 vccd1 _08572_/X sky130_fd_sc_hd__and3_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12988__A1 _10819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07523_ _07524_/A _07524_/B vssd1 vssd1 vccd1 vccd1 _07523_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07454_ _10155_/A _07454_/B vssd1 vssd1 vccd1 vccd1 _07458_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08408__A2 _09618_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07385_ _07385_/A _07385_/B vssd1 vssd1 vccd1 vccd1 _07694_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09124_ reg1_val[5] reg1_val[26] _09173_/S vssd1 vssd1 vccd1 vccd1 _09124_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11412__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11412__A1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09055_ _09055_/A _09055_/B vssd1 vssd1 vccd1 vccd1 _10859_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08006_ _08007_/A _08007_/B vssd1 vssd1 vccd1 vccd1 _08006_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08041__B1 _07181_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09957_ _09958_/A _09958_/B vssd1 vssd1 vccd1 vccd1 _09957_/X sky130_fd_sc_hd__and2_1
X_08908_ _08908_/A _08908_/B _08908_/C vssd1 vssd1 vccd1 vccd1 _08910_/B sky130_fd_sc_hd__nand3_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _10064_/B2 _07278_/B fanout7/X _09888_/B2 vssd1 vssd1 vccd1 vccd1 _09889_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12140__A2 fanout15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08839_ _08840_/A _08840_/B vssd1 vssd1 vccd1 vccd1 _08899_/A sky130_fd_sc_hd__nand2_1
X_11850_ fanout35/X _12203_/A fanout19/X fanout37/X vssd1 vssd1 vccd1 vccd1 _11851_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09844__A1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08647__A2 _09925_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11781_ _10565_/A _06987_/B fanout9/X _10555_/A vssd1 vssd1 vccd1 vccd1 _11783_/B
+ sky130_fd_sc_hd__o31a_1
X_10801_ _10801_/A _10801_/B vssd1 vssd1 vccd1 vccd1 _10802_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11100__B1 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10732_ _10732_/A _10960_/A vssd1 vssd1 vccd1 vccd1 _10732_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_36_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07231__A _10658_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08046__B _09752_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10663_ _10663_/A _10663_/B vssd1 vssd1 vccd1 vccd1 _10664_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11403__A1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12402_ _12408_/B _12402_/B vssd1 vssd1 vccd1 vccd1 new_PC[3] sky130_fd_sc_hd__and2_4
XFILLER_0_51_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10594_ _10592_/A _10592_/B _10595_/B vssd1 vssd1 vccd1 vccd1 _10594_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12333_ _06631_/A _09383_/B _09191_/X vssd1 vssd1 vccd1 vccd1 _12333_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_35_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11688__A _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12264_ _12264_/A _12264_/B _12264_/C vssd1 vssd1 vccd1 vccd1 _12266_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_120_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12195_ _11381_/A _12174_/X _12182_/X _12194_/X vssd1 vssd1 vccd1 vccd1 _12195_/X
+ sky130_fd_sc_hd__a211o_1
X_11215_ _11215_/A _11215_/B _11215_/C _11215_/D vssd1 vssd1 vccd1 vccd1 _11316_/C
+ sky130_fd_sc_hd__or4_1
XFILLER_0_128_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11146_ _11028_/A _11028_/B _11025_/A vssd1 vssd1 vccd1 vccd1 _11148_/A sky130_fd_sc_hd__a21oi_1
X_11077_ _09059_/A _09059_/B _12131_/A vssd1 vssd1 vccd1 vccd1 _11077_/X sky130_fd_sc_hd__a21o_1
XANTENNA__06948__C _09679_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _10161_/A _10028_/B vssd1 vssd1 vccd1 vccd1 _10030_/C sky130_fd_sc_hd__and2_1
XANTENNA__07125__B _07126_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09621__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11979_ _11906_/A _11904_/X _11922_/A vssd1 vssd1 vccd1 vccd1 _11979_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08237__A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07141__A _08595_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07170_ reg1_val[12] _07170_/B vssd1 vssd1 vccd1 vccd1 _07172_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_54_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08271__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10905__B1 fanout70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout306 instruction[6] vssd1 vssd1 vccd1 vccd1 _09198_/C sky130_fd_sc_hd__buf_2
X_09811_ _09811_/A _09811_/B vssd1 vssd1 vccd1 vccd1 _09814_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07019__C _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ _09742_/A _09742_/B vssd1 vssd1 vccd1 vccd1 _09746_/A sky130_fd_sc_hd__xnor2_1
X_06954_ reg1_val[24] _07087_/B _07087_/C _07165_/A vssd1 vssd1 vccd1 vccd1 _06955_/B
+ sky130_fd_sc_hd__o31a_2
X_06885_ reg1_idx[2] reg1_idx[3] _06885_/C _06885_/D vssd1 vssd1 vccd1 vccd1 int_return
+ sky130_fd_sc_hd__and4_4
XFILLER_0_118_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09673_ _09352_/X _09362_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09673_/X sky130_fd_sc_hd__mux2_1
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _08338_/X _08626_/B _08295_/X vssd1 vssd1 vccd1 vccd1 _08624_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10684__A2 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _08559_/A _08555_/B vssd1 vssd1 vccd1 vccd1 _08568_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_77_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10677__A _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07506_ _07506_/A _07506_/B vssd1 vssd1 vccd1 vccd1 _07527_/A sky130_fd_sc_hd__xnor2_1
X_08486_ _08614_/A vssd1 vssd1 vccd1 vccd1 _08486_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_4_13_0_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _13296_/CLK sky130_fd_sc_hd__clkbuf_8
X_07437_ _08758_/A2 _12786_/A fanout9/X _06864_/A vssd1 vssd1 vccd1 vccd1 _07438_/B
+ sky130_fd_sc_hd__o22a_2
XANTENNA__09677__S _10249_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07368_ _08841_/A1 fanout46/X _11603_/A _08841_/B2 vssd1 vssd1 vccd1 vccd1 _07369_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_33_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09107_ _12131_/A wire3/X vssd1 vssd1 vccd1 vccd1 _09108_/B sky130_fd_sc_hd__or2_1
XFILLER_0_115_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07299_ reg1_val[19] _07299_/B vssd1 vssd1 vccd1 vccd1 _08842_/A sky130_fd_sc_hd__xor2_4
X_09038_ _09668_/B _09668_/C vssd1 vssd1 vccd1 vccd1 _09821_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12897__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07368__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09762__B1 fanout18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11000_ _11000_/A _11316_/A _11215_/A _11215_/B vssd1 vssd1 vccd1 vccd1 _11000_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__12132__A _12133_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12951_ hold165/X _12955_/A2 _13168_/B1 _13246_/Q vssd1 vssd1 vccd1 vccd1 hold166/A
+ sky130_fd_sc_hd__a22o_1
X_12882_ hold68/X hold264/X vssd1 vssd1 vccd1 vccd1 _13148_/B sky130_fd_sc_hd__nand2b_1
X_11902_ _12131_/A _09075_/Y _09076_/Y _11381_/A _11901_/Y vssd1 vssd1 vccd1 vccd1
+ _11902_/X sky130_fd_sc_hd__o311a_1
X_11833_ _12119_/B1 _11989_/C hold293/A vssd1 vssd1 vccd1 vccd1 _11833_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09817__A1 _09511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ curr_PC[21] _11764_/B vssd1 vssd1 vccd1 vccd1 _11929_/C sky130_fd_sc_hd__and2_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11695_ _11695_/A _11695_/B vssd1 vssd1 vccd1 vccd1 _11699_/B sky130_fd_sc_hd__xnor2_1
X_10715_ _10533_/A _10533_/B _10530_/Y vssd1 vssd1 vccd1 vccd1 _10718_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_126_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07896__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10646_ curr_PC[9] curr_PC[10] _10646_/C vssd1 vssd1 vccd1 vccd1 _10887_/C sky130_fd_sc_hd__and3_1
XFILLER_0_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10577_ _10677_/A _08134_/B _10677_/B fanout58/X vssd1 vssd1 vccd1 vccd1 _10578_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13296_ _13296_/CLK _13296_/D vssd1 vssd1 vccd1 vccd1 hold258/A sky130_fd_sc_hd__dfxtp_1
X_12316_ _12316_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12319_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_11_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12247_ _12241_/Y _12242_/X _12246_/Y vssd1 vssd1 vccd1 vccd1 _12247_/X sky130_fd_sc_hd__o21a_1
XANTENNA__07359__A2 _08825_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09753__B1 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12178_ _12176_/Y _12178_/B vssd1 vssd1 vccd1 vccd1 _12179_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11129_ _11129_/A _11129_/B vssd1 vssd1 vccd1 vccd1 _11131_/B sky130_fd_sc_hd__xnor2_1
X_06670_ _06687_/A _12573_/B vssd1 vssd1 vccd1 vccd1 _06670_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_59_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08340_ _08340_/A vssd1 vssd1 vccd1 vccd1 _09061_/A sky130_fd_sc_hd__inv_2
XANTENNA__07819__B1 _11147_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08271_ _10144_/B2 _08774_/B1 _08835_/B1 _08774_/A2 vssd1 vssd1 vccd1 vccd1 _08272_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__10969__A3 _09059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07222_ _07222_/A _07222_/B vssd1 vssd1 vccd1 vccd1 _07379_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07153_ _07153_/A _07153_/B vssd1 vssd1 vccd1 vccd1 _07153_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ _07084_/A vssd1 vssd1 vccd1 vccd1 _07409_/B sky130_fd_sc_hd__inv_2
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout103 _07035_/X vssd1 vssd1 vccd1 vccd1 _10527_/A sky130_fd_sc_hd__buf_8
XANTENNA__08547__A1 _09478_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08547__B2 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout125 _07319_/Y vssd1 vssd1 vccd1 vccd1 _08672_/B sky130_fd_sc_hd__buf_4
Xfanout136 _07057_/X vssd1 vssd1 vccd1 vccd1 _07058_/A sky130_fd_sc_hd__buf_6
Xfanout147 _06952_/Y vssd1 vssd1 vccd1 vccd1 _09772_/A sky130_fd_sc_hd__clkbuf_8
Xfanout114 _10015_/A vssd1 vssd1 vccd1 vccd1 _10555_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07986_ _12768_/A _08692_/A2 _08692_/B1 _12766_/A vssd1 vssd1 vccd1 vccd1 _07987_/B
+ sky130_fd_sc_hd__o22a_2
Xfanout158 _08681_/B vssd1 vssd1 vccd1 vccd1 _12730_/A sky130_fd_sc_hd__buf_6
Xfanout169 _07093_/Y vssd1 vssd1 vccd1 vccd1 _08748_/B1 sky130_fd_sc_hd__buf_6
XANTENNA__07046__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06937_ reg1_val[20] reg1_val[21] reg1_val[22] vssd1 vssd1 vccd1 vccd1 _06940_/B
+ sky130_fd_sc_hd__or3_1
X_09725_ _09725_/A _09725_/B vssd1 vssd1 vccd1 vccd1 _09726_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_96_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09656_ _09656_/A _09656_/B vssd1 vssd1 vccd1 vccd1 _09659_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_97_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06868_ _10108_/A _09970_/A _06868_/C _06868_/D vssd1 vssd1 vccd1 vccd1 _06870_/C
+ sky130_fd_sc_hd__and4bb_1
X_08607_ _08609_/A _08609_/B _09047_/A vssd1 vssd1 vccd1 vccd1 _09049_/B sky130_fd_sc_hd__a21o_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07522__A2 _12349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06799_ _06986_/A reg1_val[7] vssd1 vssd1 vccd1 vccd1 _06799_/X sky130_fd_sc_hd__and2b_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ _09588_/A _09588_/B vssd1 vssd1 vccd1 vccd1 _09736_/B sky130_fd_sc_hd__nor2_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _08538_/A _08538_/B vssd1 vssd1 vccd1 vccd1 _08609_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_49_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10409__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08469_ _08589_/A _08469_/B vssd1 vssd1 vccd1 vccd1 _08492_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07286__A1 _07179_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07286__B2 fanout54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10500_ _10392_/A _10389_/Y _10391_/B vssd1 vssd1 vccd1 vccd1 _10504_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_52_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11480_ hold178/A hold207/A _11480_/C vssd1 vssd1 vccd1 vccd1 _11573_/B sky130_fd_sc_hd__or3_1
XFILLER_0_80_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10431_ _10432_/A _10432_/B vssd1 vssd1 vccd1 vccd1 _10586_/B sky130_fd_sc_hd__nand2b_1
X_13150_ hold264/A _13149_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13150_/X sky130_fd_sc_hd__mux2_1
X_10362_ _10609_/B _10609_/C vssd1 vssd1 vccd1 vccd1 _10362_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10042__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13081_ _13086_/A hold275/X vssd1 vssd1 vccd1 vccd1 _13293_/D sky130_fd_sc_hd__and2_1
X_12101_ _12101_/A _12101_/B _12163_/A vssd1 vssd1 vccd1 vccd1 _12101_/X sky130_fd_sc_hd__and3_1
X_10293_ _10435_/A _10293_/B vssd1 vssd1 vccd1 vccd1 _10295_/B sky130_fd_sc_hd__nand2_1
X_12032_ _12032_/A _12032_/B _12032_/C vssd1 vssd1 vccd1 vccd1 _12033_/B sky130_fd_sc_hd__nand3_1
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
X_12934_ _12946_/A hold235/X vssd1 vssd1 vccd1 vccd1 hold236/A sky130_fd_sc_hd__and2_1
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07513__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12865_ _13112_/A _13113_/A _13112_/B vssd1 vssd1 vccd1 vccd1 _13117_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12796_ hold79/X hold286/A vssd1 vssd1 vccd1 vccd1 _12796_/X sky130_fd_sc_hd__and2b_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11816_ _11967_/A _11816_/B vssd1 vssd1 vccd1 vccd1 _11972_/C sky130_fd_sc_hd__xnor2_2
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11747_ _11746_/A _10642_/Y _11746_/Y _09205_/B vssd1 vssd1 vccd1 vccd1 _11747_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_56_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07122__C _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10820__A2 _07435_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11678_ _12022_/A _11678_/B vssd1 vssd1 vccd1 vccd1 _11680_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10629_ _09971_/Y _10628_/Y _10752_/S vssd1 vssd1 vccd1 vccd1 _10629_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11781__B1 _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13279_ _13280_/CLK hold50/X vssd1 vssd1 vccd1 vccd1 hold296/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12325__A2 _12279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09065__B _11379_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _07840_/A _07840_/B vssd1 vssd1 vccd1 vccd1 _07841_/B sky130_fd_sc_hd__xor2_2
XANTENNA__07201__B2 _10452_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07201__A1 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ _08420_/B fanout82/X _09295_/B _08854_/B2 vssd1 vssd1 vccd1 vccd1 _07772_/B
+ sky130_fd_sc_hd__o22a_1
X_06722_ _06722_/A _06722_/B vssd1 vssd1 vccd1 vccd1 _06866_/A sky130_fd_sc_hd__or2_1
X_09510_ _09100_/B wire5/X _09508_/Y wire4/X vssd1 vssd1 vccd1 vccd1 _09511_/B sky130_fd_sc_hd__a211oi_4
XFILLER_0_79_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06653_ reg1_val[20] _06653_/B vssd1 vssd1 vccd1 vccd1 _06654_/B sky130_fd_sc_hd__or2_1
XFILLER_0_78_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09441_ _09442_/A _09442_/B vssd1 vssd1 vccd1 vccd1 _09575_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09372_ _12563_/A curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09373_/B sky130_fd_sc_hd__and2_1
X_06584_ reg1_val[29] _07243_/A vssd1 vssd1 vccd1 vccd1 _06585_/B sky130_fd_sc_hd__nand2b_1
X_08323_ _09888_/B2 _08772_/B2 _08772_/A2 _07969_/A vssd1 vssd1 vccd1 vccd1 _08324_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__08465__B1 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07268__B2 fanout57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07268__A1 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09662__C1 _09816_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08254_ _08294_/A _08294_/B _08214_/Y vssd1 vssd1 vccd1 vccd1 _08259_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_117_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08185_ _08244_/A _08195_/B vssd1 vssd1 vccd1 vccd1 _08185_/X sky130_fd_sc_hd__or2_1
XFILLER_0_105_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07205_ _07205_/A _07205_/B vssd1 vssd1 vccd1 vccd1 _07209_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_40_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07136_ _07153_/A _07129_/B _07129_/C _07129_/D _07434_/A vssd1 vssd1 vccd1 vccd1
+ _07136_/X sky130_fd_sc_hd__o41a_1
XANTENNA__10024__B1 fanout14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07067_ _07303_/B _07129_/B _06653_/B vssd1 vssd1 vccd1 vccd1 _07821_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_70_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10575__A1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10575__B2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10690__A _12255_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06599__B _06633_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07991__A2 _08774_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07969_ _07969_/A _09752_/B vssd1 vssd1 vccd1 vccd1 _07971_/B sky130_fd_sc_hd__or2_1
X_09708_ _09183_/Y _09682_/X _12235_/B _09158_/S _09707_/X vssd1 vssd1 vccd1 vccd1
+ _09708_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_4_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10980_ _11194_/S _09974_/X _10979_/X _10752_/S vssd1 vssd1 vccd1 vccd1 _10980_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_fanout52_A _08134_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09639_ _09640_/A _09640_/B vssd1 vssd1 vccd1 vccd1 _09641_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07504__A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12650_ _12648_/X _12650_/B vssd1 vssd1 vccd1 vccd1 _12657_/C sky130_fd_sc_hd__nand2b_2
XFILLER_0_93_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12252__A1 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11601_ fanout33/X fanout19/X _12301_/A _10553_/A vssd1 vssd1 vccd1 vccd1 _11602_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12556__S _12556_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12252__B2 _12301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12581_ _12580_/A _12577_/Y _12579_/B vssd1 vssd1 vccd1 vccd1 _12585_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_108_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11532_ _11532_/A _11532_/B vssd1 vssd1 vccd1 vccd1 _11535_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11463_ _11073_/B _11462_/Y _11461_/Y vssd1 vssd1 vccd1 vccd1 _11464_/B sky130_fd_sc_hd__a21o_1
X_13202_ _13309_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ _10415_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10416_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13133_ hold256/X _13165_/A2 _13132_/X _13146_/B2 vssd1 vssd1 vccd1 vccd1 hold257/A
+ sky130_fd_sc_hd__a22o_1
X_11394_ _06684_/B _06928_/X _09197_/B _06683_/X _11393_/Y vssd1 vssd1 vccd1 vccd1
+ _11394_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10345_ _10175_/A _10175_/B _10173_/X vssd1 vssd1 vccd1 vccd1 _10348_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_21_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13064_ hold268/X _13063_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _13064_/X sky130_fd_sc_hd__mux2_1
XANTENNA__12304__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10276_ _10218_/A _10218_/B _10219_/Y vssd1 vssd1 vccd1 vccd1 _10357_/A sky130_fd_sc_hd__o21ai_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10105__A _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ _11935_/A _12304_/B _12011_/A _11939_/A vssd1 vssd1 vccd1 vccd1 _12027_/A
+ sky130_fd_sc_hd__o31ai_2
X_12917_ hold219/A _12947_/A2 _12947_/B1 hold195/X vssd1 vssd1 vccd1 vccd1 hold196/A
+ sky130_fd_sc_hd__a22o_1
X_12848_ _13067_/A _13068_/A _13067_/B vssd1 vssd1 vccd1 vccd1 _13073_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_61_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07133__B _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12779_ _12087_/A _12781_/A2 hold80/X _13147_/A vssd1 vssd1 vccd1 vccd1 _13211_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10254__B1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07670__A1 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07670__B2 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09990_ reg1_val[5] curr_PC[5] vssd1 vssd1 vccd1 vccd1 _09991_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07973__A2 _07322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08941_ _08941_/A _08941_/B vssd1 vssd1 vccd1 vccd1 _08944_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11506__B1 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08872_ _08872_/A _08872_/B vssd1 vssd1 vccd1 vccd1 _08873_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__07308__B _07308_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07823_ _07824_/B _07824_/C _08394_/A vssd1 vssd1 vccd1 vccd1 _07825_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__10015__A _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout187_A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07754_ _07754_/A _07754_/B _07754_/C vssd1 vssd1 vccd1 vccd1 _07756_/A sky130_fd_sc_hd__and3_1
XANTENNA__12230__A _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09478__A2 _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06705_ _06705_/A vssd1 vssd1 vccd1 vccd1 _06867_/B sky130_fd_sc_hd__inv_2
XFILLER_0_79_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07685_ _07686_/A _08813_/A _07685_/C vssd1 vssd1 vccd1 vccd1 _08908_/A sky130_fd_sc_hd__nand3_2
XANTENNA__07489__B2 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07489__A1 fanout81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06636_ _06634_/Y _06680_/B1 _06729_/B reg2_val[23] vssd1 vssd1 vccd1 vccd1 _07112_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_35_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09424_ _09580_/A _09424_/B vssd1 vssd1 vccd1 vccd1 _09428_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_87_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06700__A3 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09355_ _09347_/X _09354_/X _10750_/S vssd1 vssd1 vccd1 vccd1 _09355_/X sky130_fd_sc_hd__mux2_1
X_06567_ _09198_/B _06567_/B vssd1 vssd1 vccd1 vccd1 is_store sky130_fd_sc_hd__nor2_8
XANTENNA__10685__A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08306_ _07313_/A _07313_/B _08758_/A2 vssd1 vssd1 vccd1 vccd1 _08308_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10796__A1 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09286_ _12349_/B _09286_/B vssd1 vssd1 vccd1 vccd1 _09288_/B sky130_fd_sc_hd__xnor2_2
X_08237_ _09452_/A _08237_/B vssd1 vssd1 vccd1 vccd1 _08285_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10796__B2 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08168_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08168_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08099_ _08099_/A _08099_/B vssd1 vssd1 vccd1 vccd1 _08154_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12405__A _12578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07119_ _07119_/A _07119_/B vssd1 vssd1 vccd1 vccd1 _07119_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10130_ reg1_val[6] curr_PC[6] vssd1 vssd1 vccd1 vccd1 _10131_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06767__A3 _12578_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10061_ _10061_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _10072_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10963_ _10729_/Y _11174_/A _10962_/Y vssd1 vssd1 vccd1 vccd1 _10963_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12702_ reg1_val[29] _12708_/B vssd1 vssd1 vccd1 vccd1 _12704_/A sky130_fd_sc_hd__or2_1
XFILLER_0_128_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_730 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10894_ _10894_/A _10894_/B vssd1 vssd1 vccd1 vccd1 _10898_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12633_ _12639_/A _12633_/B vssd1 vssd1 vccd1 vccd1 _12635_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10236__B1 _09110_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12564_ _12564_/A _12564_/B vssd1 vssd1 vccd1 vccd1 _12565_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_65_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11515_ _11516_/A _11516_/B vssd1 vssd1 vccd1 vccd1 _11515_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_19_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12495_ _12500_/B _12495_/B vssd1 vssd1 vccd1 vccd1 new_PC[17] sky130_fd_sc_hd__xnor2_4
XFILLER_0_53_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ _11446_/A _11446_/B vssd1 vssd1 vccd1 vccd1 _11449_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07404__B2 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07404__A1 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11377_ _11317_/X _11730_/B _12223_/B1 vssd1 vssd1 vccd1 vccd1 _11377_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13116_ _13116_/A hold281/X vssd1 vssd1 vccd1 vccd1 _13300_/D sky130_fd_sc_hd__and2_1
X_10328_ _12774_/A fanout52/X _10677_/B _12772_/A vssd1 vssd1 vccd1 vccd1 _10329_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13047_/A _13047_/B vssd1 vssd1 vccd1 vccd1 _13048_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09157__A1 _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _06744_/B _12243_/B1 _10257_/Y _10258_/X vssd1 vssd1 vccd1 vccd1 _10259_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__09624__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09062__C _11285_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08668__B1 _10694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07340__B1 _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07470_ _07471_/A _07471_/B vssd1 vssd1 vccd1 vccd1 _07472_/A sky130_fd_sc_hd__or2_1
XFILLER_0_118_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11019__A2 _10557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09140_ _09138_/X _09139_/X _09359_/S vssd1 vssd1 vccd1 vccd1 _09140_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_127_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09071_ _09022_/A _09023_/Y _09070_/Y _09063_/B _09025_/X vssd1 vssd1 vccd1 vccd1
+ _09072_/B sky130_fd_sc_hd__o221a_2
XFILLER_0_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10778__A1 fanout27/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10778__B2 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08022_ _08023_/A _08023_/B vssd1 vssd1 vccd1 vccd1 _08022_/X sky130_fd_sc_hd__and2_1
XFILLER_0_112_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout102_A _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09973_ _09346_/X _09350_/X _10247_/S vssd1 vssd1 vccd1 vccd1 _09973_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08924_ _08873_/A _08873_/B _08871_/X vssd1 vssd1 vccd1 vccd1 _08925_/B sky130_fd_sc_hd__a21oi_4
X_08855_ _08855_/A _08855_/B vssd1 vssd1 vccd1 vccd1 _08859_/A sky130_fd_sc_hd__xnor2_1
X_07806_ _08855_/A _07806_/B vssd1 vssd1 vccd1 vccd1 _07809_/A sky130_fd_sc_hd__xnor2_2
X_08786_ _08703_/A _08703_/C _08703_/B vssd1 vssd1 vccd1 vccd1 _08796_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__09253__B _12087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07737_ _07737_/A _07737_/B vssd1 vssd1 vccd1 vccd1 _07738_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__08659__B1 fanout51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ fanout77/X _09618_/B2 _09618_/A1 _12768_/A vssd1 vssd1 vccd1 vccd1 _07669_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07331__B1 fanout33/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09871__A2 _07197_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06619_ _06619_/A _06619_/B vssd1 vssd1 vccd1 vccd1 _06620_/B sky130_fd_sc_hd__nand2_2
X_09407_ _09888_/B2 _07389_/B fanout26/X _12736_/A vssd1 vssd1 vccd1 vccd1 _09408_/B
+ sky130_fd_sc_hd__o22a_1
X_07599_ _07599_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07601_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09338_ reg1_val[0] _09362_/S _09283_/A _09620_/A _09337_/X vssd1 vssd1 vccd1 vccd1
+ _09338_/X sky130_fd_sc_hd__a41o_1
XFILLER_0_124_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10769__A1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout15_A _07278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09623__A2 fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11300_ _06693_/B wire201/X _09197_/B _06691_/Y _11299_/X vssd1 vssd1 vccd1 vccd1
+ _11300_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09269_ _10184_/A _09269_/B vssd1 vssd1 vccd1 vccd1 _09271_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12280_ _12279_/A _12279_/B _12279_/Y _11184_/A vssd1 vssd1 vccd1 vccd1 _12280_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_31_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09387__A1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11231_ _11354_/A _11231_/B vssd1 vssd1 vccd1 vccd1 _11235_/B sky130_fd_sc_hd__or2_1
XFILLER_0_15_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11162_ _11162_/A _11162_/B vssd1 vssd1 vccd1 vccd1 _11164_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__07229__A _09610_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ _10246_/S _09521_/X _10112_/X _11089_/A vssd1 vssd1 vccd1 vccd1 _10113_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__06987__C_N _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11093_ _11088_/Y _11092_/A _11197_/S vssd1 vssd1 vccd1 vccd1 _11093_/X sky130_fd_sc_hd__mux2_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
X_10044_ _10452_/B2 _12782_/A fanout22/X _10527_/A vssd1 vssd1 vccd1 vccd1 _10045_/B
+ sky130_fd_sc_hd__o22a_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06787__B _09679_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
X_11995_ _11995_/A _11995_/B vssd1 vssd1 vccd1 vccd1 _12000_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10946_ _10834_/A _10833_/B _10831_/Y vssd1 vssd1 vccd1 vccd1 _10947_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_128_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10877_ hold291/A _10877_/B vssd1 vssd1 vccd1 vccd1 _10986_/B sky130_fd_sc_hd__or2_1
XANTENNA__07873__A1 _12760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07873__B2 _09925_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12749__A2 _12980_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12616_ _12617_/A _12617_/B _12617_/C vssd1 vssd1 vccd1 vccd1 _12623_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_115_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12547_ _12557_/A _12538_/B _12542_/A _12542_/B vssd1 vssd1 vccd1 vccd1 _12548_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_108_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12478_ _12478_/A _12478_/B _12478_/C vssd1 vssd1 vccd1 vccd1 _12479_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12126__A2_N _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09619__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_3 _12786_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11868__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13174__A2 _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11429_ _11429_/A _11429_/B fanout9/X vssd1 vssd1 vccd1 vccd1 _11429_/X sky130_fd_sc_hd__or3_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12382__A0 _12563_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ _07087_/B _06940_/B _12658_/B _07165_/A vssd1 vssd1 vccd1 vccd1 _06971_/B
+ sky130_fd_sc_hd__o31a_2
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11488__A2 _09188_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08640_ _08641_/A _08641_/B vssd1 vssd1 vccd1 vccd1 _09074_/B sky130_fd_sc_hd__xor2_4
XANTENNA__06697__B _07178_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09073__B _11559_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__B2 _09201_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11823__S _11823_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08571_ _09362_/S _08572_/B vssd1 vssd1 vccd1 vccd1 _08583_/B sky130_fd_sc_hd__nand2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12988__A2 _13020_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07522_ _06864_/A _12349_/A _08595_/A vssd1 vssd1 vccd1 vccd1 _07524_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__10999__A1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11660__A2 _11838_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09853__A2 _09383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07453_ _07058_/A _10557_/A fanout58/X _08532_/B vssd1 vssd1 vccd1 vccd1 _07454_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_91_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11124__A _11125_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07384_ _07384_/A _07384_/B vssd1 vssd1 vccd1 vccd1 _07694_/A sky130_fd_sc_hd__nor2_1
X_09123_ reg1_val[4] reg1_val[27] _09173_/S vssd1 vssd1 vccd1 vccd1 _09123_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11412__A2 _11935_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09054_ _09054_/A _09054_/B vssd1 vssd1 vccd1 vccd1 _10740_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_32_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13165__A2 _13165_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08005_ _08004_/B _07753_/B _08004_/Y vssd1 vssd1 vccd1 vccd1 _08007_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08041__A1 _08837_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12373__B1 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap250 _09620_/A vssd1 vssd1 vccd1 vccd1 _08394_/A sky130_fd_sc_hd__buf_6
XFILLER_0_4_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08041__B2 _07969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12125__B1 _10638_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11794__A _11794_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ _09958_/A _09958_/B vssd1 vssd1 vccd1 vccd1 _09956_/X sky130_fd_sc_hd__or2_1
X_08907_ _08907_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08908_/C sky130_fd_sc_hd__and2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ _09887_/A _09887_/B vssd1 vssd1 vccd1 vccd1 _09891_/A sky130_fd_sc_hd__xor2_1
X_08838_ _10565_/A _08838_/B vssd1 vssd1 vccd1 vccd1 _08840_/B sky130_fd_sc_hd__xnor2_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10203__A _11695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ _08768_/A _08768_/B _08768_/C vssd1 vssd1 vccd1 vccd1 _08770_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__11100__A1 _07192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11780_ _11780_/A _11780_/B vssd1 vssd1 vccd1 vccd1 _11783_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__10439__B1 _11603_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ _10801_/A _10801_/B vssd1 vssd1 vccd1 vccd1 _10802_/A sky130_fd_sc_hd__and2_1
XFILLER_0_95_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10731_ _10488_/Y _10960_/A _10729_/Y vssd1 vssd1 vccd1 vccd1 _10734_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_55_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ _12401_/A _12401_/B _12401_/C vssd1 vssd1 vccd1 vccd1 _12402_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_36_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10662_ _10662_/A _10662_/B _10662_/C vssd1 vssd1 vccd1 vccd1 _10663_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_106_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10593_ _10463_/A _10463_/B _10462_/A vssd1 vssd1 vccd1 vccd1 _10595_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_23_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12332_ hold231/A _12332_/B _12332_/C vssd1 vssd1 vccd1 vccd1 _12332_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_51_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11688__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12263_ _12263_/A _12263_/B vssd1 vssd1 vccd1 vccd1 _12264_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11214_ _12556_/S _11212_/Y _11314_/C _11211_/X vssd1 vssd1 vccd1 vccd1 dest_val[15]
+ sky130_fd_sc_hd__o31ai_4
X_12194_ _12194_/A _12194_/B _12185_/X vssd1 vssd1 vccd1 vccd1 _12194_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_31_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11145_ _11143_/Y _11145_/B vssd1 vssd1 vccd1 vccd1 _11152_/A sky130_fd_sc_hd__nand2b_1
X_11076_ _11076_/A _11076_/B vssd1 vssd1 vccd1 vccd1 _11076_/X sky130_fd_sc_hd__or2_4
X_10027_ _10027_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10028_/B sky130_fd_sc_hd__or2_1
XANTENNA__06948__D _08588_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__B1 _12736_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06751__D1 _06898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09902__A _10894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11978_ _11977_/A _11977_/B _11977_/Y _11381_/A vssd1 vssd1 vccd1 vccd1 _11978_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08518__A _10155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10929_ _10930_/A _10930_/B vssd1 vssd1 vccd1 vccd1 _10929_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08271__A1 _10144_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08271__B2 _08774_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12355__B1 _09968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10905__A1 fanout35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__B2 fanout37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09810_ _09810_/A _09810_/B vssd1 vssd1 vccd1 vccd1 _09811_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_10_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07019__D _07303_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06953_ _07087_/B _07087_/C _07165_/A vssd1 vssd1 vccd1 vccd1 _06997_/B sky130_fd_sc_hd__o21ai_2
X_09741_ _10557_/A fanout98/X fanout56/X fanout62/X vssd1 vssd1 vccd1 vccd1 _09742_/B
+ sky130_fd_sc_hd__o22a_1
X_06884_ reg1_idx[5] _06898_/C vssd1 vssd1 vccd1 vccd1 _06885_/D sky130_fd_sc_hd__and2_1
XFILLER_0_118_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10133__A2 _09851_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09672_ _09349_/X _09351_/X _09678_/S vssd1 vssd1 vccd1 vccd1 _09672_/X sky130_fd_sc_hd__mux2_1
XANTENNA__10023__A _10180_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08623_ _08295_/A _08295_/B _08295_/C vssd1 vssd1 vccd1 vccd1 _08626_/B sky130_fd_sc_hd__a21o_1
XANTENNA_fanout267_A _12955_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _08542_/Y _08551_/X _08552_/X _08538_/B vssd1 vssd1 vccd1 vccd1 _08608_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07332__A _10015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10677__B _10677_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07505_ _07506_/B vssd1 vssd1 vccd1 vccd1 _07505_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_92_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08485_ _08485_/A _08485_/B _08485_/C vssd1 vssd1 vccd1 vccd1 _08614_/A sky130_fd_sc_hd__or3_1
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07436_ _09968_/A _07434_/X _06622_/X vssd1 vssd1 vccd1 vccd1 fanout9/A sky130_fd_sc_hd__a21o_1
XFILLER_0_18_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07367_ _11429_/A _07367_/B vssd1 vssd1 vccd1 vccd1 _07371_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11789__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10693__A _10694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ _12278_/B _12279_/A _12326_/A _12360_/A vssd1 vssd1 vccd1 vccd1 wire3/A sky130_fd_sc_hd__nor4_1
XFILLER_0_33_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09037_ _09037_/A _09037_/B vssd1 vssd1 vccd1 vccd1 _09668_/C sky130_fd_sc_hd__xor2_1
X_07298_ reg1_val[18] _07087_/B _06939_/C _07165_/A vssd1 vssd1 vccd1 vccd1 _07299_/B
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_103_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09762__A1 _07058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09762__B2 _08532_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout82_A _07312_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__B1 _11012_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ _09939_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09940_/B sky130_fd_sc_hd__nand2_2
X_12950_ _13169_/A hold214/X vssd1 vssd1 vccd1 vccd1 _13245_/D sky130_fd_sc_hd__and2_1
X_12881_ _12798_/B _13144_/B _12796_/X vssd1 vssd1 vccd1 vccd1 _13149_/A sky130_fd_sc_hd__a21o_1
X_11901_ _12131_/A _09075_/Y _09076_/Y vssd1 vssd1 vccd1 vccd1 _11901_/Y sky130_fd_sc_hd__o21ai_1
X_11832_ hold252/A _11832_/B vssd1 vssd1 vccd1 vccd1 _11989_/C sky130_fd_sc_hd__or2_1
XFILLER_0_68_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11763_ curr_PC[21] _11764_/B vssd1 vssd1 vccd1 vccd1 _11765_/B sky130_fd_sc_hd__nor2_1
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11694_ _11695_/A _11695_/B vssd1 vssd1 vccd1 vccd1 _11791_/A sky130_fd_sc_hd__and2_1
X_10714_ _10588_/A _10588_/B _10587_/A vssd1 vssd1 vccd1 vccd1 _10719_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_126_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10645_ _10614_/Y _10615_/X _10618_/Y _11184_/A _10644_/X vssd1 vssd1 vccd1 vccd1
+ _10645_/X sky130_fd_sc_hd__o221a_2
XFILLER_0_36_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08073__A _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12315_ _12105_/B _12313_/Y _12314_/Y _12266_/B vssd1 vssd1 vccd1 vccd1 _12316_/B
+ sky130_fd_sc_hd__a211o_1
X_10576_ _10894_/A _10576_/B vssd1 vssd1 vccd1 vccd1 _10580_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13295_ _13296_/CLK _13295_/D vssd1 vssd1 vccd1 vccd1 hold282/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12246_ _09158_/S _09682_/X _12245_/X vssd1 vssd1 vccd1 vccd1 _12246_/Y sky130_fd_sc_hd__a21oi_2
X_12177_ reg1_val[27] curr_PC[27] vssd1 vssd1 vccd1 vccd1 _12178_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09753__A1 _07308_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10899__B1 _12205_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07764__B1 _12768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06811__A_N _07197_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ _11429_/A _11128_/B vssd1 vssd1 vccd1 vccd1 _11129_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11312__A1 _10400_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059_ _11060_/A _11060_/B vssd1 vssd1 vccd1 vccd1 _11167_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__13065__B2 _12722_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07152__A _07153_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07819__A1 _08572_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08270_ _10819_/A _08329_/A vssd1 vssd1 vccd1 vccd1 _08270_/X sky130_fd_sc_hd__and2_1
XFILLER_0_104_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06991__A _10555_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07221_ _07221_/A _07221_/B vssd1 vssd1 vccd1 vccd1 _07222_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_13_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09079__A _09079_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07152_ _07153_/A _07153_/B vssd1 vssd1 vccd1 vccd1 _12087_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_13_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11305__A1_N _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ _10458_/A _07083_/B vssd1 vssd1 vccd1 vccd1 _07084_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08547__A2 _08588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout104 _12760_/A vssd1 vssd1 vccd1 vccd1 _11347_/A sky130_fd_sc_hd__buf_6
XFILLER_0_10_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout137 _07057_/X vssd1 vssd1 vccd1 vccd1 _08772_/A2 sky130_fd_sc_hd__buf_4
Xfanout115 _06999_/A vssd1 vssd1 vccd1 vccd1 _10015_/A sky130_fd_sc_hd__buf_8
XANTENNA__07327__A _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout126 _10184_/A vssd1 vssd1 vccd1 vccd1 _11125_/A sky130_fd_sc_hd__buf_12
XFILLER_0_1_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07985_ _07737_/A _07737_/B _07733_/X vssd1 vssd1 vccd1 vccd1 _07997_/A sky130_fd_sc_hd__o21a_2
Xfanout159 _08681_/B vssd1 vssd1 vccd1 vccd1 _09476_/A sky130_fd_sc_hd__clkbuf_8
Xfanout148 _11973_/A vssd1 vssd1 vccd1 vccd1 _10617_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__07046__B _07046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06936_ reg1_val[13] reg1_val[14] reg1_val[15] _07165_/B vssd1 vssd1 vccd1 vccd1
+ _07087_/B sky130_fd_sc_hd__or4_4
XFILLER_0_38_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09724_ _09725_/A _09725_/B vssd1 vssd1 vccd1 vccd1 _09726_/A sky130_fd_sc_hd__or2_1
XANTENNA__07507__B1 fanout56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06867_ _11187_/A _06867_/B _10972_/A _10863_/A vssd1 vssd1 vccd1 vccd1 _06871_/B
+ sky130_fd_sc_hd__and4_1
X_09655_ _09655_/A _09655_/B vssd1 vssd1 vccd1 vccd1 _09656_/B sky130_fd_sc_hd__xor2_4
XANTENNA__08180__B1 fanout84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10511__C1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _08608_/B _09045_/A _08553_/X vssd1 vssd1 vccd1 vccd1 _09047_/A sky130_fd_sc_hd__a21o_1
X_06798_ _10108_/A _06796_/X _06797_/Y vssd1 vssd1 vccd1 vccd1 _06798_/Y sky130_fd_sc_hd__o21ai_1
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09586_ _11695_/A _09586_/B vssd1 vssd1 vccd1 vccd1 _09588_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _08538_/A _08537_/B _08537_/C vssd1 vssd1 vccd1 vccd1 _08538_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_37_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08468_ _08837_/B2 _08588_/B _09273_/A1 _07969_/A vssd1 vssd1 vccd1 vccd1 _08469_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__07286__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07419_ _07417_/A _07417_/B _07418_/Y vssd1 vssd1 vccd1 vccd1 _07426_/B sky130_fd_sc_hd__o21a_2
XANTENNA__10290__A1 _10458_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08399_ _08399_/A _08399_/B vssd1 vssd1 vccd1 vccd1 _08407_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10627__S _11194_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ _10586_/A _10430_/B vssd1 vssd1 vccd1 vccd1 _10432_/B sky130_fd_sc_hd__and2_1
XFILLER_0_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10042__A1 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10042__B2 fanout58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10361_ _10361_/A _10486_/A vssd1 vssd1 vccd1 vccd1 _10609_/C sky130_fd_sc_hd__nor2_1
X_13080_ hold274/X _12721_/B _13079_/X _12722_/A vssd1 vssd1 vccd1 vccd1 hold275/A
+ sky130_fd_sc_hd__a22o_1
X_12100_ _12101_/A _12035_/A _12102_/C vssd1 vssd1 vccd1 vccd1 _12100_/Y sky130_fd_sc_hd__a21oi_1
X_10292_ _10292_/A _10292_/B vssd1 vssd1 vccd1 vccd1 _10293_/B sky130_fd_sc_hd__nand2_1
Xhold180 hold180/A vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
X_12031_ _12032_/A _12032_/B _12032_/C vssd1 vssd1 vccd1 vccd1 _12098_/B sky130_fd_sc_hd__a21o_1
Xhold191 hold191/A vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12143__A _12143_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12933_ _13236_/Q _13146_/B2 _13168_/B1 hold234/X vssd1 vssd1 vccd1 vccd1 hold235/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__09452__A _09452_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12864_ hold88/X hold289/A vssd1 vssd1 vccd1 vccd1 _13112_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12795_ hold264/X hold68/X vssd1 vssd1 vccd1 vccd1 _13148_/A sky130_fd_sc_hd__nand2b_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11815_ _11464_/B _11814_/Y _11813_/Y vssd1 vssd1 vccd1 vccd1 _11816_/B sky130_fd_sc_hd__a21o_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11746_ _11746_/A _11746_/B vssd1 vssd1 vccd1 vccd1 _11746_/Y sky130_fd_sc_hd__nor2_1
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11677_ fanout37/X _12150_/A _12150_/B fanout35/X vssd1 vssd1 vccd1 vccd1 _11678_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11222__A _11222_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10628_ _10628_/A vssd1 vssd1 vccd1 vccd1 _10628_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09423__B1 fanout13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10559_ _10559_/A _10559_/B _10559_/C vssd1 vssd1 vccd1 vccd1 _10562_/C sky130_fd_sc_hd__and3_1
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_251 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13278_ _13280_/CLK _13278_/D vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11781__A1 _10565_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12229_ _06605_/B _12227_/X _12228_/Y vssd1 vssd1 vccd1 vccd1 _12229_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_20_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11533__A1 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09065__C _11468_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07147__A _09621_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07201__A2 _10527_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ _07770_/A _07770_/B vssd1 vssd1 vccd1 vccd1 _07780_/A sky130_fd_sc_hd__xnor2_4
X_06721_ _06722_/A _06722_/B vssd1 vssd1 vccd1 vccd1 _10743_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_79_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09440_ _09258_/B _09261_/B _09258_/A vssd1 vssd1 vccd1 vccd1 _09442_/B sky130_fd_sc_hd__o21bai_2
XANTENNA__06712__A1 _06898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06652_ reg1_val[20] _06653_/B vssd1 vssd1 vccd1 vccd1 _06654_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10301__A _10301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09371_ _12563_/A curr_PC[1] vssd1 vssd1 vccd1 vccd1 _09373_/A sky130_fd_sc_hd__nor2_1
X_06583_ _07243_/A reg1_val[29] vssd1 vssd1 vccd1 vccd1 _06583_/X sky130_fd_sc_hd__and2b_1
X_08322_ _08334_/B _08334_/A vssd1 vssd1 vccd1 vccd1 _08336_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__08465__A1 _06864_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09111__C1 _12223_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07268__A2 fanout95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08253_ _08253_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _08294_/B sky130_fd_sc_hd__xor2_1
XANTENNA__06681__A2_N _06680_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08465__B2 _08758_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10272__A1 _12005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout132_A _10156_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07204_ _09610_/A _07204_/B vssd1 vssd1 vccd1 vccd1 _07205_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_755 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08184_ _08182_/Y _08245_/B _08179_/Y vssd1 vssd1 vccd1 vccd1 _08195_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__09414__B1 _10064_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07135_ _07434_/A _07135_/B vssd1 vssd1 vccd1 vccd1 _07139_/A sky130_fd_sc_hd__nand2_2
XANTENNA__10024__A1 _10553_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10024__B2 fanout69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07066_ _07066_/A _07066_/B vssd1 vssd1 vccd1 vccd1 _07409_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11786__B _11786_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10575__A2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10980__C1 _10752_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07968_ _07968_/A _07968_/B vssd1 vssd1 vccd1 vccd1 _07978_/A sky130_fd_sc_hd__xnor2_1
X_09707_ _09707_/A _09707_/B _09707_/C _09706_/X vssd1 vssd1 vccd1 vccd1 _09707_/X
+ sky130_fd_sc_hd__or4b_1
X_06919_ _09198_/C instruction[4] _09198_/B _09200_/B vssd1 vssd1 vccd1 vccd1 _06919_/X
+ sky130_fd_sc_hd__and4b_1
X_07899_ _08772_/B2 fanout84/X fanout82/X _08772_/A2 vssd1 vssd1 vccd1 vccd1 _07900_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09638_ _09638_/A _09638_/B vssd1 vssd1 vccd1 vccd1 _09640_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_38_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09569_ _09569_/A _09569_/B vssd1 vssd1 vccd1 vccd1 _09570_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12580_ _12580_/A _12580_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[4] sky130_fd_sc_hd__xnor2_4
X_11600_ _11706_/B _11600_/B vssd1 vssd1 vccd1 vccd1 _11614_/A sky130_fd_sc_hd__or2_1
XFILLER_0_93_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12252__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11531_ _11414_/A _11414_/B _11415_/Y vssd1 vssd1 vccd1 vccd1 _11536_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_92_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11462_ _11462_/A _11462_/B _11636_/A vssd1 vssd1 vccd1 vccd1 _11462_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_123_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13201_ _13309_/CLK hold60/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dfxtp_1
X_11393_ reg1_val[17] _11099_/B _12487_/S vssd1 vssd1 vccd1 vccd1 _11393_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__11977__A _11977_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ _11429_/A _10413_/B vssd1 vssd1 vccd1 vccd1 _10415_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12960__B1 _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ hold293/A _13131_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _13132_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_103_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10344_ _10208_/A _10208_/B _10207_/A vssd1 vssd1 vccd1 vccd1 _10349_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09708__A1 _09183_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13063_ _13063_/A _13063_/B vssd1 vssd1 vccd1 vccd1 _13063_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__07719__B1 _07179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10275_ _10224_/A _10222_/X _10221_/X vssd1 vssd1 vccd1 vccd1 _10360_/A sky130_fd_sc_hd__a21oi_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12014_ _12014_/A _12014_/B vssd1 vssd1 vccd1 vccd1 _12029_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_88_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12916_ _12946_/A hold220/X vssd1 vssd1 vccd1 vccd1 _13228_/D sky130_fd_sc_hd__and2_1
X_12847_ hold54/X hold272/X vssd1 vssd1 vccd1 vccd1 _13067_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_68_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12778_ hold79/X _12778_/B vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__or2_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07430__A _09622_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11729_ _11892_/A _11729_/B vssd1 vssd1 vccd1 vccd1 _11767_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07670__A2 _10677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10791__A _11499_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12951__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07973__A3 _07322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08940_ _08940_/A _08940_/B vssd1 vssd1 vccd1 vccd1 _08946_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11506__A1 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08871_ _08870_/A _08870_/B _08872_/A vssd1 vssd1 vccd1 vccd1 _08871_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11506__B2 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07822_ _07079_/A _07079_/B _08758_/A2 vssd1 vssd1 vccd1 vccd1 _07824_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__08135__A0 _08836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _08004_/B _07753_/B vssd1 vssd1 vccd1 vccd1 _07754_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__12230__B _12230_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06704_ _06704_/A _06704_/B vssd1 vssd1 vccd1 vccd1 _06705_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_79_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06866__D _06866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07684_ _07678_/A _07678_/B _07678_/C vssd1 vssd1 vccd1 vccd1 _07685_/C sky130_fd_sc_hd__a21o_1
XANTENNA__09883__B1 _10433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07489__A2 fanout46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06635_ reg2_val[23] _06729_/B _06680_/B1 _06634_/Y vssd1 vssd1 vccd1 vccd1 _07119_/A
+ sky130_fd_sc_hd__o2bb2a_2
X_09423_ _11134_/B2 _09752_/B fanout13/X fanout57/X vssd1 vssd1 vccd1 vccd1 _09424_/B
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__11561__S _11738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09354_ _09350_/X _09353_/X _10246_/S vssd1 vssd1 vccd1 vccd1 _09354_/X sky130_fd_sc_hd__mux2_1
X_06566_ instruction[3] _06567_/B vssd1 vssd1 vccd1 vccd1 is_load sky130_fd_sc_hd__nor2_8
X_08305_ _09180_/A _08305_/B _08305_/C vssd1 vssd1 vccd1 vccd1 _08308_/B sky130_fd_sc_hd__and3_1
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09285_ _09478_/B2 _07278_/B _09476_/A fanout7/X vssd1 vssd1 vccd1 vccd1 _09286_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_105_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08236_ _09888_/B2 _08477_/B _08776_/B1 _12736_/A vssd1 vssd1 vccd1 vccd1 _08237_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_34_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10796__A2 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08167_ _08167_/A _08167_/B vssd1 vssd1 vccd1 vccd1 _08207_/B sky130_fd_sc_hd__xor2_4
X_07118_ _07111_/B _07128_/B _07111_/C _07135_/B vssd1 vssd1 vccd1 vccd1 _07119_/B
+ sky130_fd_sc_hd__a31o_1
X_08098_ _08853_/A _08098_/B vssd1 vssd1 vccd1 vccd1 _08154_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__08171__A _08733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07049_ _07077_/A _07075_/A _07049_/C _07167_/A vssd1 vssd1 vccd1 vccd1 _07050_/C
+ sky130_fd_sc_hd__and4_1
XFILLER_0_101_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10060_ _10061_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _10060_/X sky130_fd_sc_hd__or2_1
XANTENNA__07177__A1 _07192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08126__B1 _08776_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11037__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ _10726_/Y _10959_/B _10846_/X vssd1 vssd1 vccd1 vccd1 _10962_/Y sky130_fd_sc_hd__a21oi_1
X_12701_ _12705_/B _12701_/B vssd1 vssd1 vccd1 vccd1 loadstore_address[28] sky130_fd_sc_hd__nor2_8
XANTENNA__06588__A2_N _06752_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10893_ _10894_/A _10894_/B vssd1 vssd1 vccd1 vccd1 _11005_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_742 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12632_ reg1_val[14] _12632_/B vssd1 vssd1 vccd1 vccd1 _12633_/B sky130_fd_sc_hd__or2_1
XFILLER_0_93_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12563_ _12563_/A _12563_/B vssd1 vssd1 vccd1 vccd1 _12564_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_26_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12494_ _12551_/A _12488_/B _12500_/A vssd1 vssd1 vccd1 vccd1 _12495_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11514_ _11618_/D _11514_/B vssd1 vssd1 vccd1 vccd1 _11516_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11445_ _11443_/X _11445_/B vssd1 vssd1 vccd1 vccd1 _11446_/B sky130_fd_sc_hd__and2b_1
XANTENNA__12933__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07404__A2 _12768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11376_ _11550_/A _11376_/B vssd1 vssd1 vccd1 vccd1 _11730_/B sky130_fd_sc_hd__xnor2_2
X_13115_ hold280/X _13165_/A2 _13114_/X _13146_/B2 vssd1 vssd1 vccd1 vccd1 hold281/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ _10027_/A _10027_/B _10161_/B _10159_/Y vssd1 vssd1 vccd1 vccd1 _10341_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _13086_/A hold285/X vssd1 vssd1 vccd1 vccd1 _13286_/D sky130_fd_sc_hd__and2_1
X_10258_ hold292/A _09385_/C _10514_/C _12339_/B1 vssd1 vssd1 vccd1 vccd1 _10258_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10189_ _10190_/A _10190_/B vssd1 vssd1 vccd1 vccd1 _10346_/B sky130_fd_sc_hd__and2b_1
XANTENNA__08668__A1 _07173_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08668__B2 _07182_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07340__B2 fanout83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07340__A1 _10927_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11424__B1 _12150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09070_ _09070_/A _09070_/B _09070_/C _09070_/D vssd1 vssd1 vccd1 vccd1 _09070_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_72_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10778__A2 _11134_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08021_ _08021_/A _08021_/B vssd1 vssd1 vccd1 vccd1 _08023_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11188__C1 _12277_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout6 fanout7/X vssd1 vssd1 vccd1 vccd1 fanout6/X sky130_fd_sc_hd__buf_6
X_09972_ _10752_/S _09971_/Y _09214_/A vssd1 vssd1 vccd1 vccd1 _09972_/Y sky130_fd_sc_hd__a21boi_2
X_08923_ _08923_/A _08923_/B vssd1 vssd1 vccd1 vccd1 _08925_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__08356__B1 _08835_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout297_A _11647_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08854_ _07031_/Y _09925_/A1 _07179_/Y _08854_/B2 vssd1 vssd1 vccd1 vccd1 _08855_/B
+ sky130_fd_sc_hd__o22a_1
X_07805_ _08420_/B _09295_/B _08835_/B1 _08854_/B2 vssd1 vssd1 vccd1 vccd1 _07806_/B
+ sky130_fd_sc_hd__o22a_1
X_08785_ _08785_/A _08785_/B vssd1 vssd1 vccd1 vccd1 _08798_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__08659__A1 _08841_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ _08857_/A _07736_/B vssd1 vssd1 vccd1 vccd1 _07737_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08659__B2 _08841_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06893__B _12721_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07667_ _07401_/A _07400_/C _07400_/B vssd1 vssd1 vccd1 vccd1 _07678_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07331__B2 _09888_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07331__A1 _08681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06618_ reg1_val[26] _07153_/A vssd1 vssd1 vccd1 vccd1 _06619_/B sky130_fd_sc_hd__or2_1
XFILLER_0_48_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07598_ _07274_/A _07273_/Y _07271_/Y vssd1 vssd1 vccd1 vccd1 _07603_/A sky130_fd_sc_hd__a21o_2
X_09406_ _09438_/B _09272_/B _09281_/B _09282_/B _09282_/A vssd1 vssd1 vccd1 vccd1
+ _09421_/A sky130_fd_sc_hd__a32o_2
X_06549_ pred_val instruction[1] vssd1 vssd1 vccd1 vccd1 _06881_/C sky130_fd_sc_hd__and2_1
XFILLER_0_75_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09337_ _08594_/B _08595_/A _08593_/X vssd1 vssd1 vccd1 vccd1 _09337_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_117_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09268_ fanout69/X fanout95/X fanout54/X _12762_/A vssd1 vssd1 vccd1 vccd1 _09269_/B
+ sky130_fd_sc_hd__o22a_1
X_08219_ _08283_/A _08283_/B vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_105_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13168__B1 _13168_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09199_ instruction[3] _09199_/B instruction[4] vssd1 vssd1 vccd1 vccd1 _09199_/X
+ sky130_fd_sc_hd__or3b_1
XFILLER_0_90_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11230_ _11229_/B _11230_/B vssd1 vssd1 vccd1 vccd1 _11231_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11320__A _11429_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ _11162_/B _11162_/A vssd1 vssd1 vccd1 vccd1 _11217_/A sky130_fd_sc_hd__nand2b_1
X_10112_ _10249_/S _10112_/B vssd1 vssd1 vccd1 vccd1 _10112_/X sky130_fd_sc_hd__or2_1
XFILLER_0_101_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11092_ _11092_/A vssd1 vssd1 vccd1 vccd1 _11092_/Y sky130_fd_sc_hd__inv_2
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12151__A _12200_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10043_ _10894_/A _10043_/B vssd1 vssd1 vccd1 vccd1 _10050_/A sky130_fd_sc_hd__xnor2_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
X_11994_ hold173/A _12124_/B _12059_/B _12290_/C1 vssd1 vssd1 vccd1 vccd1 _11995_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_98_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10945_ _10945_/A _10945_/B vssd1 vssd1 vccd1 vccd1 _10947_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07873__A2 _08692_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08076__A _08394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ hold195/A _11559_/A _10983_/B _12290_/C1 vssd1 vssd1 vccd1 vccd1 _10876_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_42_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11406__B1 _12230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12615_ _12623_/A _12615_/B vssd1 vssd1 vccd1 vccd1 _12617_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_109_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12546_ _12546_/A _12546_/B vssd1 vssd1 vccd1 vccd1 _12548_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_109_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12477_ _12478_/A _12478_/B _12478_/C vssd1 vssd1 vccd1 vccd1 _12485_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _10694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11428_ _11532_/B _11428_/B vssd1 vssd1 vccd1 vccd1 _11437_/A sky130_fd_sc_hd__and2_1
XFILLER_0_22_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08586__B1 _09476_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11359_ _11264_/A _11264_/B _11261_/X vssd1 vssd1 vccd1 vccd1 _11360_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12134__A1 _11381_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ _13029_/A _13029_/B vssd1 vssd1 vccd1 vccd1 _13030_/B sky130_fd_sc_hd__nand2_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09073__C _09073_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09550__A2 _10377_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08570_ _08570_/A _08570_/B vssd1 vssd1 vccd1 vccd1 _08583_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07521_ _09898_/A _07521_/B vssd1 vssd1 vccd1 vccd1 _07524_/A sky130_fd_sc_hd__xor2_2
XANTENNA__11645__B1 _11184_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08510__B1 _09273_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07452_ _07464_/A _07464_/B vssd1 vssd1 vccd1 vccd1 _07452_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07383_ _07383_/A _07383_/B _07383_/C vssd1 vssd1 vccd1 vccd1 _07384_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09122_ _09118_/X _09121_/X _09676_/S vssd1 vssd1 vccd1 vccd1 _09122_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09053_ _10617_/B _10617_/C vssd1 vssd1 vccd1 vccd1 _10740_/B sky130_fd_sc_hd__and2_1
XANTENNA_fanout212_A _09362_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08004_ _10015_/A _08004_/B vssd1 vssd1 vccd1 vccd1 _08004_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap240 _09194_/Y vssd1 vssd1 vccd1 vccd1 _11838_/A2 sky130_fd_sc_hd__buf_4
XANTENNA__12373__A1 _12373_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08041__A2 _08348_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_6_0_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11794__B _12304_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09955_ _09955_/A _09955_/B vssd1 vssd1 vccd1 vccd1 _09958_/B sky130_fd_sc_hd__xnor2_4
X_08906_ _08906_/A _08906_/B vssd1 vssd1 vccd1 vccd1 _08907_/B sky130_fd_sc_hd__or2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ _09887_/A _09887_/B vssd1 vssd1 vccd1 vccd1 _10030_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_99_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08837_ _07969_/A _07322_/A _07322_/B fanout47/X _08837_/B2 vssd1 vssd1 vccd1 vccd1
+ _08838_/B sky130_fd_sc_hd__o32a_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _08768_/A _08768_/B _08768_/C vssd1 vssd1 vccd1 vccd1 _08768_/Y sky130_fd_sc_hd__nor3_1
X_08699_ _08699_/A _08699_/B vssd1 vssd1 vccd1 vccd1 _08700_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07719_ _09252_/A _11222_/A _07179_/A _09253_/A vssd1 vssd1 vccd1 vccd1 _07720_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10439__B2 _11688_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10439__A1 _11704_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11100__A2 _06928_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10730_ _10730_/A _10730_/B vssd1 vssd1 vccd1 vccd1 _10960_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10661_ _10662_/A _10662_/B _10662_/C vssd1 vssd1 vccd1 vccd1 _10663_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_82_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12400_ _12401_/A _12401_/B _12401_/C vssd1 vssd1 vccd1 vccd1 _12408_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_118_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12061__B1 _12290_/C1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10592_ _10592_/A _10592_/B vssd1 vssd1 vccd1 vccd1 _10595_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_8_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12331_ _12332_/B _12332_/C hold231/A vssd1 vssd1 vccd1 vccd1 _12331_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_23_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12262_ _12263_/A _12263_/B vssd1 vssd1 vccd1 vccd1 _12308_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11213_ curr_PC[15] _11213_/B vssd1 vssd1 vccd1 vccd1 _11314_/C sky130_fd_sc_hd__and2_2
XFILLER_0_31_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11572__C1 _11400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12193_ _09183_/Y _12181_/B _09835_/X _09158_/S _12192_/Y vssd1 vssd1 vccd1 vccd1
+ _12194_/A sky130_fd_sc_hd__a221o_1
X_11144_ _11262_/B _11143_/B _11143_/C vssd1 vssd1 vccd1 vccd1 _11145_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10127__B1 _11838_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11075_ _12278_/A _11000_/X _11215_/C _09110_/X vssd1 vssd1 vccd1 vccd1 _11076_/B
+ sky130_fd_sc_hd__a31o_1
X_10026_ _10027_/A _10027_/B vssd1 vssd1 vccd1 vccd1 _10161_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07543__A1 _09772_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07543__B2 _08821_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06751__C1 _12588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11977_ _11977_/A _11977_/B vssd1 vssd1 vccd1 vccd1 _11977_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10928_ _10928_/A _10928_/B vssd1 vssd1 vccd1 vccd1 _10930_/B sky130_fd_sc_hd__xnor2_1
X_10859_ _10859_/A _10859_/B vssd1 vssd1 vccd1 vccd1 _10860_/B sky130_fd_sc_hd__xnor2_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08534__A _09898_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12529_ _12529_/A _12529_/B vssd1 vssd1 vccd1 vccd1 _12530_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08271__A2 _08774_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06989__A _06989_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10905__A2 _11431_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06952_ _08544_/A _08544_/B vssd1 vssd1 vccd1 vccd1 _06952_/Y sky130_fd_sc_hd__nand2_2
X_09740_ _10658_/A _09740_/B vssd1 vssd1 vccd1 vccd1 _09748_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
.ends

