// This is the unpowered netlist.
module execution_unit (busy,
    dest_pred_val,
    int_return,
    is_load,
    is_store,
    pred_val,
    rst,
    sign_extend,
    take_branch,
    wb_clk_i,
    curr_PC,
    dest_idx,
    dest_mask,
    dest_pred,
    dest_val,
    instruction,
    loadstore_address,
    loadstore_dest,
    loadstore_size,
    new_PC,
    pred_idx,
    reg1_idx,
    reg1_val,
    reg2_idx,
    reg2_val);
 output busy;
 output dest_pred_val;
 output int_return;
 output is_load;
 output is_store;
 input pred_val;
 input rst;
 output sign_extend;
 output take_branch;
 input wb_clk_i;
 input [27:0] curr_PC;
 output [5:0] dest_idx;
 output [1:0] dest_mask;
 output [2:0] dest_pred;
 output [31:0] dest_val;
 input [41:0] instruction;
 output [31:0] loadstore_address;
 output [5:0] loadstore_dest;
 output [1:0] loadstore_size;
 output [27:0] new_PC;
 output [2:0] pred_idx;
 output [5:0] reg1_idx;
 input [31:0] reg1_val;
 output [5:0] reg2_idx;
 input [31:0] reg2_val;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire busy_l;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire div_complete;
 wire \div_counter[0] ;
 wire \div_counter[1] ;
 wire \div_counter[2] ;
 wire \div_counter[3] ;
 wire \div_counter[4] ;
 wire \div_res[0] ;
 wire \div_res[10] ;
 wire \div_res[11] ;
 wire \div_res[12] ;
 wire \div_res[13] ;
 wire \div_res[14] ;
 wire \div_res[15] ;
 wire \div_res[16] ;
 wire \div_res[17] ;
 wire \div_res[18] ;
 wire \div_res[19] ;
 wire \div_res[1] ;
 wire \div_res[20] ;
 wire \div_res[21] ;
 wire \div_res[22] ;
 wire \div_res[23] ;
 wire \div_res[24] ;
 wire \div_res[25] ;
 wire \div_res[26] ;
 wire \div_res[27] ;
 wire \div_res[28] ;
 wire \div_res[29] ;
 wire \div_res[2] ;
 wire \div_res[30] ;
 wire \div_res[31] ;
 wire \div_res[3] ;
 wire \div_res[4] ;
 wire \div_res[5] ;
 wire \div_res[6] ;
 wire \div_res[7] ;
 wire \div_res[8] ;
 wire \div_res[9] ;
 wire \div_shifter[0] ;
 wire \div_shifter[10] ;
 wire \div_shifter[11] ;
 wire \div_shifter[12] ;
 wire \div_shifter[13] ;
 wire \div_shifter[14] ;
 wire \div_shifter[15] ;
 wire \div_shifter[16] ;
 wire \div_shifter[17] ;
 wire \div_shifter[18] ;
 wire \div_shifter[19] ;
 wire \div_shifter[1] ;
 wire \div_shifter[20] ;
 wire \div_shifter[21] ;
 wire \div_shifter[22] ;
 wire \div_shifter[23] ;
 wire \div_shifter[24] ;
 wire \div_shifter[25] ;
 wire \div_shifter[26] ;
 wire \div_shifter[27] ;
 wire \div_shifter[28] ;
 wire \div_shifter[29] ;
 wire \div_shifter[2] ;
 wire \div_shifter[30] ;
 wire \div_shifter[31] ;
 wire \div_shifter[32] ;
 wire \div_shifter[33] ;
 wire \div_shifter[34] ;
 wire \div_shifter[35] ;
 wire \div_shifter[36] ;
 wire \div_shifter[37] ;
 wire \div_shifter[38] ;
 wire \div_shifter[39] ;
 wire \div_shifter[3] ;
 wire \div_shifter[40] ;
 wire \div_shifter[41] ;
 wire \div_shifter[42] ;
 wire \div_shifter[43] ;
 wire \div_shifter[44] ;
 wire \div_shifter[45] ;
 wire \div_shifter[46] ;
 wire \div_shifter[47] ;
 wire \div_shifter[48] ;
 wire \div_shifter[49] ;
 wire \div_shifter[4] ;
 wire \div_shifter[50] ;
 wire \div_shifter[51] ;
 wire \div_shifter[52] ;
 wire \div_shifter[53] ;
 wire \div_shifter[54] ;
 wire \div_shifter[55] ;
 wire \div_shifter[56] ;
 wire \div_shifter[57] ;
 wire \div_shifter[58] ;
 wire \div_shifter[59] ;
 wire \div_shifter[5] ;
 wire \div_shifter[60] ;
 wire \div_shifter[61] ;
 wire \div_shifter[62] ;
 wire \div_shifter[63] ;
 wire \div_shifter[6] ;
 wire \div_shifter[7] ;
 wire \div_shifter[8] ;
 wire \div_shifter[9] ;
 wire divi1_sign;
 wire \divi2_l[0] ;
 wire \divi2_l[10] ;
 wire \divi2_l[11] ;
 wire \divi2_l[12] ;
 wire \divi2_l[13] ;
 wire \divi2_l[14] ;
 wire \divi2_l[15] ;
 wire \divi2_l[16] ;
 wire \divi2_l[17] ;
 wire \divi2_l[18] ;
 wire \divi2_l[19] ;
 wire \divi2_l[1] ;
 wire \divi2_l[20] ;
 wire \divi2_l[21] ;
 wire \divi2_l[22] ;
 wire \divi2_l[23] ;
 wire \divi2_l[24] ;
 wire \divi2_l[25] ;
 wire \divi2_l[26] ;
 wire \divi2_l[27] ;
 wire \divi2_l[28] ;
 wire \divi2_l[29] ;
 wire \divi2_l[2] ;
 wire \divi2_l[30] ;
 wire \divi2_l[31] ;
 wire \divi2_l[3] ;
 wire \divi2_l[4] ;
 wire \divi2_l[5] ;
 wire \divi2_l[6] ;
 wire \divi2_l[7] ;
 wire \divi2_l[8] ;
 wire \divi2_l[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(reg1_val[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(reg1_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(reg1_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(reg1_val[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(reg1_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(reg1_val[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(reg1_val[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(reg1_val[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(reg1_val[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(reg1_val[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_00360_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(reg1_val[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(reg1_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(reg1_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(reg1_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(reg1_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(reg1_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(reg1_val[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(reg2_val[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(reg2_val[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(reg2_val[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(reg2_val[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(reg2_val[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(reg2_val[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(reg2_val[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(reg2_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(reg2_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(reg2_val[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(reg2_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(reg2_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(reg2_val[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(instruction[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(reg2_val[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(instruction[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(instruction[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(reg1_val[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(reg1_val[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(reg1_val[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(reg1_val[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(instruction[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(reg1_val[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(reg1_val[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(reg1_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(reg1_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(reg1_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(reg2_val[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(reg1_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(reg1_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(instruction[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(reg1_val[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(instruction[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(reg1_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(reg1_val[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06577__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__06584__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__06591__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06593__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06595__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06597__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06601__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__C1 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06611__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06616__A2 (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06617__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06618__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06619__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06619__B (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06620__A2_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06621__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06626__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__B (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06628__A2_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06629__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06633__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06634__B (.DIODE(_05067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06635__A2_N (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06636__B1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06640__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06641__B (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06642__A2_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06647__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06648__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06648__B (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06649__A2_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06650__A_N (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06651__B (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06653__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06654__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06654__B (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06655__A2_N (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06656__B1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06660__B (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06662__A2 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06663__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06663__B (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__B (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06665__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__B (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__A2_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06675__B (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__06676__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06676__B (.DIODE(_05523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__A2_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__A_N (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__B (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06682__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06682__B (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06683__A2_N (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06684__A_N (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06685__B (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06688__B (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__A2_N (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06690__A_N (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06691__B (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06692__B (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06694__B (.DIODE(_05706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06695__A2_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06696__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06699__B (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06703__B (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06704__A2_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06705__A_N (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06706__B (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06710__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06710__B (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06711__A2_N (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06712__B1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06717__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06717__B (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06718__A2_N (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06719__A_N (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06720__B (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06723__A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06723__B (.DIODE(_05962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06724__A2_N (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06725__B1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06726__B (.DIODE(_05980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06727__B (.DIODE(_05980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06729__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06730__A2 (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06731__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06731__B (.DIODE(_06031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06732__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06732__B (.DIODE(_06031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06734__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06735__A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06735__A3 (.DIODE(_05067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__B (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06737__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06737__B (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06740__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06740__A3 (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06741__B (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06742__B (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06744__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__A3 (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06746__B (.DIODE(_06151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06747__B (.DIODE(_06151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06749__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06750__A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06750__A3 (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06755__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06756__A1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06756__A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06756__A3 (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06757__B (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06758__B (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__A3 (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__B1 (.DIODE(_06274_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06766__B (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06767__A3 (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06771__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06772__A3 (.DIODE(_05523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06772__B1 (.DIODE(_06319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06776__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__A3 (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__B1 (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__C1 (.DIODE(_05706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__D1 (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__C_N (.DIODE(_05706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06784__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06784__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__A2 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__06791__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06792__A3 (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06792__B1 (.DIODE(_06339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__A3 (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__B1 (.DIODE(_06339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06794__B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__06795__B (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__06797__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06798__A3 (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06798__B1 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06799__A3 (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06799__B1 (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__B (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06801__B (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06803__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06804__A3 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06804__B1 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06805__A3 (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06805__B1 (.DIODE(_06351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06806__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__06807__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__06808__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__06810__B (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__06811__A3 (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06811__B1 (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06812__A3 (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06812__B1 (.DIODE(_06358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__B (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__B (.DIODE(_05962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06816__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__06818__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06819__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06819__B (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06821__B (.DIODE(_06352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06823__B (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__06825__B (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__06837__A_N (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06841__A_N (.DIODE(_06151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06843__A_N (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06845__A_N (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06845__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__06847__A_N (.DIODE(_06031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06847__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__B (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06855__B (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06857__B (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__B (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06861__B (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__A2 (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06870__B (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__B (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__B (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__06912__A1 (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06912__B1 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__B (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06919__A1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__B (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06924__B (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__B (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__B (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__C (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__B (.DIODE(_04596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__A2 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__B1 (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__06955__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__C (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__C (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__B (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06969__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__06969__B (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__B (.DIODE(_06352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__C (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__D (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__A (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__C (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__D (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__06972__D (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__06976__B (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06977__A (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06977__B (.DIODE(_06151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06977__D (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06978__A (.DIODE(_06031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06978__B (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__A (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__A (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__C (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__A (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__B (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__A (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__B (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__A (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__B (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__A (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__A (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__A (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__B1 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__B (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__07005__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__A2 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__07009__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07010__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__A (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__S (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__A (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07017__A1 (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__C1 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__B (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07020__A (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07020__B (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__B1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07022__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07024__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07026__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07027__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07028__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07029__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07034__A1 (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__A (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__A (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07037__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__S (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07040__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07044__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__A2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__B2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07067__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07069__B1 (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__A (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__B (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__A (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__B (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07073__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07073__C_N (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__B1 (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07078__A (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__A (.DIODE(_00169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__B (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__A (.DIODE(_00169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__B (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__A (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__A (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07098__S (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07107__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07107__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07109__C (.DIODE(_00200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A4 (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07117__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__07117__B (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07117__C (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__A3 (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__A (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__A2 (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07132__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__07136__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__S (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__B1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__B (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__B (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__D (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__A (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07143__B (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__B (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__C (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07148__A (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__A (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A4 (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__A_N (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__S (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__A1 (.DIODE(_00240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__A1 (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__A2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__B1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__C1 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__A2 (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__A3 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__B1 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__C1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__07165__A (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07172__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__A (.DIODE(_06352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07174__S (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__A1 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__B1 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07186__A1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__07187__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__07189__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07190__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__A (.DIODE(_06151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__A (.DIODE(_06151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A1 (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__B (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__A2 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07205__A4 (.DIODE(_00200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__C (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__S (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A3 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__A2 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__B2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07229__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07232__A (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07233__A (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__C1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07253__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__S (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__A1 (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__A (.DIODE(_06031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__A (.DIODE(_06031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__B (.DIODE(_00357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__A (.DIODE(_00338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__B (.DIODE(_00357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__A (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__A (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__A1 (.DIODE(_06151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__A (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07274__A (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__B2 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__B1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A1 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__B2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07305__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__A (.DIODE(_00405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__B (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__A (.DIODE(_00405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__B (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__A1 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__B2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07332__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07334__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__07337__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07337__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07337__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07337__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07338__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__A1 (.DIODE(_00240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__B1 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__B1 (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__A1 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__B2 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__C (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__A2 (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07360__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__B2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__B2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07390__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A1 (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__B1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07396__A1 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07396__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07396__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07396__B2 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__B (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07422__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07422__A2 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07422__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07422__B2 (.DIODE(_00240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__A1 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07449__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07449__A2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07449__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07449__B2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07450__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__A2 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__B1 (.DIODE(_00330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07471__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__A1 (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__B2 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07476__A1 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07476__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07476__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07476__B2 (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07477__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__B1 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__A1 (.DIODE(_00240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07510__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07510__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07510__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07510__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__B2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07525__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__A2 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__A1 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__B2 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__B1 (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__B1 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07553__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__A1 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__B1 (.DIODE(_00330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__A1 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07583__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07585__A3 (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__B (.DIODE(_00678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__B1 (.DIODE(_00678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__B1 (.DIODE(_00678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__B2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__A (.DIODE(_00678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__B (.DIODE(_00698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07608__A (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07608__B (.DIODE(_00698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__A2 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__B1 (.DIODE(_00700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__B1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07612__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07616__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07616__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07616__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07616__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07622__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A2 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__B1 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__A2 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07632__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07636__A1 (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07636__A2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07636__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07636__B2 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07637__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__B2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07685__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07685__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07685__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07685__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__A1 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__B1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__B2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07695__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__B2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__B1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07719__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__A1 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__B2 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__B1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__B2 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__B1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07786__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__B1 (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__B2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__A1 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__B2 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__A1 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__B2 (.DIODE(_00240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A1 (.DIODE(_06544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A2 (.DIODE(_06545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__B1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__B (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__C (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07840__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__A0 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__B2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07847__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07849__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__07851__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07851__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07851__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07851__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07852__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A1 (.DIODE(_00240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__B2 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07907__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__07907__B (.DIODE(_00161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07907__C (.DIODE(_00162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__A1 (.DIODE(_00169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__A2 (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__B1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__B2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__A (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__A2 (.DIODE(_00179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__B1 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__A1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__B2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07923__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__A1 (.DIODE(_00169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__A2 (.DIODE(_00170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__B1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__B (.DIODE(_00179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07984__B1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__07985__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__A2 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__B1 (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07995__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08019__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08021__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08031__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08033__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08035__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__A2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08045__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__B2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__B1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08092__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08102__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08106__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08106__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08106__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08106__B2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__B (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__A0 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__B2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__B1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08129__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__B2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08147__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08149__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08199__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08199__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08203__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08205__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08207__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08237__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08238__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08238__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08238__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08238__B2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08239__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08242__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08244__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08248__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08252__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08253__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08253__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08253__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08253__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08293__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08299__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08331__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08333__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08334__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__A2 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__B1 (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__B2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__A (.DIODE(_01428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__A (.DIODE(_01428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08344__B1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08369__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__B2 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__A (.DIODE(_00342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08380__B (.DIODE(_01471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__B2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__B (.DIODE(_01471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08390__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08411__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__A1 (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08416__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08418__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08440__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08442__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08453__B2 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08456__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__A2 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08458__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08473__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08474__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08474__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08474__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08474__B2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08484__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08484__B (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__08487__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08501__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08501__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08501__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08501__B2 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08502__A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08504__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__B1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08508__A (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08508__B (.DIODE(_01599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__B2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08514__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__08515__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08515__A2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08515__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08515__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08516__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08529__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08539__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__B (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__A_N (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__B1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__08559__B2 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__A2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A2 (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__B1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__A2 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__B1 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08575__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08577__A (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08579__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08598__B (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__B2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08602__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__08612__B1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08613__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__08614__B1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__A2 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08616__B1 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__08627__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08627__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08627__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08627__B2 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08628__A (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__A2 (.DIODE(_00240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__B1 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__08633__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__08633__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08633__B2 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08641__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__A0 (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__A1 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__A2 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08647__B1 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__B1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__A (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__A2 (.DIODE(_00240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__B1 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08655__B2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__08657__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08657__B (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__A (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__B1 (.DIODE(_00240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__A0 (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08713__A1 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__08716__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__A2 (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__C (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__A2 (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08816__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__08816__A2 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08816__B1 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08816__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08818__A1 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08818__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__08818__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__08818__B2 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08819__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__A1 (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__B1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__B2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__08836__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__08838__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__08842__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__08846__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__08848__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__A2 (.DIODE(_00700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__B1 (.DIODE(_01951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__A2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__B1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08864__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__B (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__D (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__A4 (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08873__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08874__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__08878__A1 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08878__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08878__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__08878__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__B2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08886__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08887__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__08887__A2 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08887__B1 (.DIODE(_00330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08887__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__08888__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__A2 (.DIODE(_01889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__A3 (.DIODE(_01959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__A2 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__A1 (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__B2 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08931__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__B1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__08936__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__08950__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__A2 (.DIODE(_00160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__08952__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__08956__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08960__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__08962__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08966__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__08966__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08966__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08966__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08972__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__08974__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__A1 (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08976__B2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__A2 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08978__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08983__B (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__08988__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__08988__B1 (.DIODE(_00678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08988__D1 (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__A2 (.DIODE(_02078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__B2 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__B2 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__A (.DIODE(_00678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__A2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__B2 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__09004__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__B2 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09006__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09010__B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09030__A (.DIODE(_02110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09031__A (.DIODE(_02110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09047__A3 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09048__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09048__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09048__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09048__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__A2 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09052__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__A1 (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__B1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09054__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09055__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__A2 (.DIODE(_00160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09071__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09073__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__09082__A1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09082__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__09082__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09082__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09083__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09087__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A2 (.DIODE(_00405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__A3 (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__B1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__09093__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__A (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__A1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__B1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__A (.DIODE(_06364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09103__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__A1 (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09115__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__A2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__B1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09117__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09145__B (.DIODE(_02236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__B (.DIODE(_02236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09148__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09155__A0 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__09156__S (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09179__A0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__A0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__09195__A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A0 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__A0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__09220__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__09230__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__A2 (.DIODE(_02325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__B (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__A1 (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__A (.DIODE(_06352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A2 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A0 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__S (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__A2 (.DIODE(_02349_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09266__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A2 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__B1 (.DIODE(_00330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__B2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__B1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09272__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__B1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__B2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09290__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__A2 (.DIODE(_00184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09298__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__A2 (.DIODE(_00698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09300__B1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__B (.DIODE(_00405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__C (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__A (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__B1 (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__B1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__B1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09306__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__B2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09326__B2 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__A2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__B1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09340__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__B1 (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__B2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A (.DIODE(_02353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__B (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__A (.DIODE(_02353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__B (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__B2 (.DIODE(_02236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__S (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09411__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__B1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09415__A1 (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09417__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__09419__A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__09420__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__A (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__B (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__C_N (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__B2 (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__A2_N (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__B2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__A2 (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__A2 (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__A (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09435__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09439__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__09439__A2 (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__A1 (.DIODE(_02531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__A1 (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09448__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__A2 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__B1 (.DIODE(_00330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09450__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__A2 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__B1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09456__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__B1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09480__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09482__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__A3 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__A (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__B1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09516__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__A2 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__B1 (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__A (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__B (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__A (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__B (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__B (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A2 (.DIODE(_02236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__B1 (.DIODE(_02353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__B2 (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A1 (.DIODE(_02353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A2 (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09556__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__09559__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__S (.DIODE(_06352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09575__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09583__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09584__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A2 (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__B1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__09587__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__09588__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__09592__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09594__B (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__B (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__C1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09598__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09598__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__A1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__B2 (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09612__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09612__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09612__B1 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09612__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__A2 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__B1 (.DIODE(_00330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09616__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__09626__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__A1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09628__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__A2 (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__B1 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__09632__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__09648__A (.DIODE(_00342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__A2 (.DIODE(_00698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__B (.DIODE(_00405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__C (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09651__B1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09652__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09656__B2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__A (.DIODE(_00338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__09666__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09666__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__09666__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__B2 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__09672__A (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09680__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A (.DIODE(_02695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__B (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09706__A (.DIODE(_02695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09706__B (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A (.DIODE(_02695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__B (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09726__S (.DIODE(_06352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09728__S (.DIODE(_06359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09730__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09732__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__09732__B (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09737__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__09744__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__A1 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__B1 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__09756__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__A1 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__A2 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__B1 (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__A3 (.DIODE(_02827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09759__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__A2 (.DIODE(_02849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__A1 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__A1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__B2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__A2 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__B1 (.DIODE(_00330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09792__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__A (.DIODE(_00338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__A2 (.DIODE(_00405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__A3 (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09796__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09802__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__A2 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09812__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09812__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09812__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09812__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09813__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09814__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09814__B1 (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__A1 (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09823__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__A1 (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__A1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__09834__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__A2 (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__B1 (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__09836__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__A (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09870__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__B1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09877__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__S (.DIODE(_06352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__09887__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__09887__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09887__B1 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09889__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__B1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__B2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__A3 (.DIODE(_02987_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__B1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A2 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__A3 (.DIODE(_02325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__A2 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__B1 (.DIODE(_02974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__B1 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__09921__A1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__09921__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09921__B1 (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09921__B2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__09922__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__A1 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__B1 (.DIODE(_00330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__A1 (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__B2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__A1 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__B2 (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09974__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09974__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__09974__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__09974__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__09975__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__A1 (.DIODE(_02695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__A2 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__B1 (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__A1 (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10006__B (.DIODE(_03092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__10012__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__A1 (.DIODE(_06352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10021__C1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__A1 (.DIODE(_06352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10024__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__B1 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__10040__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__10040__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__10041__A2 (.DIODE(_03113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10042__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10049__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__10052__A1 (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__B1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__C1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__A1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10058__A (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__A2 (.DIODE(_00405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__A3 (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__B1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10059__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10070__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__10070__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10070__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10070__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__10071__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__10073__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__10073__B2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__10079__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__A1 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__B2 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10081__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__B1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__A2 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__B1 (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__A (.DIODE(_00245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__B2 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__A (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__A1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__B1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10115__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__A (.DIODE(_03136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__B (.DIODE(_03221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__A1 (.DIODE(_02855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__A (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__B1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__B (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__S (.DIODE(_06352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10164__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10172__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__10173__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10173__B1 (.DIODE(_02325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10174__A2 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10174__B1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__A1 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__10181__A2 (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10183__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10187__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10193__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A1 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__A2 (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__B1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10207__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10209__A (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__10222__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__A (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__A1 (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__A1 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__A (.DIODE(_00678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__A2 (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__B1 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A (.DIODE(_00245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__B1 (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__A2 (.DIODE(_00698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__B (.DIODE(_00405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__C (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10241__B1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__10244__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__10246__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__A (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__B (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__B1 (.DIODE(_03136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__B2 (.DIODE(_03221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10280__A1 (.DIODE(_03136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10280__A2 (.DIODE(_03221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__B (.DIODE(_03367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__A2 (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__10285__A2 (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10289__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__S (.DIODE(_06352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__S (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__10301__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__A2_N (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__10308__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__A2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10317__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__B (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__A1 (.DIODE(_03136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__A2 (.DIODE(_03221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__B1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__B2 (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__A2 (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__B2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__A (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__B (.DIODE(_02078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__A (.DIODE(_00342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__B1_N (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__10350__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A2 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__B1 (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__A2 (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__B1 (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__A (.DIODE(_00245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__A2 (.DIODE(_00405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__A3 (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__10371__A (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__B2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10384__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__A1 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10386__B2 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10392__A (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__A (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__B (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__A (.DIODE(_03417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__A2 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__A2 (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__C1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__S (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__A2 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__B1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__10442__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__A1 (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__A1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__A1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10451__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__B (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__A (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__A (.DIODE(_00342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__A1 (.DIODE(_00697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__A2 (.DIODE(_00698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__B (.DIODE(_00405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__C (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__10480__B1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A1 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__B2 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__A2 (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__B1 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__A1 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__B2 (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__A (.DIODE(_00245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__A1 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10507__B2 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10539__A (.DIODE(_03620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__B1 (.DIODE(_03625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__A1 (.DIODE(_03273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__A2 (.DIODE(_03360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__B1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__B2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__A1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__A2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__C1 (.DIODE(_03629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__A (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__B (.DIODE(_03630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10549__C (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__B1 (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__S (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__10566__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__A2 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__B1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__10572__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__10572__C1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__A1 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__10578__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__A (.DIODE(_03368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__B (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__C (.DIODE(_03631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__D_N (.DIODE(_03500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__B1 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__B2 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A (.DIODE(_00245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__A2 (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__B1 (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__B2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10599__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10599__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10602__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10603__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10603__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10603__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10603__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__A (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__A1 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__B2 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__B1 (.DIODE(_00342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__A1 (.DIODE(_00342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__A3 (.DIODE(_02067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10616__B (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__B2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10623__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10625__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__A1 (.DIODE(_03418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__A2 (.DIODE(_03498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__B1 (.DIODE(_03620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__B (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10661__D (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10664__A (.DIODE(_03738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__B1 (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A3 (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10683__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__C1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10686__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__A0 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__A1 (.DIODE(_06238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10694__B1 (.DIODE(_03774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10696__A1 (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10696__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__B2 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10702__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__A2 (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__A (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__A (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10713__A1 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10713__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10713__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10713__B2 (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10714__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__A1 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__B2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__A1 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__B2 (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__A (.DIODE(_00678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10725__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__10725__B (.DIODE(_02078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__A1 (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__B2 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10732__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10735__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10735__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10735__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10735__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10736__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10744__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10744__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10744__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10744__B2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10745__A (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__10747__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10748__A (.DIODE(_00342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10749__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__A2 (.DIODE(_03697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__A (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__B (.DIODE(_03738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__A1 (.DIODE(_03620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__A1 (.DIODE(_03367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__A (.DIODE(_03859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__A2 (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__A2 (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10788__A (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__10792__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__B1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10800__B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__10808__A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__10808__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__10809__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__10812__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__10813__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__10817__A1 (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10817__B2 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__B (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__C (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__B1 (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__A1 (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__A3 (.DIODE(_02067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__B2 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10840__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10842__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__A1 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__B2 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10847__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__A2 (.DIODE(_00405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__A3 (.DIODE(_00407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__A1 (.DIODE(_06559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__B2 (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__10856__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10862__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__A (.DIODE(_03738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__B (.DIODE(_03859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10903__A1 (.DIODE(_03417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__A2 (.DIODE(_03984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__A2 (.DIODE(_03984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10908__B1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10910__S (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__10914__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__B1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10923__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__10923__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__A1 (.DIODE(_06151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__A1 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__B2 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__10933__C (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10937__A2 (.DIODE(_03984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A1 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__B2 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__A1 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__B2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__A (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__B1 (.DIODE(_02067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10952__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__A1 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__B2 (.DIODE(_06559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10965__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10970__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__A (.DIODE(_03859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__A1 (.DIODE(_03629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__A1 (.DIODE(_03092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__A2 (.DIODE(_03625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__A2 (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__A2 (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__B1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__S (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__11029__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__11030__A (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__A1 (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__A (.DIODE(_06121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__B (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__A1 (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__A (.DIODE(_03746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__B (.DIODE(_03865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__C (.DIODE(_03984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__D (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__B1 (.DIODE(_04134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__B (.DIODE(_04134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11062__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__A2 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11064__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__A1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__B2 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__A1 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__B2 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11072__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__A1 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__B2 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11074__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11079__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__11080__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11082__S (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__A2 (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11092__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__11093__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__11093__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11123__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__A2 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11126__A2 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__S (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__11132__C1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__11134__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__11138__A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__C1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11149__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__11151__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__A1 (.DIODE(_06086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A1 (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__S (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11163__A2 (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__B2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A1 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B2 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__B2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__A1 (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__B2 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__A1 (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__A2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__B2 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__11198__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__11198__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__A2 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__A1 (.DIODE(_03367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__B (.DIODE(_04309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__B (.DIODE(_04309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11236__B1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__S (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__C1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__11242__A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__C1 (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11254__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11257__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__A1 (.DIODE(_06031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__A1_N (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__11269__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__B (.DIODE(_04309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__D_N (.DIODE(_04202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__B (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11274__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11274__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11274__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11274__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11275__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__A1 (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__B1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11277__A (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__B2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__A (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11285__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11285__B1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__B (.DIODE(_04362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__B (.DIODE(_04362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__A1 (.DIODE(_06559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__B2 (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__A (.DIODE(_00245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__A1 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__B2 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11300__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11306__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11310__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__11310__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11338__A1 (.DIODE(_03417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11339__B (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__B (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__A2 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__A2 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__S (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__11355__S (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__11358__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11360__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__11360__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__A1 (.DIODE(_05980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11361__B1 (.DIODE(_02325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11366__A1_N (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__11368__A1 (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11369__A1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11370__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11372__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11376__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A1 (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A2 (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11378__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11378__A2 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11378__B1 (.DIODE(_00700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11378__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__B1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11382__B2 (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11390__A1 (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11390__A2 (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11390__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__11390__B2 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__A2 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__A1 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__B2 (.DIODE(_06559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11398__A (.DIODE(_00245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__A1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11402__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11403__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__B (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11433__B (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11439__A1 (.DIODE(_03630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11441__A (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__A2 (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__A2 (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11447__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__11448__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__A (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__C1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__A1 (.DIODE(_05934_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__B1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__11459__A2 (.DIODE(_02325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11460__A1 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11465__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__11469__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__A1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__A (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__B (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__B1 (.DIODE(_04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__C (.DIODE(_04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__A1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__B2 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__A2 (.DIODE(_00700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__B1 (.DIODE(_01951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__A (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__A2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11497__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__A1 (.DIODE(_06559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__B2 (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__A2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__11526__A (.DIODE(_04409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11532__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11534__B1 (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11535__A3 (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11535__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__11540__S (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__B1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11548__S (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__A0 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__A1 (.DIODE(_02325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__A (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__B2 (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__A1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__A1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__B1 (.DIODE(_04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11566__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__A (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__B (.DIODE(_04419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__D (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__A1 (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__B2 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11571__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__A1 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__B2 (.DIODE(_06559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11579__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11579__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11579__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11579__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__11583__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11583__A2 (.DIODE(_01951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11583__B1 (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11583__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__A (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11590__A (.DIODE(_04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11591__A (.DIODE(_04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11592__A (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11592__B (.DIODE(_02078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11626__A (.DIODE(_04724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11628__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__11632__A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__11634__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__11643__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__11644__C1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11648__A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__A0 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__11654__A1 (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11654__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__B2 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__B2 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__C1 (.DIODE(_04757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11659__B1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11661__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__A1 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__A2 (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__B1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11666__A1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11666__A3 (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11679__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__A1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__B2 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11683__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__A (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__A (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__B (.DIODE(_04823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__A2 (.DIODE(_04823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__S (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__11727__C1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11733__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__C1 (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11737__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11741__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__B (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11743__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__11743__C1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__11744__A1 (.DIODE(_05668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11744__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__B2 (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__B2 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__C1 (.DIODE(_04854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11752__S (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11753__A3 (.DIODE(_04823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__A1 (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__B1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__B2 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11759__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__A (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__B1 (.DIODE(_00699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11779__A (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11779__B (.DIODE(_02078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11799__B (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11807__B (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__A2 (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__S (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__11820__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__A1 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__C1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11827__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11829__B (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11830__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__11830__C1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__11831__A1 (.DIODE(_05725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11831__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11832__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__11832__B2 (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__B2 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__C1 (.DIODE(_04949_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__C (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__D_N (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11841__A (.DIODE(_04724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11841__D_N (.DIODE(_04918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__A (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__A (.DIODE(_00678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11845__A1 (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11845__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11845__B1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11845__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11846__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__A1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__A2 (.DIODE(_00700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__B1 (.DIODE(_01951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11853__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__11854__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__A1 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11864__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11864__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11864__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11864__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__A (.DIODE(_04813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11891__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__11891__B1 (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__C (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__B1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__S (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__11899__B1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__S (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__11909__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11913__A0 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__A1 (.DIODE(_05609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11915__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11916__B2 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11919__A1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__11920__A1 (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11920__B1 (.DIODE(_05015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11922__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__11923__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__A1 (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__A3 (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__11926__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11926__A2 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11926__B1 (.DIODE(_00700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11926__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11927__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__11928__A_N (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11929__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11943__A (.DIODE(_02079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11945__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__11946__B (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11946__C (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__A1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__A2 (.DIODE(_02079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11973__B (.DIODE(_05098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11974__A2 (.DIODE(_05098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11974__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11976__B1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11978__C1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__11980__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__B1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11988__S (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11990__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__11994__C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__B (.DIODE(_02325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__A2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__C1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A1 (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__11998__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__11998__B2 (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__A1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12001__B1 (.DIODE(_05104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__A1 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A3 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__12007__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__12007__B (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12009__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__12009__B (.DIODE(_02079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12010__A (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__A2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__12017__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__A2 (.DIODE(_00700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__B1 (.DIODE(_01951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__12019__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__A1 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__A (.DIODE(_05009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__B (.DIODE(_05098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__A (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12051__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__B1 (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__S (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__12055__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__12057__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__B1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__S (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__12066__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12070__C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__A0 (.DIODE(_02325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__A1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12072__A1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__A2 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__B1 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12074__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__A1 (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__C1 (.DIODE(_05192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12080__A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12081__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__12084__B (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12085__A_N (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12087__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__12087__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__A3 (.DIODE(_05137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__B1 (.DIODE(_00699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12091__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__A2 (.DIODE(_01951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__B1 (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__12096__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__12121__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__S (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__12126__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__A0 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__S (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12138__B1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__A0 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12144__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12145__A1 (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12145__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12145__B1 (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12145__B2 (.DIODE(_03244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12146__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12146__A2 (.DIODE(_03251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12148__A1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__B1 (.DIODE(_05290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__A1 (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__C1 (.DIODE(_05291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12152__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12153__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__A2 (.DIODE(_00699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__B1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__12158__B (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__12168__A1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12168__B2 (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__A (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__A1 (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__S (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__12190__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__12196__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__12198__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12198__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12204__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__B1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__A0 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12208__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12210__A1 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12210__B1 (.DIODE(_03113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12210__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12212__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__D_N (.DIODE(_05362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12218__A (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__B1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__A1 (.DIODE(_00699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__B2 (.DIODE(_00409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12222__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__B1 (.DIODE(_02067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__B2 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__12227__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__12232__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__12232__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__12233__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__12233__B (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__12233__C (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12253__B1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__B1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__A2 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12272__C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__A2 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__B1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__B1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__C1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__A1 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__A2 (.DIODE(_02968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__B1 (.DIODE(_02974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__A1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__B1 (.DIODE(_05430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__B2 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__B2 (.DIODE(_00699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12282__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__A (.DIODE(_00409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12288__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__12288__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12288__B1 (.DIODE(_00678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12289__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__12289__A3 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__12308__B1 (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__S (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__C1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__B (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__A1 (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__C1 (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12322__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__A2 (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__A2 (.DIODE(_02325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__C1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__A1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__A2 (.DIODE(_02820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__B1 (.DIODE(_02830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__B2 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12331__B (.DIODE(_05472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12332__C1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__B2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12334__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12335__A (.DIODE(_00699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12335__B (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__12356__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12360__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__B1 (.DIODE(_02317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__A (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12368__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__A1 (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12369__C1 (.DIODE(_06476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12371__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__C1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__12377__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12377__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__A2 (.DIODE(_02325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__C1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12379__A1 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12379__B1 (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12379__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__C1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12383__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__A1 (.DIODE(_01951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12387__A1 (.DIODE(_01951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12387__A2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__12401__B1 (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__S (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__12405__B1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__12409__B1 (.DIODE(_02324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12412__A (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12412__B (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12413__A1 (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12413__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__C1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__12419__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__12419__B1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__A0 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12421__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12423__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__12423__B1 (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12423__B2 (.DIODE(_02314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__C1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12427__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__B (.DIODE(_02078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12436__B1 (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12438__A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__B1 (.DIODE(_02323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12444__B (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12446__C1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__B1 (.DIODE(_02330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12452__A2 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12452__B1 (.DIODE(_02315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__A2 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__A3 (.DIODE(_02325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__C1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__A2 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__B2 (.DIODE(_02313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__A1 (.DIODE(_05382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__A2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12460__A0 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__12460__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__A (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12462__A (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12464__A0 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__12464__S (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__12465__A (.DIODE(_05962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12466__A (.DIODE(_05962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12471__S (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12473__A (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12479__A (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12480__A (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12485__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__A (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12487__A (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12493__A (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__A (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__A (.DIODE(_05706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12501__A (.DIODE(_05706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__A (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12508__A (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12514__A (.DIODE(_05523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__A (.DIODE(_05523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12520__S (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__A (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12522__A (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12527__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12528__A (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__A (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__A (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12542__A (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12543__A (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12548__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12549__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12550__A (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12555__A0 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__12555__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12556__A (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12557__A (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__A0 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__12562__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__A (.DIODE(_05067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__A (.DIODE(_05067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12574__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12587__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12593__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__S (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__S (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__S (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__12638__S (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__B (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__B (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__B (.DIODE(_05962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__B (.DIODE(_05962_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12649__B (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__B (.DIODE(_05916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__B (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12655__B (.DIODE(_05854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12659__B (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__B (.DIODE(_05791_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__B (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12665__B (.DIODE(_05649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12669__B (.DIODE(_05706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__B (.DIODE(_05706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__B (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__B (.DIODE(_05588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__B (.DIODE(_05523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12680__B (.DIODE(_05523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12684__B (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__B (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12688__B (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__B (.DIODE(_05219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12695__B (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12696__B (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__B (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12702__B (.DIODE(_05143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__B (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12708__B (.DIODE(_04991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12713__B (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__B (.DIODE(_04904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12719__B (.DIODE(_05067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__A2 (.DIODE(_05067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12733__A2_N (.DIODE(_00200_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__B (.DIODE(_00201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12761__B2 (.DIODE(_00232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12771__A2 (.DIODE(_00234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__B (.DIODE(_00449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12795__A (.DIODE(_04531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__A (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12803__B (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__12807__A1 (.DIODE(_02078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__12809__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__12811__A1 (.DIODE(_00240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12811__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__12812__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__A1 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__12813__C1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12814__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__12815__A1 (.DIODE(_00258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12815__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__12815__C1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12816__B (.DIODE(_05944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12817__A1 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12817__A2 (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12817__C1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12818__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__A1 (.DIODE(_00213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__12819__C1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12820__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__12821__A1 (.DIODE(_00374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12821__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__12821__C1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12822__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__12823__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__12823__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__12823__C1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12824__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__12825__A1 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12825__C1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__12826__B (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__12827__A1 (.DIODE(_00330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12827__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__12827__C1 (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__12828__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__12829__A1 (.DIODE(_00324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12830__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12831__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12832__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__A1 (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12833__C1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__12834__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__A1 (.DIODE(_00366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12836__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12837__A1 (.DIODE(_00361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12837__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__A1 (.DIODE(_00354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12839__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12841__A1 (.DIODE(_00348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12841__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__A1 (.DIODE(_00189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12843__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12845__A1 (.DIODE(_00179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12845__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12847__A1 (.DIODE(_00172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12847__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12847__C1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12849__A1 (.DIODE(_00163_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12849__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12850__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12851__A1 (.DIODE(_06547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12851__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__A1 (.DIODE(_06540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12853__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12855__A1 (.DIODE(_06563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12855__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12856__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__A1 (.DIODE(_06559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12857__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12859__A1 (.DIODE(_06525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12860__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12861__A1 (.DIODE(_06517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12861__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12862__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__12863__A1 (.DIODE(_00143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12863__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__12864__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__12865__A1 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12866__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__12867__A1 (.DIODE(_00700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12868__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__12869__A1 (.DIODE(_01951_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12870__B (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__12871__A1 (.DIODE(_02066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__B1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__B2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12976__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12977__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12979__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12981__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12982__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12982__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12985__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12987__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12988__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12988__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12989__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12990__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12991__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12993__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12994__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12995__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12996__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__12998__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__12999__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__A2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__13000__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13001__A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13003__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13004__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13005__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13007__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13008__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13009__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13010__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13014__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13015__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__13016__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13016__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13018__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13019__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__13020__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13020__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13021__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13024__B1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__A2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__A2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13028__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13029__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__13035__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__B1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__B2 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__13043__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13044__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__13045__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13047__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__B1 (.DIODE(_06532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13049__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__13053__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__13055__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__13057__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__13057__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__13059__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__13061__A1 (.DIODE(_00342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13061__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__13063__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__A1 (.DIODE(_00339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__A1 (.DIODE(_00357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__13069__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__13069__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__13071__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__13073__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__13074__C1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__13075__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__13077__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__13077__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__13081__A1 (.DIODE(_00216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13082__C1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__13089__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__13091__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__13095__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__13096__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13096__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13098__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13099__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__13100__A2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13101__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__13101__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__13102__C (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13103__A2 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__13104__B1 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13105__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13107__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13109__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13112__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13113__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13113__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13114__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13117__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13118__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13118__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13121__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13122__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13122__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13123__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13125__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13126__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13126__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13127__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13130__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13131__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13131__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13132__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13135__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13136__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13136__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13137__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13140__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13141__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13141__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__13142__A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA__13145__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13146__A2 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13146__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__13147__A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA__13150__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13160__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13161__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13161__B2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13162__A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__13165__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13166__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13166__B2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13170__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13171__B2 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__13175__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13176__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13180__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13181__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13185__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13186__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13190__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13191__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13195__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13196__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13199__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13200__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13204__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13205__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13205__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13208__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__A2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__13209__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13213__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13214__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13214__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13217__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13218__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13222__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13223__A2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__13223__B2 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__13226__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13231__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13240__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13244__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13251__A2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__13252__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13252__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13254__A2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__13254__B2 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__13257__A2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__13257__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__A2 (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__13260__B2 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__13262__B1 (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout101_A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout104_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(_00375_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout10_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(_00329_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(_00325_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(_00313_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout117_A (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(_00286_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(_00276_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout12_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(_00190_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(_00190_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout134_A (.DIODE(_00184_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(_00338_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(_00264_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(_00160_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout14_A (.DIODE(_00699_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(_06542_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout15_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(_05945_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(_05944_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(_05944_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout17_A (.DIODE(_00409_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout18_A (.DIODE(_02079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(_06465_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout19_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(_02241_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(_06534_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout20_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(_06475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_A (.DIODE(_06364_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(_06360_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout21_A (.DIODE(_02079_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout220_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(_06347_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(_06331_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_A (.DIODE(_02078_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_A (.DIODE(_02514_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(_02514_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(_06520_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(_06494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout23_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout248_A (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout251_A (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout25_A (.DIODE(_00327_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout264_A (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout265_A (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_A (.DIODE(_00327_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout27_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(net283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout28_A (.DIODE(_00323_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout29_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout30_A (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout31_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout32_A (.DIODE(_00305_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout33_A (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_A (.DIODE(_00293_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout35_A (.DIODE(_00284_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_A (.DIODE(_00284_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout41_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout43_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_A (.DIODE(_00249_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout49_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(_00217_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout51_A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(_00171_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_A (.DIODE(_06562_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(_06562_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout59_A (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(_06560_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout61_A (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(_06546_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(_06541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(_06541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_A (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout66_A (.DIODE(_06524_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout69_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout72_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(_00365_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(_00362_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout7_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout81_A (.DIODE(_00353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout8_A (.DIODE(_02067_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout91_A (.DIODE(_00245_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap102_A (.DIODE(_00179_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap113_A (.DIODE(_00314_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap118_A (.DIODE(_00287_));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap9_A (.DIODE(_02066_));
 sky130_fd_sc_hd__fill_2 FILLER_0_0_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_728 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_628 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_756 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_403 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_710 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_638 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_308 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_22 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_695 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_535 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_543 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_89 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _06571_ (.A(net591),
    .Y(_04400_));
 sky130_fd_sc_hd__inv_2 _06572_ (.A(net300),
    .Y(_04411_));
 sky130_fd_sc_hd__inv_2 _06573_ (.A(net351),
    .Y(_04422_));
 sky130_fd_sc_hd__inv_2 _06574_ (.A(net337),
    .Y(_04433_));
 sky130_fd_sc_hd__inv_2 _06575_ (.A(net333),
    .Y(_04444_));
 sky130_fd_sc_hd__inv_2 _06576_ (.A(\div_shifter[2] ),
    .Y(_04454_));
 sky130_fd_sc_hd__inv_2 _06577_ (.A(net255),
    .Y(_04465_));
 sky130_fd_sc_hd__inv_2 _06578_ (.A(instruction[3]),
    .Y(_04476_));
 sky130_fd_sc_hd__inv_2 _06579_ (.A(instruction[6]),
    .Y(_04487_));
 sky130_fd_sc_hd__clkinv_4 _06580_ (.A(instruction[5]),
    .Y(_04498_));
 sky130_fd_sc_hd__inv_2 _06581_ (.A(net292),
    .Y(_04509_));
 sky130_fd_sc_hd__inv_2 _06582_ (.A(instruction[41]),
    .Y(_04520_));
 sky130_fd_sc_hd__clkinv_4 _06583_ (.A(reg1_val[31]),
    .Y(_04531_));
 sky130_fd_sc_hd__inv_2 _06584_ (.A(net294),
    .Y(_04542_));
 sky130_fd_sc_hd__inv_2 _06585_ (.A(rst),
    .Y(_04553_));
 sky130_fd_sc_hd__nand2_1 _06586_ (.A(instruction[0]),
    .B(pred_val),
    .Y(_04563_));
 sky130_fd_sc_hd__and2_1 _06587_ (.A(pred_val),
    .B(instruction[1]),
    .X(_04574_));
 sky130_fd_sc_hd__o31a_1 _06588_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(pred_val),
    .X(_04585_));
 sky130_fd_sc_hd__and4b_4 _06589_ (.A_N(instruction[1]),
    .B(instruction[2]),
    .C(instruction[0]),
    .D(pred_val),
    .X(_04596_));
 sky130_fd_sc_hd__or3b_4 _06590_ (.A(_04574_),
    .B(_04563_),
    .C_N(instruction[2]),
    .X(_04607_));
 sky130_fd_sc_hd__or2_1 _06591_ (.A(instruction[23]),
    .B(_04596_),
    .X(_04618_));
 sky130_fd_sc_hd__o211a_4 _06592_ (.A1(instruction[16]),
    .A2(_04607_),
    .B1(_04618_),
    .C1(net272),
    .X(reg1_idx[5]));
 sky130_fd_sc_hd__or2_1 _06593_ (.A(instruction[20]),
    .B(_04596_),
    .X(_04639_));
 sky130_fd_sc_hd__o211a_4 _06594_ (.A1(instruction[13]),
    .A2(_04607_),
    .B1(_04639_),
    .C1(net272),
    .X(reg1_idx[2]));
 sky130_fd_sc_hd__or2_1 _06595_ (.A(instruction[21]),
    .B(_04596_),
    .X(_04660_));
 sky130_fd_sc_hd__o211a_4 _06596_ (.A1(instruction[14]),
    .A2(_04607_),
    .B1(_04660_),
    .C1(net272),
    .X(reg1_idx[3]));
 sky130_fd_sc_hd__or2_1 _06597_ (.A(instruction[18]),
    .B(_04596_),
    .X(_04680_));
 sky130_fd_sc_hd__o211a_4 _06598_ (.A1(instruction[11]),
    .A2(_04607_),
    .B1(_04680_),
    .C1(net272),
    .X(reg1_idx[0]));
 sky130_fd_sc_hd__or2_1 _06599_ (.A(instruction[19]),
    .B(_04596_),
    .X(_04701_));
 sky130_fd_sc_hd__o211a_4 _06600_ (.A1(instruction[12]),
    .A2(_04607_),
    .B1(_04701_),
    .C1(net272),
    .X(reg1_idx[1]));
 sky130_fd_sc_hd__or2_1 _06601_ (.A(instruction[22]),
    .B(_04596_),
    .X(_04722_));
 sky130_fd_sc_hd__o211a_4 _06602_ (.A1(instruction[15]),
    .A2(_04607_),
    .B1(_04722_),
    .C1(net273),
    .X(reg1_idx[4]));
 sky130_fd_sc_hd__or4bb_4 _06603_ (.A(instruction[0]),
    .B(instruction[1]),
    .C_N(instruction[2]),
    .D_N(pred_val),
    .X(_04743_));
 sky130_fd_sc_hd__nor2_8 _06604_ (.A(instruction[3]),
    .B(_04743_),
    .Y(is_load));
 sky130_fd_sc_hd__nor2_8 _06605_ (.A(_04476_),
    .B(_04743_),
    .Y(is_store));
 sky130_fd_sc_hd__and4bb_1 _06606_ (.A_N(instruction[0]),
    .B_N(instruction[2]),
    .C(instruction[1]),
    .D(pred_val),
    .X(_04773_));
 sky130_fd_sc_hd__or4bb_1 _06607_ (.A(instruction[0]),
    .B(instruction[2]),
    .C_N(instruction[1]),
    .D_N(pred_val),
    .X(_04784_));
 sky130_fd_sc_hd__o311a_4 _06608_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[41]),
    .C1(pred_val),
    .X(_04795_));
 sky130_fd_sc_hd__and4bb_2 _06609_ (.A_N(instruction[1]),
    .B_N(instruction[2]),
    .C(instruction[0]),
    .D(pred_val),
    .X(_04806_));
 sky130_fd_sc_hd__or4bb_4 _06610_ (.A(instruction[1]),
    .B(instruction[2]),
    .C_N(instruction[0]),
    .D_N(pred_val),
    .X(_04817_));
 sky130_fd_sc_hd__and2_4 _06611_ (.A(instruction[25]),
    .B(net273),
    .X(_04828_));
 sky130_fd_sc_hd__o211a_1 _06612_ (.A1(instruction[1]),
    .A2(instruction[2]),
    .B1(instruction[25]),
    .C1(pred_val),
    .X(_04839_));
 sky130_fd_sc_hd__o211ai_1 _06613_ (.A1(instruction[1]),
    .A2(instruction[2]),
    .B1(instruction[25]),
    .C1(pred_val),
    .Y(_04850_));
 sky130_fd_sc_hd__a21o_1 _06614_ (.A1(instruction[41]),
    .A2(_04806_),
    .B1(_04839_),
    .X(_04860_));
 sky130_fd_sc_hd__a21oi_4 _06615_ (.A1(instruction[41]),
    .A2(_04806_),
    .B1(_04839_),
    .Y(_04871_));
 sky130_fd_sc_hd__a221o_1 _06616_ (.A1(instruction[24]),
    .A2(_04795_),
    .B1(_04806_),
    .B2(instruction[41]),
    .C1(_04839_),
    .X(_04882_));
 sky130_fd_sc_hd__nand2_1 _06617_ (.A(net271),
    .B(_04882_),
    .Y(_04893_));
 sky130_fd_sc_hd__and2_4 _06618_ (.A(instruction[39]),
    .B(net273),
    .X(_04904_));
 sky130_fd_sc_hd__nor2_1 _06619_ (.A(net252),
    .B(_04904_),
    .Y(_04915_));
 sky130_fd_sc_hd__o2bb2a_1 _06620_ (.A1_N(reg2_val[29]),
    .A2_N(net267),
    .B1(net230),
    .B2(_04915_),
    .X(_04926_));
 sky130_fd_sc_hd__a2bb2o_2 _06621_ (.A1_N(_04915_),
    .A2_N(net230),
    .B1(net267),
    .B2(reg2_val[29]),
    .X(_04937_));
 sky130_fd_sc_hd__and2_1 _06622_ (.A(reg1_val[29]),
    .B(_04937_),
    .X(_04948_));
 sky130_fd_sc_hd__or2_1 _06623_ (.A(reg1_val[29]),
    .B(_04937_),
    .X(_04958_));
 sky130_fd_sc_hd__and2b_1 _06624_ (.A_N(_04948_),
    .B(_04958_),
    .X(_04969_));
 sky130_fd_sc_hd__inv_2 _06625_ (.A(_04969_),
    .Y(_04980_));
 sky130_fd_sc_hd__and2_4 _06626_ (.A(instruction[38]),
    .B(net273),
    .X(_04991_));
 sky130_fd_sc_hd__nor2_1 _06627_ (.A(net252),
    .B(_04991_),
    .Y(_05002_));
 sky130_fd_sc_hd__o2bb2a_1 _06628_ (.A1_N(reg2_val[28]),
    .A2_N(net267),
    .B1(net230),
    .B2(_05002_),
    .X(_05013_));
 sky130_fd_sc_hd__a2bb2o_4 _06629_ (.A1_N(_05002_),
    .A2_N(net230),
    .B1(net267),
    .B2(reg2_val[28]),
    .X(_05024_));
 sky130_fd_sc_hd__and2_1 _06630_ (.A(reg1_val[28]),
    .B(_05024_),
    .X(_05035_));
 sky130_fd_sc_hd__or2_1 _06631_ (.A(reg1_val[28]),
    .B(_05024_),
    .X(_05045_));
 sky130_fd_sc_hd__and2b_1 _06632_ (.A_N(_05035_),
    .B(_05045_),
    .X(_05056_));
 sky130_fd_sc_hd__and2_4 _06633_ (.A(instruction[40]),
    .B(net273),
    .X(_05067_));
 sky130_fd_sc_hd__nor2_1 _06634_ (.A(_04871_),
    .B(_05067_),
    .Y(_05078_));
 sky130_fd_sc_hd__o2bb2a_1 _06635_ (.A1_N(reg2_val[30]),
    .A2_N(net268),
    .B1(net230),
    .B2(_05078_),
    .X(_05089_));
 sky130_fd_sc_hd__a2bb2o_4 _06636_ (.A1_N(_05078_),
    .A2_N(net230),
    .B1(net268),
    .B2(reg2_val[30]),
    .X(_05100_));
 sky130_fd_sc_hd__and2_1 _06637_ (.A(reg1_val[30]),
    .B(_05100_),
    .X(_05111_));
 sky130_fd_sc_hd__nor2_1 _06638_ (.A(reg1_val[30]),
    .B(_05100_),
    .Y(_05122_));
 sky130_fd_sc_hd__or2_2 _06639_ (.A(_05111_),
    .B(_05122_),
    .X(_05133_));
 sky130_fd_sc_hd__and2_4 _06640_ (.A(instruction[37]),
    .B(net273),
    .X(_05143_));
 sky130_fd_sc_hd__nor2_1 _06641_ (.A(_04871_),
    .B(_05143_),
    .Y(_05154_));
 sky130_fd_sc_hd__o2bb2a_2 _06642_ (.A1_N(reg2_val[27]),
    .A2_N(net267),
    .B1(net231),
    .B2(_05154_),
    .X(_05165_));
 sky130_fd_sc_hd__and2b_1 _06643_ (.A_N(reg1_val[27]),
    .B(_05165_),
    .X(_05176_));
 sky130_fd_sc_hd__nand2b_2 _06644_ (.A_N(_05165_),
    .B(reg1_val[27]),
    .Y(_05187_));
 sky130_fd_sc_hd__nand2b_2 _06645_ (.A_N(_05176_),
    .B(_05187_),
    .Y(_05198_));
 sky130_fd_sc_hd__nand2_1 _06646_ (.A(_05133_),
    .B(_05198_),
    .Y(_05209_));
 sky130_fd_sc_hd__and2_4 _06647_ (.A(instruction[35]),
    .B(net273),
    .X(_05219_));
 sky130_fd_sc_hd__nor2_1 _06648_ (.A(net252),
    .B(_05219_),
    .Y(_05230_));
 sky130_fd_sc_hd__o2bb2a_4 _06649_ (.A1_N(reg2_val[25]),
    .A2_N(net267),
    .B1(net231),
    .B2(_05230_),
    .X(_05241_));
 sky130_fd_sc_hd__and2b_1 _06650_ (.A_N(_05241_),
    .B(reg1_val[25]),
    .X(_05252_));
 sky130_fd_sc_hd__and2b_1 _06651_ (.A_N(reg1_val[25]),
    .B(_05241_),
    .X(_05263_));
 sky130_fd_sc_hd__or2_2 _06652_ (.A(_05252_),
    .B(_05263_),
    .X(_05274_));
 sky130_fd_sc_hd__and2_4 _06653_ (.A(instruction[34]),
    .B(net273),
    .X(_05285_));
 sky130_fd_sc_hd__nor2_1 _06654_ (.A(net252),
    .B(_05285_),
    .Y(_05295_));
 sky130_fd_sc_hd__o2bb2a_2 _06655_ (.A1_N(reg2_val[24]),
    .A2_N(net268),
    .B1(net231),
    .B2(_05295_),
    .X(_05306_));
 sky130_fd_sc_hd__a2bb2o_1 _06656_ (.A1_N(_05295_),
    .A2_N(net231),
    .B1(net268),
    .B2(reg2_val[24]),
    .X(_05317_));
 sky130_fd_sc_hd__nand2_1 _06657_ (.A(reg1_val[24]),
    .B(_05317_),
    .Y(_05328_));
 sky130_fd_sc_hd__or2_1 _06658_ (.A(reg1_val[24]),
    .B(_05317_),
    .X(_05339_));
 sky130_fd_sc_hd__nand2_2 _06659_ (.A(_05328_),
    .B(_05339_),
    .Y(_05350_));
 sky130_fd_sc_hd__and2_1 _06660_ (.A(reg2_val[31]),
    .B(net268),
    .X(_05361_));
 sky130_fd_sc_hd__o21ba_1 _06661_ (.A1(_04520_),
    .A2(net231),
    .B1_N(_05361_),
    .X(_05371_));
 sky130_fd_sc_hd__a31o_4 _06662_ (.A1(instruction[41]),
    .A2(net271),
    .A3(_04882_),
    .B1(_05361_),
    .X(_05382_));
 sky130_fd_sc_hd__xnor2_2 _06663_ (.A(_04531_),
    .B(_05382_),
    .Y(_05393_));
 sky130_fd_sc_hd__xnor2_2 _06664_ (.A(reg1_val[31]),
    .B(_05382_),
    .Y(_05404_));
 sky130_fd_sc_hd__and2_4 _06665_ (.A(instruction[36]),
    .B(net273),
    .X(_05415_));
 sky130_fd_sc_hd__nor2_1 _06666_ (.A(net252),
    .B(_05415_),
    .Y(_05426_));
 sky130_fd_sc_hd__o2bb2a_4 _06667_ (.A1_N(reg2_val[26]),
    .A2_N(net267),
    .B1(net231),
    .B2(_05426_),
    .X(_05436_));
 sky130_fd_sc_hd__and2b_1 _06668_ (.A_N(_05436_),
    .B(reg1_val[26]),
    .X(_05447_));
 sky130_fd_sc_hd__inv_2 _06669_ (.A(_05447_),
    .Y(_05458_));
 sky130_fd_sc_hd__and2b_1 _06670_ (.A_N(reg1_val[26]),
    .B(_05436_),
    .X(_05469_));
 sky130_fd_sc_hd__or2_2 _06671_ (.A(_05447_),
    .B(_05469_),
    .X(_05480_));
 sky130_fd_sc_hd__and4_1 _06672_ (.A(_05274_),
    .B(_05350_),
    .C(_05404_),
    .D(_05480_),
    .X(_05490_));
 sky130_fd_sc_hd__or4b_1 _06673_ (.A(_04969_),
    .B(_05056_),
    .C(_05209_),
    .D_N(_05490_),
    .X(_05501_));
 sky130_fd_sc_hd__inv_2 _06674_ (.A(_05501_),
    .Y(_05512_));
 sky130_fd_sc_hd__and2_4 _06675_ (.A(instruction[33]),
    .B(net273),
    .X(_05523_));
 sky130_fd_sc_hd__nor2_1 _06676_ (.A(net252),
    .B(_05523_),
    .Y(_05534_));
 sky130_fd_sc_hd__o2bb2a_4 _06677_ (.A1_N(reg2_val[23]),
    .A2_N(net267),
    .B1(net231),
    .B2(_05534_),
    .X(_05544_));
 sky130_fd_sc_hd__and2b_1 _06678_ (.A_N(_05544_),
    .B(reg1_val[23]),
    .X(_05555_));
 sky130_fd_sc_hd__and2b_1 _06679_ (.A_N(reg1_val[23]),
    .B(_05544_),
    .X(_05566_));
 sky130_fd_sc_hd__nor2_1 _06680_ (.A(_05555_),
    .B(_05566_),
    .Y(_05577_));
 sky130_fd_sc_hd__and2_4 _06681_ (.A(instruction[32]),
    .B(net272),
    .X(_05588_));
 sky130_fd_sc_hd__nor2_1 _06682_ (.A(net252),
    .B(_05588_),
    .Y(_05598_));
 sky130_fd_sc_hd__o2bb2a_4 _06683_ (.A1_N(reg2_val[22]),
    .A2_N(net269),
    .B1(net230),
    .B2(_05598_),
    .X(_05609_));
 sky130_fd_sc_hd__and2b_1 _06684_ (.A_N(_05609_),
    .B(reg1_val[22]),
    .X(_05620_));
 sky130_fd_sc_hd__and2b_1 _06685_ (.A_N(reg1_val[22]),
    .B(_05609_),
    .X(_05629_));
 sky130_fd_sc_hd__nor2_2 _06686_ (.A(_05620_),
    .B(_05629_),
    .Y(_05639_));
 sky130_fd_sc_hd__and2_4 _06687_ (.A(instruction[30]),
    .B(net272),
    .X(_05649_));
 sky130_fd_sc_hd__nor2_1 _06688_ (.A(_04871_),
    .B(_05649_),
    .Y(_05658_));
 sky130_fd_sc_hd__o2bb2a_4 _06689_ (.A1_N(reg2_val[20]),
    .A2_N(net269),
    .B1(net230),
    .B2(_05658_),
    .X(_05668_));
 sky130_fd_sc_hd__nand2b_1 _06690_ (.A_N(_05668_),
    .B(reg1_val[20]),
    .Y(_05677_));
 sky130_fd_sc_hd__and2b_1 _06691_ (.A_N(reg1_val[20]),
    .B(_05668_),
    .X(_05687_));
 sky130_fd_sc_hd__xnor2_2 _06692_ (.A(reg1_val[20]),
    .B(_05668_),
    .Y(_05696_));
 sky130_fd_sc_hd__o311a_4 _06693_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[31]),
    .C1(pred_val),
    .X(_05706_));
 sky130_fd_sc_hd__nor2_1 _06694_ (.A(_04871_),
    .B(_05706_),
    .Y(_05716_));
 sky130_fd_sc_hd__o2bb2a_2 _06695_ (.A1_N(reg2_val[21]),
    .A2_N(net267),
    .B1(net230),
    .B2(_05716_),
    .X(_05725_));
 sky130_fd_sc_hd__a2bb2o_2 _06696_ (.A1_N(_05716_),
    .A2_N(net230),
    .B1(net267),
    .B2(reg2_val[21]),
    .X(_05734_));
 sky130_fd_sc_hd__nand2_1 _06697_ (.A(reg1_val[21]),
    .B(_05734_),
    .Y(_05744_));
 sky130_fd_sc_hd__nor2_1 _06698_ (.A(reg1_val[21]),
    .B(_05734_),
    .Y(_05753_));
 sky130_fd_sc_hd__xnor2_2 _06699_ (.A(reg1_val[21]),
    .B(_05725_),
    .Y(_05763_));
 sky130_fd_sc_hd__nor4_1 _06700_ (.A(_05577_),
    .B(_05639_),
    .C(_05696_),
    .D(_05763_),
    .Y(_05773_));
 sky130_fd_sc_hd__inv_2 _06701_ (.A(_05773_),
    .Y(_05782_));
 sky130_fd_sc_hd__and2_4 _06702_ (.A(instruction[29]),
    .B(net272),
    .X(_05791_));
 sky130_fd_sc_hd__nor2_1 _06703_ (.A(_04871_),
    .B(_05791_),
    .Y(_05799_));
 sky130_fd_sc_hd__o2bb2a_4 _06704_ (.A1_N(reg2_val[19]),
    .A2_N(net267),
    .B1(net230),
    .B2(_05799_),
    .X(_05808_));
 sky130_fd_sc_hd__and2b_1 _06705_ (.A_N(_05808_),
    .B(reg1_val[19]),
    .X(_05817_));
 sky130_fd_sc_hd__and2b_1 _06706_ (.A_N(reg1_val[19]),
    .B(_05808_),
    .X(_05826_));
 sky130_fd_sc_hd__nor2_1 _06707_ (.A(_05817_),
    .B(_05826_),
    .Y(_05835_));
 sky130_fd_sc_hd__inv_2 _06708_ (.A(_05835_),
    .Y(_05845_));
 sky130_fd_sc_hd__and2_4 _06709_ (.A(instruction[28]),
    .B(net272),
    .X(_05854_));
 sky130_fd_sc_hd__nor2_1 _06710_ (.A(net252),
    .B(_05854_),
    .Y(_05863_));
 sky130_fd_sc_hd__o2bb2a_4 _06711_ (.A1_N(reg2_val[18]),
    .A2_N(net268),
    .B1(net230),
    .B2(_05863_),
    .X(_05872_));
 sky130_fd_sc_hd__a2bb2o_2 _06712_ (.A1_N(_05863_),
    .A2_N(net230),
    .B1(net268),
    .B2(reg2_val[18]),
    .X(_05881_));
 sky130_fd_sc_hd__and2_1 _06713_ (.A(reg1_val[18]),
    .B(_05881_),
    .X(_05889_));
 sky130_fd_sc_hd__nor2_1 _06714_ (.A(reg1_val[18]),
    .B(_05881_),
    .Y(_05898_));
 sky130_fd_sc_hd__or2_2 _06715_ (.A(_05889_),
    .B(_05898_),
    .X(_05907_));
 sky130_fd_sc_hd__and2_4 _06716_ (.A(instruction[27]),
    .B(net272),
    .X(_05916_));
 sky130_fd_sc_hd__nor2_1 _06717_ (.A(net252),
    .B(_05916_),
    .Y(_05925_));
 sky130_fd_sc_hd__o2bb2a_4 _06718_ (.A1_N(reg2_val[17]),
    .A2_N(net267),
    .B1(net230),
    .B2(_05925_),
    .X(_05934_));
 sky130_fd_sc_hd__and2b_1 _06719_ (.A_N(_05934_),
    .B(reg1_val[17]),
    .X(_05943_));
 sky130_fd_sc_hd__nand2b_1 _06720_ (.A_N(reg1_val[17]),
    .B(_05934_),
    .Y(_05950_));
 sky130_fd_sc_hd__nand2b_1 _06721_ (.A_N(_05943_),
    .B(_05950_),
    .Y(_05956_));
 sky130_fd_sc_hd__o311a_4 _06722_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[26]),
    .C1(pred_val),
    .X(_05962_));
 sky130_fd_sc_hd__nor2_1 _06723_ (.A(net252),
    .B(_05962_),
    .Y(_05968_));
 sky130_fd_sc_hd__o2bb2a_2 _06724_ (.A1_N(reg2_val[16]),
    .A2_N(net268),
    .B1(net230),
    .B2(_05968_),
    .X(_05974_));
 sky130_fd_sc_hd__a2bb2o_2 _06725_ (.A1_N(_05968_),
    .A2_N(net230),
    .B1(net268),
    .B2(reg2_val[16]),
    .X(_05980_));
 sky130_fd_sc_hd__and2_1 _06726_ (.A(reg1_val[16]),
    .B(_05980_),
    .X(_05987_));
 sky130_fd_sc_hd__or2_1 _06727_ (.A(reg1_val[16]),
    .B(_05980_),
    .X(_05998_));
 sky130_fd_sc_hd__and2b_1 _06728_ (.A_N(_05987_),
    .B(_05998_),
    .X(_06009_));
 sky130_fd_sc_hd__and2_1 _06729_ (.A(reg2_val[15]),
    .B(net269),
    .X(_06020_));
 sky130_fd_sc_hd__a31o_4 _06730_ (.A1(net270),
    .A2(_04795_),
    .A3(net251),
    .B1(_06020_),
    .X(_06031_));
 sky130_fd_sc_hd__and2_1 _06731_ (.A(net290),
    .B(_06031_),
    .X(_06042_));
 sky130_fd_sc_hd__nor2_1 _06732_ (.A(net290),
    .B(_06031_),
    .Y(_06053_));
 sky130_fd_sc_hd__nor2_2 _06733_ (.A(_06042_),
    .B(_06053_),
    .Y(_06064_));
 sky130_fd_sc_hd__and2_1 _06734_ (.A(reg2_val[14]),
    .B(net269),
    .X(_06075_));
 sky130_fd_sc_hd__a31o_4 _06735_ (.A1(net270),
    .A2(net252),
    .A3(_05067_),
    .B1(_06075_),
    .X(_06086_));
 sky130_fd_sc_hd__nor2_1 _06736_ (.A(net291),
    .B(_06086_),
    .Y(_06097_));
 sky130_fd_sc_hd__and2_1 _06737_ (.A(net291),
    .B(_06086_),
    .X(_06103_));
 sky130_fd_sc_hd__nor2_1 _06738_ (.A(_06097_),
    .B(_06103_),
    .Y(_06109_));
 sky130_fd_sc_hd__and2_1 _06739_ (.A(reg2_val[13]),
    .B(net269),
    .X(_06115_));
 sky130_fd_sc_hd__a31o_4 _06740_ (.A1(net271),
    .A2(net251),
    .A3(_04904_),
    .B1(_06115_),
    .X(_06121_));
 sky130_fd_sc_hd__and2_1 _06741_ (.A(reg1_val[13]),
    .B(_06121_),
    .X(_06127_));
 sky130_fd_sc_hd__nor2_1 _06742_ (.A(reg1_val[13]),
    .B(_06121_),
    .Y(_06133_));
 sky130_fd_sc_hd__or2_2 _06743_ (.A(_06127_),
    .B(_06133_),
    .X(_06139_));
 sky130_fd_sc_hd__and2_1 _06744_ (.A(reg2_val[12]),
    .B(net269),
    .X(_06145_));
 sky130_fd_sc_hd__a31o_4 _06745_ (.A1(net271),
    .A2(net252),
    .A3(_04991_),
    .B1(_06145_),
    .X(_06151_));
 sky130_fd_sc_hd__and2_1 _06746_ (.A(reg1_val[12]),
    .B(_06151_),
    .X(_06157_));
 sky130_fd_sc_hd__nor2_1 _06747_ (.A(reg1_val[12]),
    .B(_06151_),
    .Y(_06163_));
 sky130_fd_sc_hd__or2_2 _06748_ (.A(_06157_),
    .B(_06163_),
    .X(_06169_));
 sky130_fd_sc_hd__and2_1 _06749_ (.A(reg2_val[11]),
    .B(net269),
    .X(_06176_));
 sky130_fd_sc_hd__a31o_4 _06750_ (.A1(net270),
    .A2(net252),
    .A3(_05143_),
    .B1(_06176_),
    .X(_06185_));
 sky130_fd_sc_hd__and2_1 _06751_ (.A(reg1_val[11]),
    .B(_06185_),
    .X(_06193_));
 sky130_fd_sc_hd__nor2_1 _06752_ (.A(reg1_val[11]),
    .B(_06185_),
    .Y(_06202_));
 sky130_fd_sc_hd__nor2_1 _06753_ (.A(_06193_),
    .B(_06202_),
    .Y(_06211_));
 sky130_fd_sc_hd__or2_1 _06754_ (.A(_06193_),
    .B(_06202_),
    .X(_06220_));
 sky130_fd_sc_hd__and2_1 _06755_ (.A(reg2_val[10]),
    .B(net267),
    .X(_06229_));
 sky130_fd_sc_hd__a31o_4 _06756_ (.A1(net271),
    .A2(net252),
    .A3(_05415_),
    .B1(_06229_),
    .X(_06238_));
 sky130_fd_sc_hd__nor2_1 _06757_ (.A(reg1_val[10]),
    .B(_06238_),
    .Y(_06247_));
 sky130_fd_sc_hd__and2_1 _06758_ (.A(reg1_val[10]),
    .B(_06238_),
    .X(_06256_));
 sky130_fd_sc_hd__nor2_1 _06759_ (.A(_06247_),
    .B(_06256_),
    .Y(_06265_));
 sky130_fd_sc_hd__and2_2 _06760_ (.A(reg2_val[9]),
    .B(net269),
    .X(_06274_));
 sky130_fd_sc_hd__a31o_4 _06761_ (.A1(net270),
    .A2(net251),
    .A3(_05219_),
    .B1(_06274_),
    .X(_06283_));
 sky130_fd_sc_hd__inv_2 _06762_ (.A(_06283_),
    .Y(_06291_));
 sky130_fd_sc_hd__nor2_1 _06763_ (.A(reg1_val[9]),
    .B(_06283_),
    .Y(_06300_));
 sky130_fd_sc_hd__nand2_1 _06764_ (.A(reg1_val[9]),
    .B(_06283_),
    .Y(_06307_));
 sky130_fd_sc_hd__nand2b_1 _06765_ (.A_N(_06300_),
    .B(_06307_),
    .Y(_06313_));
 sky130_fd_sc_hd__and2_1 _06766_ (.A(reg2_val[8]),
    .B(net267),
    .X(_06314_));
 sky130_fd_sc_hd__a31o_4 _06767_ (.A1(net270),
    .A2(net251),
    .A3(_05285_),
    .B1(_06314_),
    .X(_06315_));
 sky130_fd_sc_hd__nor2_1 _06768_ (.A(reg1_val[8]),
    .B(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__nand2_1 _06769_ (.A(reg1_val[8]),
    .B(_06315_),
    .Y(_06317_));
 sky130_fd_sc_hd__nand2b_1 _06770_ (.A_N(_06316_),
    .B(_06317_),
    .Y(_06318_));
 sky130_fd_sc_hd__and2_2 _06771_ (.A(reg2_val[7]),
    .B(net269),
    .X(_06319_));
 sky130_fd_sc_hd__a31o_4 _06772_ (.A1(net270),
    .A2(net251),
    .A3(_05523_),
    .B1(_06319_),
    .X(_06320_));
 sky130_fd_sc_hd__nor2_1 _06773_ (.A(reg1_val[7]),
    .B(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__nand2_1 _06774_ (.A(reg1_val[7]),
    .B(_06320_),
    .Y(_06322_));
 sky130_fd_sc_hd__nand2b_2 _06775_ (.A_N(_06321_),
    .B(_06322_),
    .Y(_06323_));
 sky130_fd_sc_hd__and2_1 _06776_ (.A(reg2_val[6]),
    .B(net269),
    .X(_06324_));
 sky130_fd_sc_hd__a31o_4 _06777_ (.A1(net270),
    .A2(net251),
    .A3(_05588_),
    .B1(_06324_),
    .X(_06325_));
 sky130_fd_sc_hd__or2_1 _06778_ (.A(reg1_val[6]),
    .B(_06325_),
    .X(_06326_));
 sky130_fd_sc_hd__and2_1 _06779_ (.A(reg1_val[6]),
    .B(_06325_),
    .X(_06327_));
 sky130_fd_sc_hd__nand2_1 _06780_ (.A(reg1_val[6]),
    .B(_06325_),
    .Y(_06328_));
 sky130_fd_sc_hd__and2_1 _06781_ (.A(_06326_),
    .B(_06328_),
    .X(_06329_));
 sky130_fd_sc_hd__o2111a_2 _06782_ (.A1(_04520_),
    .A2(_04817_),
    .B1(_04850_),
    .C1(_05706_),
    .D1(net271),
    .X(_06330_));
 sky130_fd_sc_hd__or3b_4 _06783_ (.A(net268),
    .B(_04860_),
    .C_N(_05706_),
    .X(_06331_));
 sky130_fd_sc_hd__a21oi_2 _06784_ (.A1(reg2_val[5]),
    .A2(net268),
    .B1(net250),
    .Y(_06332_));
 sky130_fd_sc_hd__a21o_2 _06785_ (.A1(reg2_val[5]),
    .A2(net268),
    .B1(net250),
    .X(_06333_));
 sky130_fd_sc_hd__nor2_1 _06786_ (.A(reg1_val[5]),
    .B(_06333_),
    .Y(_06334_));
 sky130_fd_sc_hd__and2_1 _06787_ (.A(reg1_val[5]),
    .B(_06333_),
    .X(_06335_));
 sky130_fd_sc_hd__nand2_1 _06788_ (.A(reg1_val[5]),
    .B(_06333_),
    .Y(_06336_));
 sky130_fd_sc_hd__nor2_1 _06789_ (.A(_06334_),
    .B(_06335_),
    .Y(_06337_));
 sky130_fd_sc_hd__or2_1 _06790_ (.A(_06334_),
    .B(_06335_),
    .X(_06338_));
 sky130_fd_sc_hd__and2_2 _06791_ (.A(reg2_val[4]),
    .B(net269),
    .X(_06339_));
 sky130_fd_sc_hd__a31o_1 _06792_ (.A1(net270),
    .A2(net251),
    .A3(_05649_),
    .B1(_06339_),
    .X(_06340_));
 sky130_fd_sc_hd__a31oi_2 _06793_ (.A1(net270),
    .A2(net251),
    .A3(_05649_),
    .B1(_06339_),
    .Y(_06341_));
 sky130_fd_sc_hd__or2_1 _06794_ (.A(reg1_val[4]),
    .B(net228),
    .X(_06342_));
 sky130_fd_sc_hd__nand2_1 _06795_ (.A(reg1_val[4]),
    .B(net228),
    .Y(_06343_));
 sky130_fd_sc_hd__nand2_2 _06796_ (.A(_06342_),
    .B(_06343_),
    .Y(_06344_));
 sky130_fd_sc_hd__and2_2 _06797_ (.A(reg2_val[3]),
    .B(net269),
    .X(_06345_));
 sky130_fd_sc_hd__a31oi_4 _06798_ (.A1(net270),
    .A2(net251),
    .A3(_05791_),
    .B1(_06345_),
    .Y(_06346_));
 sky130_fd_sc_hd__a31o_4 _06799_ (.A1(net270),
    .A2(net251),
    .A3(_05791_),
    .B1(_06345_),
    .X(_06347_));
 sky130_fd_sc_hd__nor2_1 _06800_ (.A(reg1_val[3]),
    .B(_06347_),
    .Y(_06348_));
 sky130_fd_sc_hd__nand2_1 _06801_ (.A(reg1_val[3]),
    .B(_06347_),
    .Y(_06349_));
 sky130_fd_sc_hd__nand2b_1 _06802_ (.A_N(_06348_),
    .B(_06349_),
    .Y(_06350_));
 sky130_fd_sc_hd__and2_2 _06803_ (.A(reg2_val[2]),
    .B(net269),
    .X(_06351_));
 sky130_fd_sc_hd__a31oi_4 _06804_ (.A1(net270),
    .A2(net251),
    .A3(_05854_),
    .B1(_06351_),
    .Y(_06352_));
 sky130_fd_sc_hd__a31o_1 _06805_ (.A1(net270),
    .A2(net251),
    .A3(_05854_),
    .B1(_06351_),
    .X(_06353_));
 sky130_fd_sc_hd__nand2_1 _06806_ (.A(reg1_val[2]),
    .B(net221),
    .Y(_06354_));
 sky130_fd_sc_hd__nor2_1 _06807_ (.A(reg1_val[2]),
    .B(net221),
    .Y(_06355_));
 sky130_fd_sc_hd__or2_1 _06808_ (.A(reg1_val[2]),
    .B(net221),
    .X(_06356_));
 sky130_fd_sc_hd__nand2_2 _06809_ (.A(_06354_),
    .B(_06356_),
    .Y(_06357_));
 sky130_fd_sc_hd__and2_2 _06810_ (.A(reg2_val[1]),
    .B(net269),
    .X(_06358_));
 sky130_fd_sc_hd__a31oi_4 _06811_ (.A1(net270),
    .A2(net251),
    .A3(_05916_),
    .B1(_06358_),
    .Y(_06359_));
 sky130_fd_sc_hd__a31o_4 _06812_ (.A1(net270),
    .A2(net251),
    .A3(_05916_),
    .B1(_06358_),
    .X(_06360_));
 sky130_fd_sc_hd__or2_1 _06813_ (.A(net289),
    .B(_06360_),
    .X(_06361_));
 sky130_fd_sc_hd__xnor2_2 _06814_ (.A(net289),
    .B(net218),
    .Y(_06362_));
 sky130_fd_sc_hd__and2_1 _06815_ (.A(net270),
    .B(_05962_),
    .X(_06363_));
 sky130_fd_sc_hd__a22oi_4 _06816_ (.A1(reg2_val[0]),
    .A2(net267),
    .B1(net251),
    .B2(_06363_),
    .Y(_06364_));
 sky130_fd_sc_hd__a22o_1 _06817_ (.A1(reg2_val[0]),
    .A2(net267),
    .B1(net251),
    .B2(_06363_),
    .X(_06365_));
 sky130_fd_sc_hd__nand2_1 _06818_ (.A(net287),
    .B(net213),
    .Y(_06366_));
 sky130_fd_sc_hd__and2_1 _06819_ (.A(net289),
    .B(_06359_),
    .X(_06367_));
 sky130_fd_sc_hd__a21o_1 _06820_ (.A1(_06362_),
    .A2(_06366_),
    .B1(_06367_),
    .X(_06368_));
 sky130_fd_sc_hd__and2_1 _06821_ (.A(reg1_val[2]),
    .B(_06352_),
    .X(_06369_));
 sky130_fd_sc_hd__a21o_1 _06822_ (.A1(_06357_),
    .A2(_06368_),
    .B1(_06369_),
    .X(_06370_));
 sky130_fd_sc_hd__and2_1 _06823_ (.A(reg1_val[3]),
    .B(net224),
    .X(_06371_));
 sky130_fd_sc_hd__a21o_1 _06824_ (.A1(_06350_),
    .A2(_06370_),
    .B1(_06371_),
    .X(_06372_));
 sky130_fd_sc_hd__and2_1 _06825_ (.A(reg1_val[4]),
    .B(net225),
    .X(_06373_));
 sky130_fd_sc_hd__a21oi_1 _06826_ (.A1(_06344_),
    .A2(_06372_),
    .B1(_06373_),
    .Y(_06374_));
 sky130_fd_sc_hd__nand2_1 _06827_ (.A(reg1_val[5]),
    .B(_06332_),
    .Y(_06375_));
 sky130_fd_sc_hd__o21a_1 _06828_ (.A1(_06337_),
    .A2(_06374_),
    .B1(_06375_),
    .X(_06376_));
 sky130_fd_sc_hd__nand2b_1 _06829_ (.A_N(_06325_),
    .B(reg1_val[6]),
    .Y(_06377_));
 sky130_fd_sc_hd__o21ai_1 _06830_ (.A1(_06329_),
    .A2(_06376_),
    .B1(_06377_),
    .Y(_06378_));
 sky130_fd_sc_hd__and2b_1 _06831_ (.A_N(_06320_),
    .B(reg1_val[7]),
    .X(_06379_));
 sky130_fd_sc_hd__a21o_1 _06832_ (.A1(_06323_),
    .A2(_06378_),
    .B1(_06379_),
    .X(_06380_));
 sky130_fd_sc_hd__and2b_1 _06833_ (.A_N(_06315_),
    .B(reg1_val[8]),
    .X(_06381_));
 sky130_fd_sc_hd__a21o_1 _06834_ (.A1(_06318_),
    .A2(_06380_),
    .B1(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__and2_1 _06835_ (.A(reg1_val[9]),
    .B(_06291_),
    .X(_06383_));
 sky130_fd_sc_hd__a21oi_1 _06836_ (.A1(_06313_),
    .A2(_06382_),
    .B1(_06383_),
    .Y(_06384_));
 sky130_fd_sc_hd__and2b_1 _06837_ (.A_N(_06238_),
    .B(reg1_val[10]),
    .X(_06385_));
 sky130_fd_sc_hd__o21bai_1 _06838_ (.A1(_06265_),
    .A2(_06384_),
    .B1_N(_06385_),
    .Y(_06386_));
 sky130_fd_sc_hd__and2b_1 _06839_ (.A_N(_06185_),
    .B(reg1_val[11]),
    .X(_06387_));
 sky130_fd_sc_hd__a21o_1 _06840_ (.A1(_06220_),
    .A2(_06386_),
    .B1(_06387_),
    .X(_06388_));
 sky130_fd_sc_hd__and2b_1 _06841_ (.A_N(_06151_),
    .B(reg1_val[12]),
    .X(_06389_));
 sky130_fd_sc_hd__a21o_1 _06842_ (.A1(_06169_),
    .A2(_06388_),
    .B1(_06389_),
    .X(_06390_));
 sky130_fd_sc_hd__and2b_1 _06843_ (.A_N(_06121_),
    .B(reg1_val[13]),
    .X(_06391_));
 sky130_fd_sc_hd__a21oi_1 _06844_ (.A1(_06139_),
    .A2(_06390_),
    .B1(_06391_),
    .Y(_06392_));
 sky130_fd_sc_hd__nand2b_1 _06845_ (.A_N(_06086_),
    .B(net291),
    .Y(_06393_));
 sky130_fd_sc_hd__o21a_1 _06846_ (.A1(_06109_),
    .A2(_06392_),
    .B1(_06393_),
    .X(_06394_));
 sky130_fd_sc_hd__and2b_1 _06847_ (.A_N(_06031_),
    .B(net290),
    .X(_06395_));
 sky130_fd_sc_hd__o21ba_1 _06848_ (.A1(_06064_),
    .A2(_06394_),
    .B1_N(_06395_),
    .X(_06396_));
 sky130_fd_sc_hd__nand2_1 _06849_ (.A(reg1_val[16]),
    .B(_05974_),
    .Y(_06397_));
 sky130_fd_sc_hd__o21ai_1 _06850_ (.A1(_06009_),
    .A2(_06396_),
    .B1(_06397_),
    .Y(_06398_));
 sky130_fd_sc_hd__and2_1 _06851_ (.A(reg1_val[17]),
    .B(_05934_),
    .X(_06399_));
 sky130_fd_sc_hd__a21o_1 _06852_ (.A1(_05956_),
    .A2(_06398_),
    .B1(_06399_),
    .X(_06400_));
 sky130_fd_sc_hd__and2_1 _06853_ (.A(reg1_val[18]),
    .B(_05872_),
    .X(_06401_));
 sky130_fd_sc_hd__a21o_1 _06854_ (.A1(_05907_),
    .A2(_06400_),
    .B1(_06401_),
    .X(_06402_));
 sky130_fd_sc_hd__and2_1 _06855_ (.A(reg1_val[19]),
    .B(_05808_),
    .X(_06403_));
 sky130_fd_sc_hd__a21oi_2 _06856_ (.A1(_05845_),
    .A2(_06402_),
    .B1(_06403_),
    .Y(_06404_));
 sky130_fd_sc_hd__nand2_1 _06857_ (.A(reg1_val[21]),
    .B(_05725_),
    .Y(_06405_));
 sky130_fd_sc_hd__nand2_1 _06858_ (.A(reg1_val[20]),
    .B(_05668_),
    .Y(_06406_));
 sky130_fd_sc_hd__o21a_1 _06859_ (.A1(_05763_),
    .A2(_06406_),
    .B1(_06405_),
    .X(_06407_));
 sky130_fd_sc_hd__or2_1 _06860_ (.A(_05639_),
    .B(_06407_),
    .X(_06408_));
 sky130_fd_sc_hd__nand2_1 _06861_ (.A(reg1_val[22]),
    .B(_05609_),
    .Y(_06409_));
 sky130_fd_sc_hd__a21oi_1 _06862_ (.A1(_06408_),
    .A2(_06409_),
    .B1(_05577_),
    .Y(_06410_));
 sky130_fd_sc_hd__a21oi_1 _06863_ (.A1(reg1_val[23]),
    .A2(_05544_),
    .B1(_06410_),
    .Y(_06411_));
 sky130_fd_sc_hd__o21ai_2 _06864_ (.A1(_05782_),
    .A2(_06404_),
    .B1(_06411_),
    .Y(_06412_));
 sky130_fd_sc_hd__and2_1 _06865_ (.A(reg1_val[30]),
    .B(_05089_),
    .X(_06413_));
 sky130_fd_sc_hd__nand2_1 _06866_ (.A(reg1_val[29]),
    .B(_04926_),
    .Y(_06414_));
 sky130_fd_sc_hd__nand2_1 _06867_ (.A(reg1_val[28]),
    .B(_05013_),
    .Y(_06415_));
 sky130_fd_sc_hd__nand2_1 _06868_ (.A(reg1_val[27]),
    .B(_05165_),
    .Y(_06416_));
 sky130_fd_sc_hd__and2_1 _06869_ (.A(reg1_val[26]),
    .B(_05436_),
    .X(_06417_));
 sky130_fd_sc_hd__and2_1 _06870_ (.A(reg1_val[25]),
    .B(_05241_),
    .X(_06418_));
 sky130_fd_sc_hd__and2_1 _06871_ (.A(reg1_val[24]),
    .B(_05306_),
    .X(_06419_));
 sky130_fd_sc_hd__a21o_1 _06872_ (.A1(_05274_),
    .A2(_06419_),
    .B1(_06418_),
    .X(_06420_));
 sky130_fd_sc_hd__a21o_1 _06873_ (.A1(_05480_),
    .A2(_06420_),
    .B1(_06417_),
    .X(_06421_));
 sky130_fd_sc_hd__nand2_1 _06874_ (.A(_05198_),
    .B(_06421_),
    .Y(_06422_));
 sky130_fd_sc_hd__a21o_1 _06875_ (.A1(_06416_),
    .A2(_06422_),
    .B1(_05056_),
    .X(_06423_));
 sky130_fd_sc_hd__a21o_1 _06876_ (.A1(_06415_),
    .A2(_06423_),
    .B1(_04969_),
    .X(_06424_));
 sky130_fd_sc_hd__nand2_1 _06877_ (.A(_06414_),
    .B(_06424_),
    .Y(_06425_));
 sky130_fd_sc_hd__a21oi_1 _06878_ (.A1(_05133_),
    .A2(_06425_),
    .B1(_06413_),
    .Y(_06426_));
 sky130_fd_sc_hd__or2_1 _06879_ (.A(_04531_),
    .B(_05382_),
    .X(_06427_));
 sky130_fd_sc_hd__a21oi_1 _06880_ (.A1(_05512_),
    .A2(_06412_),
    .B1(instruction[6]),
    .Y(_06428_));
 sky130_fd_sc_hd__o211a_1 _06881_ (.A1(_05393_),
    .A2(_06426_),
    .B1(_06427_),
    .C1(_06428_),
    .X(_06429_));
 sky130_fd_sc_hd__a21o_1 _06882_ (.A1(_05350_),
    .A2(_06412_),
    .B1(_06419_),
    .X(_06430_));
 sky130_fd_sc_hd__a21o_1 _06883_ (.A1(_05274_),
    .A2(_06430_),
    .B1(_06418_),
    .X(_06431_));
 sky130_fd_sc_hd__a21o_1 _06884_ (.A1(_05480_),
    .A2(_06431_),
    .B1(_06417_),
    .X(_06432_));
 sky130_fd_sc_hd__a21boi_1 _06885_ (.A1(_05198_),
    .A2(_06432_),
    .B1_N(_06416_),
    .Y(_06433_));
 sky130_fd_sc_hd__o21ai_1 _06886_ (.A1(_05056_),
    .A2(_06433_),
    .B1(_06415_),
    .Y(_06434_));
 sky130_fd_sc_hd__a21bo_1 _06887_ (.A1(_04980_),
    .A2(_06434_),
    .B1_N(_06414_),
    .X(_06435_));
 sky130_fd_sc_hd__a21o_1 _06888_ (.A1(_05133_),
    .A2(_06435_),
    .B1(_06413_),
    .X(_06436_));
 sky130_fd_sc_hd__o21ai_1 _06889_ (.A1(_05393_),
    .A2(_06436_),
    .B1(_06427_),
    .Y(_06437_));
 sky130_fd_sc_hd__a21o_1 _06890_ (.A1(instruction[6]),
    .A2(_06437_),
    .B1(_06429_),
    .X(_06438_));
 sky130_fd_sc_hd__nor2_1 _06891_ (.A(instruction[3]),
    .B(instruction[4]),
    .Y(_06439_));
 sky130_fd_sc_hd__or2_4 _06892_ (.A(instruction[3]),
    .B(instruction[4]),
    .X(_06440_));
 sky130_fd_sc_hd__nor2_2 _06893_ (.A(net287),
    .B(net216),
    .Y(_06441_));
 sky130_fd_sc_hd__nor2_1 _06894_ (.A(net293),
    .B(net213),
    .Y(_06442_));
 sky130_fd_sc_hd__and3_1 _06895_ (.A(_05845_),
    .B(_05907_),
    .C(_05956_),
    .X(_06443_));
 sky130_fd_sc_hd__and4bb_1 _06896_ (.A_N(_06211_),
    .B_N(_06265_),
    .C(_06313_),
    .D(_06323_),
    .X(_06444_));
 sky130_fd_sc_hd__and4bb_1 _06897_ (.A_N(_06064_),
    .B_N(_06109_),
    .C(_06139_),
    .D(_06169_),
    .X(_06445_));
 sky130_fd_sc_hd__and4b_1 _06898_ (.A_N(_06329_),
    .B(_06338_),
    .C(_06344_),
    .D(_06350_),
    .X(_06446_));
 sky130_fd_sc_hd__o2111a_1 _06899_ (.A1(_06441_),
    .A2(_06442_),
    .B1(_06318_),
    .C1(_06357_),
    .D1(_06362_),
    .X(_06447_));
 sky130_fd_sc_hd__and3_1 _06900_ (.A(_06444_),
    .B(_06445_),
    .C(_06447_),
    .X(_06448_));
 sky130_fd_sc_hd__and4b_1 _06901_ (.A_N(_06009_),
    .B(_06443_),
    .C(_06446_),
    .D(_06448_),
    .X(_06449_));
 sky130_fd_sc_hd__and3_1 _06902_ (.A(_05512_),
    .B(net103),
    .C(_06449_),
    .X(_06450_));
 sky130_fd_sc_hd__nand2_1 _06903_ (.A(instruction[6]),
    .B(_05393_),
    .Y(_06451_));
 sky130_fd_sc_hd__o211a_1 _06904_ (.A1(instruction[6]),
    .A2(_06450_),
    .B1(_06451_),
    .C1(_06439_),
    .X(_06452_));
 sky130_fd_sc_hd__nand2_4 _06905_ (.A(instruction[3]),
    .B(instruction[4]),
    .Y(_06453_));
 sky130_fd_sc_hd__inv_2 _06906_ (.A(_06453_),
    .Y(_06454_));
 sky130_fd_sc_hd__or2_2 _06907_ (.A(_04476_),
    .B(instruction[4]),
    .X(_06455_));
 sky130_fd_sc_hd__a221o_2 _06908_ (.A1(instruction[3]),
    .A2(_06438_),
    .B1(_06450_),
    .B2(_06454_),
    .C1(_06452_),
    .X(_06456_));
 sky130_fd_sc_hd__xnor2_4 _06909_ (.A(_04498_),
    .B(_06456_),
    .Y(dest_pred_val));
 sky130_fd_sc_hd__and3_4 _06910_ (.A(instruction[2]),
    .B(_04563_),
    .C(_04574_),
    .X(_06457_));
 sky130_fd_sc_hd__nand3_1 _06911_ (.A(instruction[2]),
    .B(_04563_),
    .C(_04574_),
    .Y(_06458_));
 sky130_fd_sc_hd__a21o_4 _06912_ (.A1(_04596_),
    .A2(dest_pred_val),
    .B1(_06457_),
    .X(take_branch));
 sky130_fd_sc_hd__and3_1 _06913_ (.A(reg1_idx[0]),
    .B(reg1_idx[1]),
    .C(reg1_idx[4]),
    .X(_06459_));
 sky130_fd_sc_hd__and2_1 _06914_ (.A(reg1_idx[5]),
    .B(_06457_),
    .X(_06460_));
 sky130_fd_sc_hd__and4_4 _06915_ (.A(reg1_idx[2]),
    .B(reg1_idx[3]),
    .C(_06459_),
    .D(_06460_),
    .X(int_return));
 sky130_fd_sc_hd__nand2_8 _06916_ (.A(instruction[6]),
    .B(_04498_),
    .Y(_06461_));
 sky130_fd_sc_hd__a21oi_2 _06917_ (.A1(instruction[6]),
    .A2(instruction[5]),
    .B1(instruction[4]),
    .Y(_06462_));
 sky130_fd_sc_hd__a221oi_4 _06918_ (.A1(net268),
    .A2(_04817_),
    .B1(_06461_),
    .B2(instruction[4]),
    .C1(_06462_),
    .Y(_06463_));
 sky130_fd_sc_hd__a221o_1 _06919_ (.A1(net268),
    .A2(_04817_),
    .B1(_06461_),
    .B2(instruction[4]),
    .C1(_06462_),
    .X(_06464_));
 sky130_fd_sc_hd__nor2_4 _06920_ (.A(net256),
    .B(_06463_),
    .Y(_06465_));
 sky130_fd_sc_hd__nand2_1 _06921_ (.A(net254),
    .B(_06464_),
    .Y(_06466_));
 sky130_fd_sc_hd__nor2_8 _06922_ (.A(div_complete),
    .B(_06465_),
    .Y(busy));
 sky130_fd_sc_hd__and4b_4 _06923_ (.A_N(instruction[2]),
    .B(instruction[1]),
    .C(pred_val),
    .D(instruction[0]),
    .X(_06467_));
 sky130_fd_sc_hd__and2_4 _06924_ (.A(instruction[11]),
    .B(_06467_),
    .X(dest_pred[0]));
 sky130_fd_sc_hd__and2_4 _06925_ (.A(instruction[12]),
    .B(_06467_),
    .X(dest_pred[1]));
 sky130_fd_sc_hd__and2_4 _06926_ (.A(instruction[13]),
    .B(_06467_),
    .X(dest_pred[2]));
 sky130_fd_sc_hd__or3_4 _06927_ (.A(net271),
    .B(_04806_),
    .C(_06457_),
    .X(_06468_));
 sky130_fd_sc_hd__and2_4 _06928_ (.A(instruction[11]),
    .B(_06468_),
    .X(dest_idx[0]));
 sky130_fd_sc_hd__and2_4 _06929_ (.A(instruction[12]),
    .B(_06468_),
    .X(dest_idx[1]));
 sky130_fd_sc_hd__and2_4 _06930_ (.A(instruction[13]),
    .B(_06468_),
    .X(dest_idx[2]));
 sky130_fd_sc_hd__and2_4 _06931_ (.A(instruction[14]),
    .B(_06468_),
    .X(dest_idx[3]));
 sky130_fd_sc_hd__and2_4 _06932_ (.A(instruction[15]),
    .B(_06468_),
    .X(dest_idx[4]));
 sky130_fd_sc_hd__and2_4 _06933_ (.A(instruction[16]),
    .B(_06468_),
    .X(dest_idx[5]));
 sky130_fd_sc_hd__or2_1 _06934_ (.A(instruction[25]),
    .B(_04596_),
    .X(_06469_));
 sky130_fd_sc_hd__o211a_4 _06935_ (.A1(instruction[18]),
    .A2(_04607_),
    .B1(_06469_),
    .C1(net272),
    .X(reg2_idx[0]));
 sky130_fd_sc_hd__or2_1 _06936_ (.A(instruction[26]),
    .B(_04596_),
    .X(_06470_));
 sky130_fd_sc_hd__o211a_4 _06937_ (.A1(instruction[19]),
    .A2(_04607_),
    .B1(_06470_),
    .C1(net272),
    .X(reg2_idx[1]));
 sky130_fd_sc_hd__or2_1 _06938_ (.A(instruction[27]),
    .B(_04596_),
    .X(_06471_));
 sky130_fd_sc_hd__o211a_4 _06939_ (.A1(instruction[20]),
    .A2(_04607_),
    .B1(_06471_),
    .C1(net272),
    .X(reg2_idx[2]));
 sky130_fd_sc_hd__or2_1 _06940_ (.A(instruction[28]),
    .B(_04596_),
    .X(_06472_));
 sky130_fd_sc_hd__o211a_4 _06941_ (.A1(instruction[21]),
    .A2(_04607_),
    .B1(_06472_),
    .C1(net272),
    .X(reg2_idx[3]));
 sky130_fd_sc_hd__or2_1 _06942_ (.A(instruction[29]),
    .B(_04596_),
    .X(_06473_));
 sky130_fd_sc_hd__o211a_4 _06943_ (.A1(instruction[22]),
    .A2(_04607_),
    .B1(_06473_),
    .C1(net272),
    .X(reg2_idx[4]));
 sky130_fd_sc_hd__or2_1 _06944_ (.A(instruction[30]),
    .B(_04596_),
    .X(_06474_));
 sky130_fd_sc_hd__o211a_4 _06945_ (.A1(instruction[23]),
    .A2(_04607_),
    .B1(_06474_),
    .C1(net272),
    .X(reg2_idx[5]));
 sky130_fd_sc_hd__and3b_4 _06946_ (.A_N(_06455_),
    .B(_04498_),
    .C(_04487_),
    .X(_06475_));
 sky130_fd_sc_hd__or3_4 _06947_ (.A(instruction[6]),
    .B(instruction[5]),
    .C(_06455_),
    .X(_06476_));
 sky130_fd_sc_hd__or2_4 _06948_ (.A(instruction[6]),
    .B(instruction[5]),
    .X(_06477_));
 sky130_fd_sc_hd__nand2_2 _06949_ (.A(_04476_),
    .B(instruction[4]),
    .Y(_06478_));
 sky130_fd_sc_hd__nor2_2 _06950_ (.A(_06477_),
    .B(_06478_),
    .Y(_06479_));
 sky130_fd_sc_hd__or2_4 _06951_ (.A(_06477_),
    .B(_06478_),
    .X(_06480_));
 sky130_fd_sc_hd__a31o_1 _06952_ (.A1(instruction[17]),
    .A2(_06476_),
    .A3(_06480_),
    .B1(net268),
    .X(_06481_));
 sky130_fd_sc_hd__nor2_1 _06953_ (.A(instruction[6]),
    .B(is_load),
    .Y(_06482_));
 sky130_fd_sc_hd__o211a_1 _06954_ (.A1(instruction[40]),
    .A2(_04817_),
    .B1(_06481_),
    .C1(_06482_),
    .X(_06483_));
 sky130_fd_sc_hd__a32o_2 _06955_ (.A1(instruction[24]),
    .A2(net295),
    .A3(is_load),
    .B1(_04860_),
    .B2(_06483_),
    .X(_06484_));
 sky130_fd_sc_hd__nand2_8 _06956_ (.A(net247),
    .B(_06484_),
    .Y(dest_mask[0]));
 sky130_fd_sc_hd__a22o_2 _06957_ (.A1(net295),
    .A2(is_load),
    .B1(net252),
    .B2(_06483_),
    .X(_06485_));
 sky130_fd_sc_hd__nand2_8 _06958_ (.A(net247),
    .B(_06485_),
    .Y(dest_mask[1]));
 sky130_fd_sc_hd__nand2_2 _06959_ (.A(_04487_),
    .B(instruction[5]),
    .Y(_06486_));
 sky130_fd_sc_hd__and4_1 _06960_ (.A(_04487_),
    .B(instruction[5]),
    .C(net294),
    .D(_06439_),
    .X(_06487_));
 sky130_fd_sc_hd__or3_4 _06961_ (.A(net284),
    .B(_06440_),
    .C(_06486_),
    .X(_06488_));
 sky130_fd_sc_hd__nor2_1 _06962_ (.A(net286),
    .B(_05404_),
    .Y(_06489_));
 sky130_fd_sc_hd__nand2_1 _06963_ (.A(net294),
    .B(_05393_),
    .Y(_06490_));
 sky130_fd_sc_hd__and2_1 _06964_ (.A(reg1_val[31]),
    .B(net295),
    .X(_06491_));
 sky130_fd_sc_hd__and3_4 _06965_ (.A(net292),
    .B(reg1_val[31]),
    .C(net295),
    .X(_06492_));
 sky130_fd_sc_hd__xor2_4 _06966_ (.A(net289),
    .B(_06492_),
    .X(_06493_));
 sky130_fd_sc_hd__xnor2_4 _06967_ (.A(net289),
    .B(_06492_),
    .Y(_06494_));
 sky130_fd_sc_hd__and2_2 _06968_ (.A(net294),
    .B(_05382_),
    .X(_06495_));
 sky130_fd_sc_hd__nand2_2 _06969_ (.A(net294),
    .B(_05382_),
    .Y(_06496_));
 sky130_fd_sc_hd__and4_1 _06970_ (.A(net224),
    .B(_06352_),
    .C(_06359_),
    .D(net216),
    .X(_06497_));
 sky130_fd_sc_hd__or4_4 _06971_ (.A(_06347_),
    .B(net221),
    .C(_06360_),
    .D(net214),
    .X(_06498_));
 sky130_fd_sc_hd__or4_4 _06972_ (.A(_06320_),
    .B(_06325_),
    .C(_06333_),
    .D(net228),
    .X(_06499_));
 sky130_fd_sc_hd__nor2_4 _06973_ (.A(_06498_),
    .B(_06499_),
    .Y(_06500_));
 sky130_fd_sc_hd__or2_2 _06974_ (.A(_06498_),
    .B(_06499_),
    .X(_06501_));
 sky130_fd_sc_hd__or2_4 _06975_ (.A(_06283_),
    .B(_06315_),
    .X(_06502_));
 sky130_fd_sc_hd__or2_1 _06976_ (.A(_06185_),
    .B(_06238_),
    .X(_06503_));
 sky130_fd_sc_hd__or4_4 _06977_ (.A(_06121_),
    .B(_06151_),
    .C(_06185_),
    .D(_06238_),
    .X(_06504_));
 sky130_fd_sc_hd__nor4_4 _06978_ (.A(_06031_),
    .B(_06086_),
    .C(_06502_),
    .D(_06504_),
    .Y(_06505_));
 sky130_fd_sc_hd__nand2_1 _06979_ (.A(_06500_),
    .B(_06505_),
    .Y(_06506_));
 sky130_fd_sc_hd__and2_1 _06980_ (.A(_05934_),
    .B(_05974_),
    .X(_06507_));
 sky130_fd_sc_hd__and4_1 _06981_ (.A(_05808_),
    .B(_05872_),
    .C(_05934_),
    .D(_05974_),
    .X(_06508_));
 sky130_fd_sc_hd__and3_4 _06982_ (.A(_06500_),
    .B(_06505_),
    .C(_06508_),
    .X(_06509_));
 sky130_fd_sc_hd__nand3_4 _06983_ (.A(_06500_),
    .B(_06505_),
    .C(_06508_),
    .Y(_06510_));
 sky130_fd_sc_hd__and2_2 _06984_ (.A(_05668_),
    .B(_05725_),
    .X(_06511_));
 sky130_fd_sc_hd__and3_1 _06985_ (.A(_05544_),
    .B(_05609_),
    .C(_06511_),
    .X(_06512_));
 sky130_fd_sc_hd__nand3_2 _06986_ (.A(_05544_),
    .B(_05609_),
    .C(_06511_),
    .Y(_06513_));
 sky130_fd_sc_hd__nand2_1 _06987_ (.A(_06509_),
    .B(_06512_),
    .Y(_06514_));
 sky130_fd_sc_hd__and2_1 _06988_ (.A(_05241_),
    .B(_05306_),
    .X(_06515_));
 sky130_fd_sc_hd__a31o_2 _06989_ (.A1(_06509_),
    .A2(_06512_),
    .A3(_06515_),
    .B1(net183),
    .X(_06516_));
 sky130_fd_sc_hd__xor2_4 _06990_ (.A(_05436_),
    .B(_06516_),
    .X(_06517_));
 sky130_fd_sc_hd__xnor2_1 _06991_ (.A(_05436_),
    .B(_06516_),
    .Y(_06518_));
 sky130_fd_sc_hd__and2_2 _06992_ (.A(net287),
    .B(net289),
    .X(_06519_));
 sky130_fd_sc_hd__nand2_8 _06993_ (.A(net288),
    .B(net289),
    .Y(_06520_));
 sky130_fd_sc_hd__a21o_1 _06994_ (.A1(_06509_),
    .A2(_06512_),
    .B1(net183),
    .X(_06521_));
 sky130_fd_sc_hd__nor2_1 _06995_ (.A(_05306_),
    .B(net183),
    .Y(_06522_));
 sky130_fd_sc_hd__a31o_2 _06996_ (.A1(_05306_),
    .A2(_06509_),
    .A3(_06512_),
    .B1(net183),
    .X(_06523_));
 sky130_fd_sc_hd__xnor2_2 _06997_ (.A(_05241_),
    .B(_06523_),
    .Y(_06524_));
 sky130_fd_sc_hd__xor2_4 _06998_ (.A(_05241_),
    .B(_06523_),
    .X(_06525_));
 sky130_fd_sc_hd__o22a_1 _06999_ (.A1(net288),
    .A2(net68),
    .B1(_06520_),
    .B2(net65),
    .X(_06526_));
 sky130_fd_sc_hd__xnor2_2 _07000_ (.A(net239),
    .B(_06526_),
    .Y(_06527_));
 sky130_fd_sc_hd__or4_2 _07001_ (.A(net292),
    .B(net289),
    .C(reg1_val[2]),
    .D(reg1_val[3]),
    .X(_06528_));
 sky130_fd_sc_hd__nand2_1 _07002_ (.A(net262),
    .B(_06528_),
    .Y(_06529_));
 sky130_fd_sc_hd__o21a_1 _07003_ (.A1(reg1_val[4]),
    .A2(_06528_),
    .B1(net262),
    .X(_06530_));
 sky130_fd_sc_hd__xnor2_2 _07004_ (.A(reg1_val[5]),
    .B(_06530_),
    .Y(_06531_));
 sky130_fd_sc_hd__inv_6 _07005_ (.A(net207),
    .Y(_06532_));
 sky130_fd_sc_hd__o31a_2 _07006_ (.A1(net292),
    .A2(net289),
    .A3(reg1_val[2]),
    .B1(net262),
    .X(_06533_));
 sky130_fd_sc_hd__xnor2_4 _07007_ (.A(reg1_val[3]),
    .B(_06533_),
    .Y(_06534_));
 sky130_fd_sc_hd__xor2_2 _07008_ (.A(reg1_val[4]),
    .B(_06529_),
    .X(_06535_));
 sky130_fd_sc_hd__or2_2 _07009_ (.A(net206),
    .B(_06535_),
    .X(_06536_));
 sky130_fd_sc_hd__nand2_1 _07010_ (.A(net205),
    .B(_06535_),
    .Y(_06537_));
 sky130_fd_sc_hd__nand2_2 _07011_ (.A(_06536_),
    .B(_06537_),
    .Y(_06538_));
 sky130_fd_sc_hd__a21o_2 _07012_ (.A1(_06509_),
    .A2(_06511_),
    .B1(net183),
    .X(_06539_));
 sky130_fd_sc_hd__xor2_4 _07013_ (.A(_05609_),
    .B(_06539_),
    .X(_06540_));
 sky130_fd_sc_hd__xnor2_4 _07014_ (.A(_05609_),
    .B(_06539_),
    .Y(_06541_));
 sky130_fd_sc_hd__mux2_2 _07015_ (.A0(_06536_),
    .A1(_06537_),
    .S(_06532_),
    .X(_06542_));
 sky130_fd_sc_hd__nor2_1 _07016_ (.A(_05668_),
    .B(net183),
    .Y(_06543_));
 sky130_fd_sc_hd__a211o_2 _07017_ (.A1(_05668_),
    .A2(_06509_),
    .B1(_06496_),
    .C1(_05734_),
    .X(_06544_));
 sky130_fd_sc_hd__a211o_2 _07018_ (.A1(net184),
    .A2(_06510_),
    .B1(_06543_),
    .C1(_05725_),
    .X(_06545_));
 sky130_fd_sc_hd__and2_2 _07019_ (.A(_06544_),
    .B(_06545_),
    .X(_06546_));
 sky130_fd_sc_hd__nand2_8 _07020_ (.A(_06544_),
    .B(_06545_),
    .Y(_06547_));
 sky130_fd_sc_hd__o22a_1 _07021_ (.A1(net156),
    .A2(net63),
    .B1(net154),
    .B2(net61),
    .X(_06548_));
 sky130_fd_sc_hd__xnor2_2 _07022_ (.A(net207),
    .B(_06548_),
    .Y(_06549_));
 sky130_fd_sc_hd__or2_1 _07023_ (.A(_06527_),
    .B(_06549_),
    .X(_06550_));
 sky130_fd_sc_hd__o21a_1 _07024_ (.A1(net292),
    .A2(reg1_val[1]),
    .B1(net262),
    .X(_06551_));
 sky130_fd_sc_hd__xnor2_2 _07025_ (.A(reg1_val[2]),
    .B(_06551_),
    .Y(_06552_));
 sky130_fd_sc_hd__and2_1 _07026_ (.A(net239),
    .B(_06552_),
    .X(_06553_));
 sky130_fd_sc_hd__nand2_1 _07027_ (.A(net239),
    .B(_06552_),
    .Y(_06554_));
 sky130_fd_sc_hd__nor2_1 _07028_ (.A(net239),
    .B(_06552_),
    .Y(_06555_));
 sky130_fd_sc_hd__or2_1 _07029_ (.A(_06494_),
    .B(_06552_),
    .X(_06556_));
 sky130_fd_sc_hd__nor2_2 _07030_ (.A(_06553_),
    .B(_06555_),
    .Y(_06557_));
 sky130_fd_sc_hd__nand2_1 _07031_ (.A(_06554_),
    .B(_06556_),
    .Y(_06558_));
 sky130_fd_sc_hd__a22oi_4 _07032_ (.A1(_05306_),
    .A2(_06521_),
    .B1(_06522_),
    .B2(_06514_),
    .Y(_06559_));
 sky130_fd_sc_hd__a22o_2 _07033_ (.A1(_05306_),
    .A2(_06521_),
    .B1(_06522_),
    .B2(_06514_),
    .X(_06560_));
 sky130_fd_sc_hd__a31oi_4 _07034_ (.A1(_05609_),
    .A2(_06509_),
    .A3(_06511_),
    .B1(net183),
    .Y(_06561_));
 sky130_fd_sc_hd__xor2_4 _07035_ (.A(_05544_),
    .B(_06561_),
    .X(_06562_));
 sky130_fd_sc_hd__xnor2_4 _07036_ (.A(_05544_),
    .B(_06561_),
    .Y(_06563_));
 sky130_fd_sc_hd__mux2_1 _07037_ (.A0(_06554_),
    .A1(_06556_),
    .S(net205),
    .X(_06564_));
 sky130_fd_sc_hd__mux2_2 _07038_ (.A0(_06553_),
    .A1(_06555_),
    .S(net205),
    .X(_06565_));
 sky130_fd_sc_hd__o22a_1 _07039_ (.A1(net151),
    .A2(net59),
    .B1(net57),
    .B2(net149),
    .X(_06566_));
 sky130_fd_sc_hd__xnor2_2 _07040_ (.A(net206),
    .B(_06566_),
    .Y(_06567_));
 sky130_fd_sc_hd__xnor2_2 _07041_ (.A(_06527_),
    .B(_06549_),
    .Y(_06568_));
 sky130_fd_sc_hd__o21a_1 _07042_ (.A1(_06567_),
    .A2(_06568_),
    .B1(_06550_),
    .X(_06569_));
 sky130_fd_sc_hd__o22a_1 _07043_ (.A1(net65),
    .A2(net151),
    .B1(net59),
    .B2(net149),
    .X(_06570_));
 sky130_fd_sc_hd__xnor2_1 _07044_ (.A(net206),
    .B(_06570_),
    .Y(_00136_));
 sky130_fd_sc_hd__a41o_1 _07045_ (.A1(_05436_),
    .A2(_06509_),
    .A3(_06512_),
    .A4(_06515_),
    .B1(_05165_),
    .X(_00137_));
 sky130_fd_sc_hd__nand3_2 _07046_ (.A(_05165_),
    .B(_05436_),
    .C(_06515_),
    .Y(_00138_));
 sky130_fd_sc_hd__nor3_4 _07047_ (.A(_06510_),
    .B(_06513_),
    .C(_00138_),
    .Y(_00139_));
 sky130_fd_sc_hd__or3_4 _07048_ (.A(_06510_),
    .B(_06513_),
    .C(_00138_),
    .X(_00140_));
 sky130_fd_sc_hd__nor2_1 _07049_ (.A(_05165_),
    .B(net184),
    .Y(_00141_));
 sky130_fd_sc_hd__a31oi_2 _07050_ (.A1(net184),
    .A2(_00137_),
    .A3(_00140_),
    .B1(_00141_),
    .Y(_00142_));
 sky130_fd_sc_hd__a31o_4 _07051_ (.A1(net184),
    .A2(_00137_),
    .A3(_00140_),
    .B1(_00141_),
    .X(_00143_));
 sky130_fd_sc_hd__o22a_1 _07052_ (.A1(net68),
    .A2(net237),
    .B1(net56),
    .B2(net288),
    .X(_00144_));
 sky130_fd_sc_hd__xnor2_2 _07053_ (.A(_06494_),
    .B(_00144_),
    .Y(_00145_));
 sky130_fd_sc_hd__o22a_1 _07054_ (.A1(net63),
    .A2(net154),
    .B1(net57),
    .B2(net156),
    .X(_00146_));
 sky130_fd_sc_hd__xnor2_1 _07055_ (.A(net207),
    .B(_00146_),
    .Y(_00147_));
 sky130_fd_sc_hd__nor2_1 _07056_ (.A(_00145_),
    .B(_00147_),
    .Y(_00148_));
 sky130_fd_sc_hd__xnor2_1 _07057_ (.A(_00145_),
    .B(_00147_),
    .Y(_00149_));
 sky130_fd_sc_hd__nor2_1 _07058_ (.A(_00136_),
    .B(_00149_),
    .Y(_00150_));
 sky130_fd_sc_hd__xor2_1 _07059_ (.A(_00136_),
    .B(_00149_),
    .X(_00151_));
 sky130_fd_sc_hd__nand2b_1 _07060_ (.A_N(_06569_),
    .B(_00151_),
    .Y(_00152_));
 sky130_fd_sc_hd__or2_1 _07061_ (.A(reg1_val[4]),
    .B(reg1_val[5]),
    .X(_00153_));
 sky130_fd_sc_hd__o31a_1 _07062_ (.A1(reg1_val[6]),
    .A2(_06528_),
    .A3(_00153_),
    .B1(net262),
    .X(_00154_));
 sky130_fd_sc_hd__xnor2_1 _07063_ (.A(reg1_val[7]),
    .B(_00154_),
    .Y(_00155_));
 sky130_fd_sc_hd__o21a_1 _07064_ (.A1(_06528_),
    .A2(_00153_),
    .B1(net262),
    .X(_00156_));
 sky130_fd_sc_hd__xnor2_2 _07065_ (.A(reg1_val[6]),
    .B(_00156_),
    .Y(_00157_));
 sky130_fd_sc_hd__nand2_1 _07066_ (.A(net207),
    .B(_00157_),
    .Y(_00158_));
 sky130_fd_sc_hd__or2_1 _07067_ (.A(net207),
    .B(_00157_),
    .X(_00159_));
 sky130_fd_sc_hd__nand2_2 _07068_ (.A(_00158_),
    .B(_00159_),
    .Y(_00160_));
 sky130_fd_sc_hd__o21ai_4 _07069_ (.A1(net183),
    .A2(_06509_),
    .B1(_05668_),
    .Y(_00161_));
 sky130_fd_sc_hd__nand2_4 _07070_ (.A(_06510_),
    .B(_06543_),
    .Y(_00162_));
 sky130_fd_sc_hd__and2_4 _07071_ (.A(_00161_),
    .B(_00162_),
    .X(_00163_));
 sky130_fd_sc_hd__nand2_4 _07072_ (.A(_00161_),
    .B(_00162_),
    .Y(_00164_));
 sky130_fd_sc_hd__or3b_1 _07073_ (.A(net207),
    .B(_00157_),
    .C_N(net203),
    .X(_00165_));
 sky130_fd_sc_hd__o21a_1 _07074_ (.A1(net202),
    .A2(_00158_),
    .B1(_00165_),
    .X(_00166_));
 sky130_fd_sc_hd__a31oi_4 _07075_ (.A1(_06500_),
    .A2(_06505_),
    .A3(_06507_),
    .B1(net183),
    .Y(_00167_));
 sky130_fd_sc_hd__nor2_1 _07076_ (.A(_05872_),
    .B(net183),
    .Y(_00168_));
 sky130_fd_sc_hd__o21ai_4 _07077_ (.A1(_00167_),
    .A2(_00168_),
    .B1(_05808_),
    .Y(_00169_));
 sky130_fd_sc_hd__or3_4 _07078_ (.A(_05808_),
    .B(_00167_),
    .C(_00168_),
    .X(_00170_));
 sky130_fd_sc_hd__and2_2 _07079_ (.A(_00169_),
    .B(_00170_),
    .X(_00171_));
 sky130_fd_sc_hd__nand2_8 _07080_ (.A(_00169_),
    .B(_00170_),
    .Y(_00172_));
 sky130_fd_sc_hd__o22a_1 _07081_ (.A1(net148),
    .A2(net53),
    .B1(net146),
    .B2(net51),
    .X(_00173_));
 sky130_fd_sc_hd__xnor2_1 _07082_ (.A(net202),
    .B(_00173_),
    .Y(_00174_));
 sky130_fd_sc_hd__or4_2 _07083_ (.A(reg1_val[6]),
    .B(reg1_val[7]),
    .C(_06528_),
    .D(_00153_),
    .X(_00175_));
 sky130_fd_sc_hd__nand2_1 _07084_ (.A(net262),
    .B(_00175_),
    .Y(_00176_));
 sky130_fd_sc_hd__o21a_1 _07085_ (.A1(reg1_val[8]),
    .A2(_00175_),
    .B1(net262),
    .X(_00177_));
 sky130_fd_sc_hd__xnor2_1 _07086_ (.A(reg1_val[9]),
    .B(_00177_),
    .Y(_00178_));
 sky130_fd_sc_hd__xnor2_4 _07087_ (.A(_05872_),
    .B(_00167_),
    .Y(_00179_));
 sky130_fd_sc_hd__xnor2_4 _07088_ (.A(_05881_),
    .B(_00167_),
    .Y(_00180_));
 sky130_fd_sc_hd__xor2_2 _07089_ (.A(reg1_val[8]),
    .B(_00176_),
    .X(_00181_));
 sky130_fd_sc_hd__or2_1 _07090_ (.A(net203),
    .B(_00181_),
    .X(_00182_));
 sky130_fd_sc_hd__nand2_1 _07091_ (.A(net203),
    .B(_00181_),
    .Y(_00183_));
 sky130_fd_sc_hd__nand2_2 _07092_ (.A(_00182_),
    .B(_00183_),
    .Y(_00184_));
 sky130_fd_sc_hd__a21o_1 _07093_ (.A1(_06500_),
    .A2(_06505_),
    .B1(net183),
    .X(_00185_));
 sky130_fd_sc_hd__nor2_1 _07094_ (.A(_05974_),
    .B(net183),
    .Y(_00186_));
 sky130_fd_sc_hd__a31o_4 _07095_ (.A1(_05974_),
    .A2(_06500_),
    .A3(_06505_),
    .B1(net183),
    .X(_00187_));
 sky130_fd_sc_hd__xnor2_4 _07096_ (.A(_05934_),
    .B(_00187_),
    .Y(_00188_));
 sky130_fd_sc_hd__xor2_4 _07097_ (.A(_05934_),
    .B(_00187_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_2 _07098_ (.A0(_00183_),
    .A1(_00182_),
    .S(net181),
    .X(_00190_));
 sky130_fd_sc_hd__o22a_1 _07099_ (.A1(net100),
    .A2(net134),
    .B1(net98),
    .B2(net132),
    .X(_00191_));
 sky130_fd_sc_hd__xnor2_1 _07100_ (.A(net181),
    .B(_00191_),
    .Y(_00192_));
 sky130_fd_sc_hd__nor2_1 _07101_ (.A(_00174_),
    .B(_00192_),
    .Y(_00193_));
 sky130_fd_sc_hd__xnor2_1 _07102_ (.A(_06569_),
    .B(_00151_),
    .Y(_00194_));
 sky130_fd_sc_hd__nand2_1 _07103_ (.A(_00193_),
    .B(_00194_),
    .Y(_00195_));
 sky130_fd_sc_hd__nand2_2 _07104_ (.A(_00152_),
    .B(_00195_),
    .Y(_00196_));
 sky130_fd_sc_hd__or4_2 _07105_ (.A(reg1_val[8]),
    .B(reg1_val[9]),
    .C(reg1_val[10]),
    .D(_00175_),
    .X(_00197_));
 sky130_fd_sc_hd__or4_4 _07106_ (.A(reg1_val[11]),
    .B(reg1_val[12]),
    .C(reg1_val[13]),
    .D(_00197_),
    .X(_00198_));
 sky130_fd_sc_hd__or3_1 _07107_ (.A(net291),
    .B(net290),
    .C(_00198_),
    .X(_00199_));
 sky130_fd_sc_hd__or2_2 _07108_ (.A(reg1_val[16]),
    .B(reg1_val[17]),
    .X(_00200_));
 sky130_fd_sc_hd__or3_4 _07109_ (.A(reg1_val[18]),
    .B(reg1_val[19]),
    .C(_00200_),
    .X(_00201_));
 sky130_fd_sc_hd__o41a_4 _07110_ (.A1(net291),
    .A2(net290),
    .A3(_00198_),
    .A4(_00201_),
    .B1(net262),
    .X(_00202_));
 sky130_fd_sc_hd__or2_1 _07111_ (.A(reg1_val[20]),
    .B(reg1_val[21]),
    .X(_00203_));
 sky130_fd_sc_hd__or2_1 _07112_ (.A(reg1_val[22]),
    .B(_00203_),
    .X(_00204_));
 sky130_fd_sc_hd__and2_1 _07113_ (.A(net262),
    .B(_00204_),
    .X(_00205_));
 sky130_fd_sc_hd__o21ai_1 _07114_ (.A1(_00202_),
    .A2(_00205_),
    .B1(reg1_val[23]),
    .Y(_00206_));
 sky130_fd_sc_hd__or3_1 _07115_ (.A(reg1_val[23]),
    .B(_00202_),
    .C(_00205_),
    .X(_00207_));
 sky130_fd_sc_hd__and2_2 _07116_ (.A(_00206_),
    .B(_00207_),
    .X(_00208_));
 sky130_fd_sc_hd__and3_1 _07117_ (.A(net294),
    .B(_05382_),
    .C(net228),
    .X(_00209_));
 sky130_fd_sc_hd__a211o_1 _07118_ (.A1(net225),
    .A2(_06497_),
    .B1(_06496_),
    .C1(_06333_),
    .X(_00210_));
 sky130_fd_sc_hd__a211o_1 _07119_ (.A1(net184),
    .A2(_06498_),
    .B1(_00209_),
    .C1(_06332_),
    .X(_00211_));
 sky130_fd_sc_hd__and2_1 _07120_ (.A(_00210_),
    .B(_00211_),
    .X(_00212_));
 sky130_fd_sc_hd__nand2_4 _07121_ (.A(_00210_),
    .B(_00211_),
    .Y(_00213_));
 sky130_fd_sc_hd__o311a_2 _07122_ (.A1(reg1_val[20]),
    .A2(_00199_),
    .A3(_00201_),
    .B1(reg1_val[21]),
    .C1(net261),
    .X(_00214_));
 sky130_fd_sc_hd__a211oi_4 _07123_ (.A1(reg1_val[20]),
    .A2(net261),
    .B1(_00202_),
    .C1(reg1_val[21]),
    .Y(_00215_));
 sky130_fd_sc_hd__nor2_4 _07124_ (.A(_00214_),
    .B(_00215_),
    .Y(_00216_));
 sky130_fd_sc_hd__clkinv_4 _07125_ (.A(_00216_),
    .Y(_00217_));
 sky130_fd_sc_hd__o311a_1 _07126_ (.A1(_00199_),
    .A2(_00201_),
    .A3(_00203_),
    .B1(net261),
    .C1(reg1_val[22]),
    .X(_00218_));
 sky130_fd_sc_hd__a211oi_2 _07127_ (.A1(net261),
    .A2(_00203_),
    .B1(_00202_),
    .C1(reg1_val[22]),
    .Y(_00219_));
 sky130_fd_sc_hd__nor2_1 _07128_ (.A(_00218_),
    .B(_00219_),
    .Y(_00220_));
 sky130_fd_sc_hd__or4_2 _07129_ (.A(_00214_),
    .B(_00215_),
    .C(_00218_),
    .D(_00219_),
    .X(_00221_));
 sky130_fd_sc_hd__o22ai_2 _07130_ (.A1(_00214_),
    .A2(_00215_),
    .B1(_00218_),
    .B2(_00219_),
    .Y(_00222_));
 sky130_fd_sc_hd__nand2_2 _07131_ (.A(_00221_),
    .B(_00222_),
    .Y(_00223_));
 sky130_fd_sc_hd__a21oi_4 _07132_ (.A1(net184),
    .A2(_06498_),
    .B1(net228),
    .Y(_00224_));
 sky130_fd_sc_hd__and2_2 _07133_ (.A(_06498_),
    .B(_00209_),
    .X(_00225_));
 sky130_fd_sc_hd__nor2_4 _07134_ (.A(_00224_),
    .B(_00225_),
    .Y(_00226_));
 sky130_fd_sc_hd__or2_1 _07135_ (.A(_00224_),
    .B(_00225_),
    .X(_00227_));
 sky130_fd_sc_hd__nor2_1 _07136_ (.A(net95),
    .B(_00221_),
    .Y(_00228_));
 sky130_fd_sc_hd__mux2_1 _07137_ (.A0(_00221_),
    .A1(_00222_),
    .S(net95),
    .X(_00229_));
 sky130_fd_sc_hd__o22a_1 _07138_ (.A1(net129),
    .A2(net48),
    .B1(net128),
    .B2(net46),
    .X(_00230_));
 sky130_fd_sc_hd__xnor2_1 _07139_ (.A(net97),
    .B(_00230_),
    .Y(_00231_));
 sky130_fd_sc_hd__or3_2 _07140_ (.A(reg1_val[23]),
    .B(_00201_),
    .C(_00204_),
    .X(_00232_));
 sky130_fd_sc_hd__or4_4 _07141_ (.A(net291),
    .B(net290),
    .C(_00198_),
    .D(_00232_),
    .X(_00233_));
 sky130_fd_sc_hd__or2_2 _07142_ (.A(reg1_val[24]),
    .B(reg1_val[25]),
    .X(_00234_));
 sky130_fd_sc_hd__or2_1 _07143_ (.A(_00232_),
    .B(_00234_),
    .X(_00235_));
 sky130_fd_sc_hd__o41a_1 _07144_ (.A1(net291),
    .A2(net290),
    .A3(_00198_),
    .A4(_00235_),
    .B1(net261),
    .X(_00236_));
 sky130_fd_sc_hd__a21oi_1 _07145_ (.A1(reg1_val[26]),
    .A2(net261),
    .B1(_00236_),
    .Y(_00237_));
 sky130_fd_sc_hd__xnor2_2 _07146_ (.A(reg1_val[27]),
    .B(_00237_),
    .Y(_00238_));
 sky130_fd_sc_hd__and3_2 _07147_ (.A(net295),
    .B(_05382_),
    .C(net214),
    .X(_00239_));
 sky130_fd_sc_hd__xnor2_4 _07148_ (.A(_06359_),
    .B(_00239_),
    .Y(_00240_));
 sky130_fd_sc_hd__xnor2_1 _07149_ (.A(_06360_),
    .B(_00239_),
    .Y(_00241_));
 sky130_fd_sc_hd__o41a_1 _07150_ (.A1(net291),
    .A2(net290),
    .A3(_00198_),
    .A4(_00232_),
    .B1(net261),
    .X(_00242_));
 sky130_fd_sc_hd__o211ai_2 _07151_ (.A1(reg1_val[24]),
    .A2(_00233_),
    .B1(net261),
    .C1(reg1_val[25]),
    .Y(_00243_));
 sky130_fd_sc_hd__a211o_1 _07152_ (.A1(reg1_val[24]),
    .A2(net261),
    .B1(_00242_),
    .C1(reg1_val[25]),
    .X(_00244_));
 sky130_fd_sc_hd__and2_4 _07153_ (.A(_00243_),
    .B(_00244_),
    .X(_00245_));
 sky130_fd_sc_hd__xor2_2 _07154_ (.A(reg1_val[26]),
    .B(_00236_),
    .X(_00246_));
 sky130_fd_sc_hd__and3_1 _07155_ (.A(_00243_),
    .B(_00244_),
    .C(_00246_),
    .X(_00247_));
 sky130_fd_sc_hd__a21oi_2 _07156_ (.A1(_00243_),
    .A2(_00244_),
    .B1(_00246_),
    .Y(_00248_));
 sky130_fd_sc_hd__nor2_2 _07157_ (.A(_00247_),
    .B(_00248_),
    .Y(_00249_));
 sky130_fd_sc_hd__and2b_1 _07158_ (.A_N(net92),
    .B(_00247_),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _07159_ (.A0(_00247_),
    .A1(_00248_),
    .S(net92),
    .X(_00251_));
 sky130_fd_sc_hd__a22o_1 _07160_ (.A1(_00240_),
    .A2(net44),
    .B1(net42),
    .B2(net214),
    .X(_00252_));
 sky130_fd_sc_hd__xor2_1 _07161_ (.A(net94),
    .B(_00252_),
    .X(_00253_));
 sky130_fd_sc_hd__xor2_1 _07162_ (.A(_00231_),
    .B(_00253_),
    .X(_00254_));
 sky130_fd_sc_hd__o211a_4 _07163_ (.A1(_06360_),
    .A2(net214),
    .B1(net294),
    .C1(_05382_),
    .X(_00255_));
 sky130_fd_sc_hd__o311a_2 _07164_ (.A1(net221),
    .A2(_06360_),
    .A3(net214),
    .B1(_05382_),
    .C1(net294),
    .X(_00256_));
 sky130_fd_sc_hd__xnor2_2 _07165_ (.A(_06347_),
    .B(_00256_),
    .Y(_00257_));
 sky130_fd_sc_hd__xnor2_4 _07166_ (.A(_06346_),
    .B(_00256_),
    .Y(_00258_));
 sky130_fd_sc_hd__xor2_2 _07167_ (.A(reg1_val[24]),
    .B(_00242_),
    .X(_00259_));
 sky130_fd_sc_hd__and3_1 _07168_ (.A(_00206_),
    .B(_00207_),
    .C(_00259_),
    .X(_00260_));
 sky130_fd_sc_hd__a21oi_1 _07169_ (.A1(_00206_),
    .A2(_00207_),
    .B1(_00259_),
    .Y(_00261_));
 sky130_fd_sc_hd__nor2_1 _07170_ (.A(_00260_),
    .B(_00261_),
    .Y(_00262_));
 sky130_fd_sc_hd__inv_2 _07171_ (.A(net40),
    .Y(_00263_));
 sky130_fd_sc_hd__xnor2_4 _07172_ (.A(net221),
    .B(_00255_),
    .Y(_00264_));
 sky130_fd_sc_hd__xnor2_4 _07173_ (.A(_06352_),
    .B(_00255_),
    .Y(_00265_));
 sky130_fd_sc_hd__mux2_2 _07174_ (.A0(_00260_),
    .A1(_00261_),
    .S(net90),
    .X(_00266_));
 sky130_fd_sc_hd__inv_2 _07175_ (.A(net37),
    .Y(_00267_));
 sky130_fd_sc_hd__a22o_1 _07176_ (.A1(_00258_),
    .A2(net39),
    .B1(_00265_),
    .B2(net37),
    .X(_00268_));
 sky130_fd_sc_hd__xor2_1 _07177_ (.A(net91),
    .B(_00268_),
    .X(_00269_));
 sky130_fd_sc_hd__nand2_1 _07178_ (.A(_00254_),
    .B(_00269_),
    .Y(_00270_));
 sky130_fd_sc_hd__a21bo_2 _07179_ (.A1(_00231_),
    .A2(_00253_),
    .B1_N(_00270_),
    .X(_00271_));
 sky130_fd_sc_hd__inv_2 _07180_ (.A(_00271_),
    .Y(_00272_));
 sky130_fd_sc_hd__o31a_1 _07181_ (.A1(net291),
    .A2(net290),
    .A3(_00198_),
    .B1(net261),
    .X(_00273_));
 sky130_fd_sc_hd__o41a_4 _07182_ (.A1(net291),
    .A2(net290),
    .A3(reg1_val[16]),
    .A4(_00198_),
    .B1(net261),
    .X(_00274_));
 sky130_fd_sc_hd__xor2_2 _07183_ (.A(reg1_val[17]),
    .B(_00274_),
    .X(_00275_));
 sky130_fd_sc_hd__xnor2_4 _07184_ (.A(reg1_val[17]),
    .B(_00274_),
    .Y(_00276_));
 sky130_fd_sc_hd__o41a_1 _07185_ (.A1(reg1_val[11]),
    .A2(reg1_val[12]),
    .A3(reg1_val[13]),
    .A4(_00197_),
    .B1(net261),
    .X(_00277_));
 sky130_fd_sc_hd__o21a_1 _07186_ (.A1(net291),
    .A2(_00198_),
    .B1(net261),
    .X(_00278_));
 sky130_fd_sc_hd__xnor2_1 _07187_ (.A(net290),
    .B(_00278_),
    .Y(_00279_));
 sky130_fd_sc_hd__xnor2_2 _07188_ (.A(reg1_val[16]),
    .B(_00273_),
    .Y(_00280_));
 sky130_fd_sc_hd__nor2_1 _07189_ (.A(net121),
    .B(_00280_),
    .Y(_00281_));
 sky130_fd_sc_hd__nand2_2 _07190_ (.A(net121),
    .B(_00280_),
    .Y(_00282_));
 sky130_fd_sc_hd__and2b_2 _07191_ (.A_N(_00281_),
    .B(_00282_),
    .X(_00283_));
 sky130_fd_sc_hd__nand2b_2 _07192_ (.A_N(_00281_),
    .B(_00282_),
    .Y(_00284_));
 sky130_fd_sc_hd__o41a_4 _07193_ (.A1(_06498_),
    .A2(_06499_),
    .A3(_06502_),
    .A4(_06503_),
    .B1(net184),
    .X(_00285_));
 sky130_fd_sc_hd__xnor2_4 _07194_ (.A(_06151_),
    .B(_00285_),
    .Y(_00286_));
 sky130_fd_sc_hd__xor2_4 _07195_ (.A(_06151_),
    .B(_00285_),
    .X(_00287_));
 sky130_fd_sc_hd__o31a_4 _07196_ (.A1(_06498_),
    .A2(_06499_),
    .A3(_06502_),
    .B1(net184),
    .X(_00288_));
 sky130_fd_sc_hd__o41a_4 _07197_ (.A1(_06238_),
    .A2(_06498_),
    .A3(_06499_),
    .A4(_06502_),
    .B1(net184),
    .X(_00289_));
 sky130_fd_sc_hd__xnor2_4 _07198_ (.A(_06185_),
    .B(_00289_),
    .Y(_00290_));
 sky130_fd_sc_hd__xor2_2 _07199_ (.A(_06185_),
    .B(_00289_),
    .X(_00291_));
 sky130_fd_sc_hd__or3_2 _07200_ (.A(net125),
    .B(net121),
    .C(_00280_),
    .X(_00292_));
 sky130_fd_sc_hd__o21a_2 _07201_ (.A1(net124),
    .A2(_00282_),
    .B1(_00292_),
    .X(_00293_));
 sky130_fd_sc_hd__o21ai_2 _07202_ (.A1(net124),
    .A2(_00282_),
    .B1(_00292_),
    .Y(_00294_));
 sky130_fd_sc_hd__a22o_1 _07203_ (.A1(_00283_),
    .A2(_00287_),
    .B1(net116),
    .B2(_00294_),
    .X(_00295_));
 sky130_fd_sc_hd__xnor2_1 _07204_ (.A(net124),
    .B(_00295_),
    .Y(_00296_));
 sky130_fd_sc_hd__o41a_2 _07205_ (.A1(reg1_val[14]),
    .A2(reg1_val[15]),
    .A3(_00198_),
    .A4(_00200_),
    .B1(net262),
    .X(_00297_));
 sky130_fd_sc_hd__and3_1 _07206_ (.A(reg1_val[18]),
    .B(reg1_val[31]),
    .C(net295),
    .X(_00298_));
 sky130_fd_sc_hd__o21ai_2 _07207_ (.A1(_00297_),
    .A2(_00298_),
    .B1(reg1_val[19]),
    .Y(_00299_));
 sky130_fd_sc_hd__or3_2 _07208_ (.A(reg1_val[19]),
    .B(_00297_),
    .C(_00298_),
    .X(_00300_));
 sky130_fd_sc_hd__and2_4 _07209_ (.A(_00299_),
    .B(_00300_),
    .X(_00301_));
 sky130_fd_sc_hd__xor2_2 _07210_ (.A(reg1_val[20]),
    .B(_00202_),
    .X(_00302_));
 sky130_fd_sc_hd__a21oi_2 _07211_ (.A1(_00299_),
    .A2(_00300_),
    .B1(_00302_),
    .Y(_00303_));
 sky130_fd_sc_hd__and3_1 _07212_ (.A(_00299_),
    .B(_00300_),
    .C(_00302_),
    .X(_00304_));
 sky130_fd_sc_hd__nor2_2 _07213_ (.A(_00303_),
    .B(_00304_),
    .Y(_00305_));
 sky130_fd_sc_hd__o21a_1 _07214_ (.A1(_06498_),
    .A2(_06499_),
    .B1(net184),
    .X(_00306_));
 sky130_fd_sc_hd__nand2_2 _07215_ (.A(_06315_),
    .B(net184),
    .Y(_00307_));
 sky130_fd_sc_hd__o22a_4 _07216_ (.A1(_06315_),
    .A2(_00306_),
    .B1(_00307_),
    .B2(_06500_),
    .X(_00308_));
 sky130_fd_sc_hd__o22ai_4 _07217_ (.A1(_06315_),
    .A2(_00306_),
    .B1(_00307_),
    .B2(_06500_),
    .Y(_00309_));
 sky130_fd_sc_hd__mux2_2 _07218_ (.A0(_00304_),
    .A1(_00303_),
    .S(_00216_),
    .X(_00310_));
 sky130_fd_sc_hd__a31o_4 _07219_ (.A1(_06332_),
    .A2(_06341_),
    .A3(_06497_),
    .B1(_06496_),
    .X(_00311_));
 sky130_fd_sc_hd__o41ai_4 _07220_ (.A1(_06325_),
    .A2(_06333_),
    .A3(net228),
    .A4(_06498_),
    .B1(net184),
    .Y(_00312_));
 sky130_fd_sc_hd__xor2_4 _07221_ (.A(_06320_),
    .B(_00312_),
    .X(_00313_));
 sky130_fd_sc_hd__xnor2_4 _07222_ (.A(_06320_),
    .B(net139),
    .Y(_00314_));
 sky130_fd_sc_hd__a22o_1 _07223_ (.A1(net31),
    .A2(_00308_),
    .B1(net29),
    .B2(net113),
    .X(_00315_));
 sky130_fd_sc_hd__xnor2_1 _07224_ (.A(net49),
    .B(_00315_),
    .Y(_00316_));
 sky130_fd_sc_hd__and2_1 _07225_ (.A(_00296_),
    .B(_00316_),
    .X(_00317_));
 sky130_fd_sc_hd__nor2_1 _07226_ (.A(_00296_),
    .B(_00316_),
    .Y(_00318_));
 sky130_fd_sc_hd__nor2_2 _07227_ (.A(_00317_),
    .B(_00318_),
    .Y(_00319_));
 sky130_fd_sc_hd__xnor2_2 _07228_ (.A(reg1_val[18]),
    .B(_00297_),
    .Y(_00320_));
 sky130_fd_sc_hd__nor2_1 _07229_ (.A(net124),
    .B(_00320_),
    .Y(_00321_));
 sky130_fd_sc_hd__and2_1 _07230_ (.A(net124),
    .B(_00320_),
    .X(_00322_));
 sky130_fd_sc_hd__or2_2 _07231_ (.A(_00321_),
    .B(_00322_),
    .X(_00323_));
 sky130_fd_sc_hd__xor2_4 _07232_ (.A(_06238_),
    .B(_00288_),
    .X(_00324_));
 sky130_fd_sc_hd__xnor2_4 _07233_ (.A(_06238_),
    .B(_00288_),
    .Y(_00325_));
 sky130_fd_sc_hd__a211oi_2 _07234_ (.A1(_00299_),
    .A2(_00300_),
    .B1(_00320_),
    .C1(net124),
    .Y(_00326_));
 sky130_fd_sc_hd__a21oi_4 _07235_ (.A1(net89),
    .A2(_00322_),
    .B1(_00326_),
    .Y(_00327_));
 sky130_fd_sc_hd__o31a_4 _07236_ (.A1(_06315_),
    .A2(_06498_),
    .A3(_06499_),
    .B1(net184),
    .X(_00328_));
 sky130_fd_sc_hd__xnor2_4 _07237_ (.A(_06283_),
    .B(_00328_),
    .Y(_00329_));
 sky130_fd_sc_hd__xnor2_4 _07238_ (.A(_06291_),
    .B(_00328_),
    .Y(_00330_));
 sky130_fd_sc_hd__o22a_2 _07239_ (.A1(net27),
    .A2(net111),
    .B1(net25),
    .B2(net109),
    .X(_00331_));
 sky130_fd_sc_hd__xnor2_4 _07240_ (.A(net88),
    .B(_00331_),
    .Y(_00332_));
 sky130_fd_sc_hd__xnor2_4 _07241_ (.A(_00319_),
    .B(_00332_),
    .Y(_00333_));
 sky130_fd_sc_hd__xor2_4 _07242_ (.A(_00271_),
    .B(_00333_),
    .X(_00334_));
 sky130_fd_sc_hd__a21o_1 _07243_ (.A1(_00152_),
    .A2(_00195_),
    .B1(_00334_),
    .X(_00335_));
 sky130_fd_sc_hd__xnor2_4 _07244_ (.A(_00196_),
    .B(_00334_),
    .Y(_00336_));
 sky130_fd_sc_hd__o31a_2 _07245_ (.A1(reg1_val[11]),
    .A2(reg1_val[12]),
    .A3(_00197_),
    .B1(net262),
    .X(_00337_));
 sky130_fd_sc_hd__xnor2_4 _07246_ (.A(reg1_val[13]),
    .B(_00337_),
    .Y(_00338_));
 sky130_fd_sc_hd__inv_6 _07247_ (.A(net138),
    .Y(_00339_));
 sky130_fd_sc_hd__nand2_2 _07248_ (.A(net262),
    .B(_00197_),
    .Y(_00340_));
 sky130_fd_sc_hd__xor2_4 _07249_ (.A(reg1_val[11]),
    .B(_00340_),
    .X(_00341_));
 sky130_fd_sc_hd__inv_6 _07250_ (.A(net135),
    .Y(_00342_));
 sky130_fd_sc_hd__o21a_1 _07251_ (.A1(reg1_val[11]),
    .A2(_00197_),
    .B1(net261),
    .X(_00343_));
 sky130_fd_sc_hd__xnor2_2 _07252_ (.A(reg1_val[12]),
    .B(_00343_),
    .Y(_00344_));
 sky130_fd_sc_hd__nand2_1 _07253_ (.A(net135),
    .B(_00344_),
    .Y(_00345_));
 sky130_fd_sc_hd__or2_1 _07254_ (.A(net135),
    .B(_00344_),
    .X(_00346_));
 sky130_fd_sc_hd__nand2_1 _07255_ (.A(_00345_),
    .B(_00346_),
    .Y(_00347_));
 sky130_fd_sc_hd__a22oi_4 _07256_ (.A1(_05974_),
    .A2(_00185_),
    .B1(_00186_),
    .B2(_06506_),
    .Y(_00348_));
 sky130_fd_sc_hd__a22o_1 _07257_ (.A1(_05974_),
    .A2(_00185_),
    .B1(_00186_),
    .B2(_06506_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _07258_ (.A0(_00345_),
    .A1(_00346_),
    .S(net137),
    .X(_00350_));
 sky130_fd_sc_hd__o31ai_4 _07259_ (.A1(_06501_),
    .A2(_06502_),
    .A3(_06504_),
    .B1(net184),
    .Y(_00351_));
 sky130_fd_sc_hd__o41a_4 _07260_ (.A1(_06086_),
    .A2(_06501_),
    .A3(_06502_),
    .A4(_06504_),
    .B1(net184),
    .X(_00352_));
 sky130_fd_sc_hd__xnor2_2 _07261_ (.A(_06031_),
    .B(_00352_),
    .Y(_00353_));
 sky130_fd_sc_hd__xor2_4 _07262_ (.A(_06031_),
    .B(_00352_),
    .X(_00354_));
 sky130_fd_sc_hd__o22a_1 _07263_ (.A1(net86),
    .A2(net84),
    .B1(net82),
    .B2(net80),
    .X(_00355_));
 sky130_fd_sc_hd__xnor2_1 _07264_ (.A(net137),
    .B(_00355_),
    .Y(_00356_));
 sky130_fd_sc_hd__xnor2_2 _07265_ (.A(reg1_val[14]),
    .B(_00277_),
    .Y(_00357_));
 sky130_fd_sc_hd__or2_2 _07266_ (.A(net137),
    .B(_00357_),
    .X(_00358_));
 sky130_fd_sc_hd__nand2_1 _07267_ (.A(_00338_),
    .B(_00357_),
    .Y(_00359_));
 sky130_fd_sc_hd__nand2_4 _07268_ (.A(_00358_),
    .B(_00359_),
    .Y(_00360_));
 sky130_fd_sc_hd__xnor2_4 _07269_ (.A(_06086_),
    .B(_00351_),
    .Y(_00361_));
 sky130_fd_sc_hd__xor2_4 _07270_ (.A(_06086_),
    .B(_00351_),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _07271_ (.A0(_00359_),
    .A1(_00358_),
    .S(net122),
    .X(_00363_));
 sky130_fd_sc_hd__a21oi_4 _07272_ (.A1(_06151_),
    .A2(net184),
    .B1(_00285_),
    .Y(_00364_));
 sky130_fd_sc_hd__xor2_2 _07273_ (.A(_06121_),
    .B(_00364_),
    .X(_00365_));
 sky130_fd_sc_hd__xnor2_4 _07274_ (.A(_06121_),
    .B(_00364_),
    .Y(_00366_));
 sky130_fd_sc_hd__o22a_1 _07275_ (.A1(net78),
    .A2(net76),
    .B1(net74),
    .B2(net72),
    .X(_00367_));
 sky130_fd_sc_hd__xnor2_1 _07276_ (.A(net121),
    .B(_00367_),
    .Y(_00368_));
 sky130_fd_sc_hd__nor2_1 _07277_ (.A(_00356_),
    .B(_00368_),
    .Y(_00369_));
 sky130_fd_sc_hd__and2_1 _07278_ (.A(_00356_),
    .B(_00368_),
    .X(_00370_));
 sky130_fd_sc_hd__nor2_1 _07279_ (.A(_00369_),
    .B(_00370_),
    .Y(_00371_));
 sky130_fd_sc_hd__a22o_1 _07280_ (.A1(_00283_),
    .A2(net116),
    .B1(_00294_),
    .B2(_00324_),
    .X(_00372_));
 sky130_fd_sc_hd__xnor2_1 _07281_ (.A(net124),
    .B(_00372_),
    .Y(_00373_));
 sky130_fd_sc_hd__xnor2_4 _07282_ (.A(_06325_),
    .B(_00311_),
    .Y(_00374_));
 sky130_fd_sc_hd__xor2_4 _07283_ (.A(_06325_),
    .B(_00311_),
    .X(_00375_));
 sky130_fd_sc_hd__a22o_1 _07284_ (.A1(net31),
    .A2(net113),
    .B1(_00374_),
    .B2(net29),
    .X(_00376_));
 sky130_fd_sc_hd__xnor2_1 _07285_ (.A(net49),
    .B(_00376_),
    .Y(_00377_));
 sky130_fd_sc_hd__and2_1 _07286_ (.A(_00373_),
    .B(_00377_),
    .X(_00378_));
 sky130_fd_sc_hd__xor2_1 _07287_ (.A(_00373_),
    .B(_00377_),
    .X(_00379_));
 sky130_fd_sc_hd__o22a_1 _07288_ (.A1(_00309_),
    .A2(net25),
    .B1(net110),
    .B2(net27),
    .X(_00380_));
 sky130_fd_sc_hd__xnor2_1 _07289_ (.A(net88),
    .B(_00380_),
    .Y(_00381_));
 sky130_fd_sc_hd__and2_1 _07290_ (.A(_00379_),
    .B(_00381_),
    .X(_00382_));
 sky130_fd_sc_hd__o21a_1 _07291_ (.A1(_00378_),
    .A2(_00382_),
    .B1(_00371_),
    .X(_00383_));
 sky130_fd_sc_hd__nor3_1 _07292_ (.A(_00371_),
    .B(_00378_),
    .C(_00382_),
    .Y(_00384_));
 sky130_fd_sc_hd__nor2_1 _07293_ (.A(_00383_),
    .B(_00384_),
    .Y(_00385_));
 sky130_fd_sc_hd__o31a_1 _07294_ (.A1(reg1_val[8]),
    .A2(reg1_val[9]),
    .A3(_00175_),
    .B1(net262),
    .X(_00386_));
 sky130_fd_sc_hd__xnor2_2 _07295_ (.A(reg1_val[10]),
    .B(_00386_),
    .Y(_00387_));
 sky130_fd_sc_hd__nand2_1 _07296_ (.A(net182),
    .B(_00387_),
    .Y(_00388_));
 sky130_fd_sc_hd__or2_1 _07297_ (.A(net182),
    .B(_00387_),
    .X(_00389_));
 sky130_fd_sc_hd__nand2_1 _07298_ (.A(_00388_),
    .B(_00389_),
    .Y(_00390_));
 sky130_fd_sc_hd__mux2_1 _07299_ (.A0(_00388_),
    .A1(_00389_),
    .S(_00341_),
    .X(_00391_));
 sky130_fd_sc_hd__o22a_1 _07300_ (.A1(net98),
    .A2(net106),
    .B1(net104),
    .B2(net84),
    .X(_00392_));
 sky130_fd_sc_hd__xnor2_1 _07301_ (.A(net135),
    .B(_00392_),
    .Y(_00393_));
 sky130_fd_sc_hd__o22a_1 _07302_ (.A1(net120),
    .A2(net74),
    .B1(net72),
    .B2(net78),
    .X(_00394_));
 sky130_fd_sc_hd__xnor2_1 _07303_ (.A(net121),
    .B(_00394_),
    .Y(_00395_));
 sky130_fd_sc_hd__o22a_1 _07304_ (.A1(net86),
    .A2(net80),
    .B1(net76),
    .B2(net82),
    .X(_00396_));
 sky130_fd_sc_hd__xnor2_1 _07305_ (.A(net137),
    .B(_00396_),
    .Y(_00397_));
 sky130_fd_sc_hd__xnor2_1 _07306_ (.A(_00393_),
    .B(_00395_),
    .Y(_00398_));
 sky130_fd_sc_hd__nor2_2 _07307_ (.A(_00397_),
    .B(_00398_),
    .Y(_00399_));
 sky130_fd_sc_hd__o21bai_1 _07308_ (.A1(_00393_),
    .A2(_00395_),
    .B1_N(_00399_),
    .Y(_00400_));
 sky130_fd_sc_hd__and2_1 _07309_ (.A(_00385_),
    .B(_00400_),
    .X(_00401_));
 sky130_fd_sc_hd__xnor2_1 _07310_ (.A(_00385_),
    .B(_00400_),
    .Y(_00402_));
 sky130_fd_sc_hd__o22a_1 _07311_ (.A1(net68),
    .A2(net151),
    .B1(net149),
    .B2(net65),
    .X(_00403_));
 sky130_fd_sc_hd__xnor2_2 _07312_ (.A(net206),
    .B(_00403_),
    .Y(_00404_));
 sky130_fd_sc_hd__a21oi_4 _07313_ (.A1(_06495_),
    .A2(_00140_),
    .B1(_05024_),
    .Y(_00405_));
 sky130_fd_sc_hd__nand2_4 _07314_ (.A(_05024_),
    .B(_06495_),
    .Y(_00406_));
 sky130_fd_sc_hd__nor2_8 _07315_ (.A(_00139_),
    .B(_00406_),
    .Y(_00407_));
 sky130_fd_sc_hd__nor2_4 _07316_ (.A(_00405_),
    .B(_00407_),
    .Y(_00408_));
 sky130_fd_sc_hd__or2_2 _07317_ (.A(_00405_),
    .B(_00407_),
    .X(_00409_));
 sky130_fd_sc_hd__o22a_1 _07318_ (.A1(_06520_),
    .A2(net56),
    .B1(net17),
    .B2(net288),
    .X(_00410_));
 sky130_fd_sc_hd__xnor2_2 _07319_ (.A(net239),
    .B(_00410_),
    .Y(_00411_));
 sky130_fd_sc_hd__o22a_1 _07320_ (.A1(net156),
    .A2(net59),
    .B1(net57),
    .B2(net154),
    .X(_00412_));
 sky130_fd_sc_hd__xnor2_2 _07321_ (.A(net207),
    .B(_00412_),
    .Y(_00413_));
 sky130_fd_sc_hd__nor2_1 _07322_ (.A(_00411_),
    .B(_00413_),
    .Y(_00414_));
 sky130_fd_sc_hd__xnor2_2 _07323_ (.A(_00411_),
    .B(_00413_),
    .Y(_00415_));
 sky130_fd_sc_hd__nor2_1 _07324_ (.A(_00404_),
    .B(_00415_),
    .Y(_00416_));
 sky130_fd_sc_hd__xnor2_2 _07325_ (.A(_00404_),
    .B(_00415_),
    .Y(_00417_));
 sky130_fd_sc_hd__o22a_1 _07326_ (.A1(net61),
    .A2(net148),
    .B1(net53),
    .B2(net146),
    .X(_00418_));
 sky130_fd_sc_hd__xnor2_1 _07327_ (.A(net202),
    .B(_00418_),
    .Y(_00419_));
 sky130_fd_sc_hd__o22a_1 _07328_ (.A1(net51),
    .A2(net134),
    .B1(net132),
    .B2(net100),
    .X(_00420_));
 sky130_fd_sc_hd__xnor2_1 _07329_ (.A(net181),
    .B(_00420_),
    .Y(_00421_));
 sky130_fd_sc_hd__nor2_1 _07330_ (.A(_00419_),
    .B(_00421_),
    .Y(_00422_));
 sky130_fd_sc_hd__o22a_1 _07331_ (.A1(net100),
    .A2(net106),
    .B1(net104),
    .B2(net98),
    .X(_00423_));
 sky130_fd_sc_hd__xnor2_2 _07332_ (.A(net135),
    .B(_00423_),
    .Y(_00424_));
 sky130_fd_sc_hd__o22a_1 _07333_ (.A1(net63),
    .A2(net148),
    .B1(net146),
    .B2(net61),
    .X(_00425_));
 sky130_fd_sc_hd__xnor2_2 _07334_ (.A(net202),
    .B(_00425_),
    .Y(_00426_));
 sky130_fd_sc_hd__nor2_1 _07335_ (.A(_00424_),
    .B(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__xor2_2 _07336_ (.A(_00424_),
    .B(_00426_),
    .X(_00428_));
 sky130_fd_sc_hd__o22a_1 _07337_ (.A1(net53),
    .A2(net134),
    .B1(net132),
    .B2(net51),
    .X(_00429_));
 sky130_fd_sc_hd__xnor2_2 _07338_ (.A(net181),
    .B(_00429_),
    .Y(_00430_));
 sky130_fd_sc_hd__inv_2 _07339_ (.A(_00430_),
    .Y(_00431_));
 sky130_fd_sc_hd__xnor2_2 _07340_ (.A(_00428_),
    .B(_00430_),
    .Y(_00432_));
 sky130_fd_sc_hd__nand2_1 _07341_ (.A(_00422_),
    .B(_00432_),
    .Y(_00433_));
 sky130_fd_sc_hd__xnor2_2 _07342_ (.A(_00422_),
    .B(_00432_),
    .Y(_00434_));
 sky130_fd_sc_hd__xnor2_2 _07343_ (.A(_00417_),
    .B(_00434_),
    .Y(_00435_));
 sky130_fd_sc_hd__a22o_1 _07344_ (.A1(_00240_),
    .A2(net42),
    .B1(_00265_),
    .B2(net44),
    .X(_00436_));
 sky130_fd_sc_hd__xor2_1 _07345_ (.A(net94),
    .B(_00436_),
    .X(_00437_));
 sky130_fd_sc_hd__o22a_1 _07346_ (.A1(net130),
    .A2(net46),
    .B1(_00375_),
    .B2(net48),
    .X(_00438_));
 sky130_fd_sc_hd__xnor2_1 _07347_ (.A(net97),
    .B(_00438_),
    .Y(_00439_));
 sky130_fd_sc_hd__nand2_1 _07348_ (.A(_00437_),
    .B(_00439_),
    .Y(_00440_));
 sky130_fd_sc_hd__xor2_1 _07349_ (.A(_00437_),
    .B(_00439_),
    .X(_00441_));
 sky130_fd_sc_hd__a22o_1 _07350_ (.A1(_00226_),
    .A2(net39),
    .B1(net37),
    .B2(_00258_),
    .X(_00442_));
 sky130_fd_sc_hd__xor2_1 _07351_ (.A(net91),
    .B(_00442_),
    .X(_00443_));
 sky130_fd_sc_hd__nand2_1 _07352_ (.A(_00441_),
    .B(_00443_),
    .Y(_00444_));
 sky130_fd_sc_hd__or2_1 _07353_ (.A(_00441_),
    .B(_00443_),
    .X(_00445_));
 sky130_fd_sc_hd__and2_1 _07354_ (.A(_00444_),
    .B(_00445_),
    .X(_00446_));
 sky130_fd_sc_hd__and2b_1 _07355_ (.A_N(_00435_),
    .B(_00446_),
    .X(_00447_));
 sky130_fd_sc_hd__xnor2_2 _07356_ (.A(_00435_),
    .B(_00446_),
    .Y(_00448_));
 sky130_fd_sc_hd__or3_4 _07357_ (.A(reg1_val[26]),
    .B(reg1_val[27]),
    .C(_00234_),
    .X(_00449_));
 sky130_fd_sc_hd__o21ai_2 _07358_ (.A1(_00233_),
    .A2(_00449_),
    .B1(net261),
    .Y(_00450_));
 sky130_fd_sc_hd__xnor2_4 _07359_ (.A(reg1_val[28]),
    .B(_00450_),
    .Y(_00451_));
 sky130_fd_sc_hd__xor2_1 _07360_ (.A(net92),
    .B(_00451_),
    .X(_00452_));
 sky130_fd_sc_hd__xnor2_1 _07361_ (.A(net92),
    .B(_00451_),
    .Y(_00453_));
 sky130_fd_sc_hd__nor2_1 _07362_ (.A(net216),
    .B(net24),
    .Y(_00454_));
 sky130_fd_sc_hd__or3b_1 _07363_ (.A(_00148_),
    .B(_00150_),
    .C_N(_00454_),
    .X(_00455_));
 sky130_fd_sc_hd__o21bai_1 _07364_ (.A1(_00148_),
    .A2(_00150_),
    .B1_N(_00454_),
    .Y(_00456_));
 sky130_fd_sc_hd__nand2_1 _07365_ (.A(_00455_),
    .B(_00456_),
    .Y(_00457_));
 sky130_fd_sc_hd__xnor2_1 _07366_ (.A(_00448_),
    .B(_00457_),
    .Y(_00458_));
 sky130_fd_sc_hd__nor2_1 _07367_ (.A(_00402_),
    .B(_00458_),
    .Y(_00459_));
 sky130_fd_sc_hd__nand2_1 _07368_ (.A(_00402_),
    .B(_00458_),
    .Y(_00460_));
 sky130_fd_sc_hd__and2b_1 _07369_ (.A_N(_00459_),
    .B(_00460_),
    .X(_00461_));
 sky130_fd_sc_hd__xor2_4 _07370_ (.A(_00336_),
    .B(_00461_),
    .X(_00462_));
 sky130_fd_sc_hd__or2_1 _07371_ (.A(_00254_),
    .B(_00269_),
    .X(_00463_));
 sky130_fd_sc_hd__nand2_1 _07372_ (.A(_00270_),
    .B(_00463_),
    .Y(_00464_));
 sky130_fd_sc_hd__nor2_1 _07373_ (.A(_00379_),
    .B(_00381_),
    .Y(_00465_));
 sky130_fd_sc_hd__or2_1 _07374_ (.A(_00382_),
    .B(_00465_),
    .X(_00466_));
 sky130_fd_sc_hd__xnor2_1 _07375_ (.A(_00193_),
    .B(_00194_),
    .Y(_00467_));
 sky130_fd_sc_hd__xnor2_1 _07376_ (.A(_00466_),
    .B(_00467_),
    .Y(_00468_));
 sky130_fd_sc_hd__xnor2_1 _07377_ (.A(_00464_),
    .B(_00468_),
    .Y(_00469_));
 sky130_fd_sc_hd__o22a_1 _07378_ (.A1(net85),
    .A2(net106),
    .B1(net104),
    .B2(net80),
    .X(_00470_));
 sky130_fd_sc_hd__xnor2_2 _07379_ (.A(net135),
    .B(_00470_),
    .Y(_00471_));
 sky130_fd_sc_hd__o22a_1 _07380_ (.A1(net120),
    .A2(net78),
    .B1(net74),
    .B2(_00290_),
    .X(_00472_));
 sky130_fd_sc_hd__xnor2_1 _07381_ (.A(net121),
    .B(_00472_),
    .Y(_00473_));
 sky130_fd_sc_hd__o22a_1 _07382_ (.A1(net86),
    .A2(net76),
    .B1(net72),
    .B2(net82),
    .X(_00474_));
 sky130_fd_sc_hd__xnor2_1 _07383_ (.A(net137),
    .B(_00474_),
    .Y(_00475_));
 sky130_fd_sc_hd__xnor2_1 _07384_ (.A(_00471_),
    .B(_00473_),
    .Y(_00476_));
 sky130_fd_sc_hd__nor2_1 _07385_ (.A(_00475_),
    .B(_00476_),
    .Y(_00477_));
 sky130_fd_sc_hd__o21bai_2 _07386_ (.A1(_00471_),
    .A2(_00473_),
    .B1_N(_00477_),
    .Y(_00478_));
 sky130_fd_sc_hd__and2_1 _07387_ (.A(_00419_),
    .B(_00421_),
    .X(_00479_));
 sky130_fd_sc_hd__nor2_1 _07388_ (.A(_00422_),
    .B(_00479_),
    .Y(_00480_));
 sky130_fd_sc_hd__o22a_1 _07389_ (.A1(net35),
    .A2(net112),
    .B1(net110),
    .B2(net33),
    .X(_00481_));
 sky130_fd_sc_hd__xnor2_1 _07390_ (.A(net125),
    .B(_00481_),
    .Y(_00482_));
 sky130_fd_sc_hd__a22o_1 _07391_ (.A1(_00213_),
    .A2(net29),
    .B1(_00374_),
    .B2(net31),
    .X(_00483_));
 sky130_fd_sc_hd__xnor2_1 _07392_ (.A(net49),
    .B(_00483_),
    .Y(_00484_));
 sky130_fd_sc_hd__and2_1 _07393_ (.A(_00482_),
    .B(_00484_),
    .X(_00485_));
 sky130_fd_sc_hd__nor2_1 _07394_ (.A(_00482_),
    .B(_00484_),
    .Y(_00486_));
 sky130_fd_sc_hd__nor2_1 _07395_ (.A(_00485_),
    .B(_00486_),
    .Y(_00487_));
 sky130_fd_sc_hd__o22a_1 _07396_ (.A1(_00309_),
    .A2(net27),
    .B1(net25),
    .B2(_00313_),
    .X(_00488_));
 sky130_fd_sc_hd__xnor2_1 _07397_ (.A(net88),
    .B(_00488_),
    .Y(_00489_));
 sky130_fd_sc_hd__and2_1 _07398_ (.A(_00487_),
    .B(_00489_),
    .X(_00490_));
 sky130_fd_sc_hd__o21a_1 _07399_ (.A1(_00485_),
    .A2(_00490_),
    .B1(_00480_),
    .X(_00491_));
 sky130_fd_sc_hd__nor3_1 _07400_ (.A(_00480_),
    .B(_00485_),
    .C(_00490_),
    .Y(_00492_));
 sky130_fd_sc_hd__nor2_2 _07401_ (.A(_00491_),
    .B(_00492_),
    .Y(_00493_));
 sky130_fd_sc_hd__xnor2_1 _07402_ (.A(_00478_),
    .B(_00493_),
    .Y(_00494_));
 sky130_fd_sc_hd__nor2_1 _07403_ (.A(_00469_),
    .B(_00494_),
    .Y(_00495_));
 sky130_fd_sc_hd__xor2_2 _07404_ (.A(_06567_),
    .B(_06568_),
    .X(_00496_));
 sky130_fd_sc_hd__and2_1 _07405_ (.A(net94),
    .B(_00496_),
    .X(_00497_));
 sky130_fd_sc_hd__o22a_1 _07406_ (.A1(net288),
    .A2(net65),
    .B1(net59),
    .B2(net237),
    .X(_00498_));
 sky130_fd_sc_hd__xnor2_1 _07407_ (.A(net239),
    .B(_00498_),
    .Y(_00499_));
 sky130_fd_sc_hd__o22a_1 _07408_ (.A1(net152),
    .A2(net57),
    .B1(net149),
    .B2(net63),
    .X(_00500_));
 sky130_fd_sc_hd__xnor2_1 _07409_ (.A(net206),
    .B(_00500_),
    .Y(_00501_));
 sky130_fd_sc_hd__or2_1 _07410_ (.A(_00499_),
    .B(_00501_),
    .X(_00502_));
 sky130_fd_sc_hd__xnor2_2 _07411_ (.A(net94),
    .B(_00496_),
    .Y(_00503_));
 sky130_fd_sc_hd__nor2_1 _07412_ (.A(_00502_),
    .B(_00503_),
    .Y(_00504_));
 sky130_fd_sc_hd__and2_1 _07413_ (.A(_00397_),
    .B(_00398_),
    .X(_00505_));
 sky130_fd_sc_hd__nor2_1 _07414_ (.A(_00399_),
    .B(_00505_),
    .Y(_00506_));
 sky130_fd_sc_hd__o22a_1 _07415_ (.A1(net48),
    .A2(net128),
    .B1(net46),
    .B2(net141),
    .X(_00507_));
 sky130_fd_sc_hd__xor2_1 _07416_ (.A(net97),
    .B(_00507_),
    .X(_00508_));
 sky130_fd_sc_hd__nand2_1 _07417_ (.A(net214),
    .B(net44),
    .Y(_00509_));
 sky130_fd_sc_hd__xor2_1 _07418_ (.A(net94),
    .B(_00509_),
    .X(_00510_));
 sky130_fd_sc_hd__nor2_1 _07419_ (.A(_00508_),
    .B(_00510_),
    .Y(_00511_));
 sky130_fd_sc_hd__and2_1 _07420_ (.A(_00508_),
    .B(_00510_),
    .X(_00512_));
 sky130_fd_sc_hd__or2_1 _07421_ (.A(_00511_),
    .B(_00512_),
    .X(_00513_));
 sky130_fd_sc_hd__a22o_1 _07422_ (.A1(net39),
    .A2(_00265_),
    .B1(net37),
    .B2(_00240_),
    .X(_00514_));
 sky130_fd_sc_hd__xor2_1 _07423_ (.A(net91),
    .B(_00514_),
    .X(_00515_));
 sky130_fd_sc_hd__and2b_1 _07424_ (.A_N(_00513_),
    .B(_00515_),
    .X(_00516_));
 sky130_fd_sc_hd__nor2_2 _07425_ (.A(_00511_),
    .B(_00516_),
    .Y(_00517_));
 sky130_fd_sc_hd__xnor2_1 _07426_ (.A(_00506_),
    .B(_00517_),
    .Y(_00518_));
 sky130_fd_sc_hd__o21ai_2 _07427_ (.A1(_00497_),
    .A2(_00504_),
    .B1(_00518_),
    .Y(_00519_));
 sky130_fd_sc_hd__or3_1 _07428_ (.A(_00497_),
    .B(_00504_),
    .C(_00518_),
    .X(_00520_));
 sky130_fd_sc_hd__and2_2 _07429_ (.A(_00519_),
    .B(_00520_),
    .X(_00521_));
 sky130_fd_sc_hd__nand2_1 _07430_ (.A(_00469_),
    .B(_00494_),
    .Y(_00522_));
 sky130_fd_sc_hd__and2b_1 _07431_ (.A_N(_00495_),
    .B(_00522_),
    .X(_00523_));
 sky130_fd_sc_hd__a21o_1 _07432_ (.A1(_00521_),
    .A2(_00522_),
    .B1(_00495_),
    .X(_00524_));
 sky130_fd_sc_hd__xnor2_2 _07433_ (.A(_00502_),
    .B(_00503_),
    .Y(_00525_));
 sky130_fd_sc_hd__nor2_1 _07434_ (.A(_00487_),
    .B(_00489_),
    .Y(_00526_));
 sky130_fd_sc_hd__nor2_1 _07435_ (.A(_00490_),
    .B(_00526_),
    .Y(_00527_));
 sky130_fd_sc_hd__and2b_1 _07436_ (.A_N(_00525_),
    .B(_00527_),
    .X(_00528_));
 sky130_fd_sc_hd__and2b_1 _07437_ (.A_N(_00515_),
    .B(_00513_),
    .X(_00529_));
 sky130_fd_sc_hd__or2_2 _07438_ (.A(_00516_),
    .B(_00529_),
    .X(_00530_));
 sky130_fd_sc_hd__inv_2 _07439_ (.A(_00530_),
    .Y(_00531_));
 sky130_fd_sc_hd__xnor2_2 _07440_ (.A(_00525_),
    .B(_00527_),
    .Y(_00532_));
 sky130_fd_sc_hd__a21o_1 _07441_ (.A1(_00531_),
    .A2(_00532_),
    .B1(_00528_),
    .X(_00533_));
 sky130_fd_sc_hd__and2_1 _07442_ (.A(_00174_),
    .B(_00192_),
    .X(_00534_));
 sky130_fd_sc_hd__nor2_1 _07443_ (.A(_00193_),
    .B(_00534_),
    .Y(_00535_));
 sky130_fd_sc_hd__o22a_1 _07444_ (.A1(net80),
    .A2(net106),
    .B1(net104),
    .B2(net76),
    .X(_00536_));
 sky130_fd_sc_hd__xnor2_1 _07445_ (.A(net135),
    .B(_00536_),
    .Y(_00537_));
 sky130_fd_sc_hd__o22a_1 _07446_ (.A1(_00290_),
    .A2(net78),
    .B1(net74),
    .B2(net112),
    .X(_00538_));
 sky130_fd_sc_hd__xnor2_1 _07447_ (.A(net121),
    .B(_00538_),
    .Y(_00539_));
 sky130_fd_sc_hd__nor2_1 _07448_ (.A(_00537_),
    .B(_00539_),
    .Y(_00540_));
 sky130_fd_sc_hd__o22a_1 _07449_ (.A1(net120),
    .A2(net82),
    .B1(net73),
    .B2(net86),
    .X(_00541_));
 sky130_fd_sc_hd__xnor2_1 _07450_ (.A(net137),
    .B(_00541_),
    .Y(_00542_));
 sky130_fd_sc_hd__xnor2_1 _07451_ (.A(_00537_),
    .B(_00539_),
    .Y(_00543_));
 sky130_fd_sc_hd__nor2_1 _07452_ (.A(_00542_),
    .B(_00543_),
    .Y(_00544_));
 sky130_fd_sc_hd__o21a_1 _07453_ (.A1(_00540_),
    .A2(_00544_),
    .B1(_00535_),
    .X(_00545_));
 sky130_fd_sc_hd__o22a_1 _07454_ (.A1(net134),
    .A2(net98),
    .B1(net132),
    .B2(net84),
    .X(_00546_));
 sky130_fd_sc_hd__xnor2_1 _07455_ (.A(net181),
    .B(_00546_),
    .Y(_00547_));
 sky130_fd_sc_hd__o22a_1 _07456_ (.A1(net156),
    .A2(net61),
    .B1(net53),
    .B2(net154),
    .X(_00548_));
 sky130_fd_sc_hd__xnor2_1 _07457_ (.A(net207),
    .B(_00548_),
    .Y(_00549_));
 sky130_fd_sc_hd__or2_1 _07458_ (.A(_00547_),
    .B(_00549_),
    .X(_00550_));
 sky130_fd_sc_hd__o22a_1 _07459_ (.A1(net148),
    .A2(net51),
    .B1(net100),
    .B2(net146),
    .X(_00551_));
 sky130_fd_sc_hd__xnor2_1 _07460_ (.A(net202),
    .B(_00551_),
    .Y(_00552_));
 sky130_fd_sc_hd__xnor2_1 _07461_ (.A(_00547_),
    .B(_00549_),
    .Y(_00553_));
 sky130_fd_sc_hd__o21ai_2 _07462_ (.A1(_00552_),
    .A2(_00553_),
    .B1(_00550_),
    .Y(_00554_));
 sky130_fd_sc_hd__nor3_1 _07463_ (.A(_00535_),
    .B(_00540_),
    .C(_00544_),
    .Y(_00555_));
 sky130_fd_sc_hd__or2_1 _07464_ (.A(_00545_),
    .B(_00555_),
    .X(_00556_));
 sky130_fd_sc_hd__and2b_1 _07465_ (.A_N(_00556_),
    .B(_00554_),
    .X(_00557_));
 sky130_fd_sc_hd__nor2_1 _07466_ (.A(_00545_),
    .B(_00557_),
    .Y(_00558_));
 sky130_fd_sc_hd__o21a_1 _07467_ (.A1(_00545_),
    .A2(_00557_),
    .B1(_00533_),
    .X(_00559_));
 sky130_fd_sc_hd__and2_1 _07468_ (.A(_00475_),
    .B(_00476_),
    .X(_00560_));
 sky130_fd_sc_hd__nor2_1 _07469_ (.A(_00477_),
    .B(_00560_),
    .Y(_00561_));
 sky130_fd_sc_hd__a22o_1 _07470_ (.A1(_00294_),
    .A2(_00308_),
    .B1(_00330_),
    .B2(_00283_),
    .X(_00562_));
 sky130_fd_sc_hd__xnor2_1 _07471_ (.A(net124),
    .B(_00562_),
    .Y(_00563_));
 sky130_fd_sc_hd__a22o_1 _07472_ (.A1(_00213_),
    .A2(net31),
    .B1(net29),
    .B2(_00226_),
    .X(_00564_));
 sky130_fd_sc_hd__xnor2_1 _07473_ (.A(net49),
    .B(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__and2_1 _07474_ (.A(_00563_),
    .B(_00565_),
    .X(_00566_));
 sky130_fd_sc_hd__xor2_1 _07475_ (.A(_00563_),
    .B(_00565_),
    .X(_00567_));
 sky130_fd_sc_hd__o22a_1 _07476_ (.A1(_00313_),
    .A2(net27),
    .B1(net25),
    .B2(_00375_),
    .X(_00568_));
 sky130_fd_sc_hd__xnor2_1 _07477_ (.A(net88),
    .B(_00568_),
    .Y(_00569_));
 sky130_fd_sc_hd__and2_1 _07478_ (.A(_00567_),
    .B(_00569_),
    .X(_00570_));
 sky130_fd_sc_hd__o21a_1 _07479_ (.A1(_00566_),
    .A2(_00570_),
    .B1(_00561_),
    .X(_00571_));
 sky130_fd_sc_hd__o22a_1 _07480_ (.A1(net63),
    .A2(net152),
    .B1(net150),
    .B2(net61),
    .X(_00572_));
 sky130_fd_sc_hd__xor2_2 _07481_ (.A(net206),
    .B(_00572_),
    .X(_00573_));
 sky130_fd_sc_hd__o22a_1 _07482_ (.A1(net288),
    .A2(net59),
    .B1(net57),
    .B2(net237),
    .X(_00574_));
 sky130_fd_sc_hd__xnor2_2 _07483_ (.A(net240),
    .B(_00574_),
    .Y(_00575_));
 sky130_fd_sc_hd__o22a_1 _07484_ (.A1(net48),
    .A2(net142),
    .B1(_00264_),
    .B2(net46),
    .X(_00576_));
 sky130_fd_sc_hd__xnor2_1 _07485_ (.A(net97),
    .B(_00576_),
    .Y(_00577_));
 sky130_fd_sc_hd__and3_1 _07486_ (.A(_00573_),
    .B(_00575_),
    .C(_00577_),
    .X(_00578_));
 sky130_fd_sc_hd__a21oi_1 _07487_ (.A1(_00573_),
    .A2(_00575_),
    .B1(_00577_),
    .Y(_00579_));
 sky130_fd_sc_hd__a22o_1 _07488_ (.A1(_00240_),
    .A2(net39),
    .B1(net37),
    .B2(net214),
    .X(_00580_));
 sky130_fd_sc_hd__xor2_1 _07489_ (.A(net91),
    .B(_00580_),
    .X(_00581_));
 sky130_fd_sc_hd__or3b_1 _07490_ (.A(_00578_),
    .B(_00579_),
    .C_N(_00581_),
    .X(_00582_));
 sky130_fd_sc_hd__nand2b_1 _07491_ (.A_N(_00578_),
    .B(_00582_),
    .Y(_00583_));
 sky130_fd_sc_hd__nor3_1 _07492_ (.A(_00561_),
    .B(_00566_),
    .C(_00570_),
    .Y(_00584_));
 sky130_fd_sc_hd__nor2_1 _07493_ (.A(_00571_),
    .B(_00584_),
    .Y(_00585_));
 sky130_fd_sc_hd__a21o_1 _07494_ (.A1(_00583_),
    .A2(_00585_),
    .B1(_00571_),
    .X(_00586_));
 sky130_fd_sc_hd__xnor2_2 _07495_ (.A(_00533_),
    .B(_00558_),
    .Y(_00587_));
 sky130_fd_sc_hd__a21o_1 _07496_ (.A1(_00586_),
    .A2(_00587_),
    .B1(_00559_),
    .X(_00588_));
 sky130_fd_sc_hd__o31ai_4 _07497_ (.A1(_00399_),
    .A2(_00505_),
    .A3(_00517_),
    .B1(_00519_),
    .Y(_00589_));
 sky130_fd_sc_hd__o32a_2 _07498_ (.A1(_00382_),
    .A2(_00465_),
    .A3(_00467_),
    .B1(_00468_),
    .B2(_00464_),
    .X(_00590_));
 sky130_fd_sc_hd__a21oi_4 _07499_ (.A1(_00478_),
    .A2(_00493_),
    .B1(_00491_),
    .Y(_00591_));
 sky130_fd_sc_hd__nor2_1 _07500_ (.A(_00590_),
    .B(_00591_),
    .Y(_00592_));
 sky130_fd_sc_hd__xor2_4 _07501_ (.A(_00590_),
    .B(_00591_),
    .X(_00593_));
 sky130_fd_sc_hd__xor2_2 _07502_ (.A(_00589_),
    .B(_00593_),
    .X(_00594_));
 sky130_fd_sc_hd__xnor2_2 _07503_ (.A(_00588_),
    .B(_00594_),
    .Y(_00595_));
 sky130_fd_sc_hd__nand2b_1 _07504_ (.A_N(_00595_),
    .B(_00524_),
    .Y(_00596_));
 sky130_fd_sc_hd__xnor2_2 _07505_ (.A(_00524_),
    .B(_00595_),
    .Y(_00597_));
 sky130_fd_sc_hd__and2_1 _07506_ (.A(_00462_),
    .B(_00597_),
    .X(_00598_));
 sky130_fd_sc_hd__xor2_1 _07507_ (.A(_00499_),
    .B(_00501_),
    .X(_00599_));
 sky130_fd_sc_hd__o22a_1 _07508_ (.A1(net76),
    .A2(net107),
    .B1(net105),
    .B2(net72),
    .X(_00600_));
 sky130_fd_sc_hd__xnor2_1 _07509_ (.A(net136),
    .B(_00600_),
    .Y(_00601_));
 sky130_fd_sc_hd__o22a_1 _07510_ (.A1(net111),
    .A2(net79),
    .B1(net75),
    .B2(net110),
    .X(_00602_));
 sky130_fd_sc_hd__xnor2_1 _07511_ (.A(net123),
    .B(_00602_),
    .Y(_00603_));
 sky130_fd_sc_hd__or2_1 _07512_ (.A(_00601_),
    .B(_00603_),
    .X(_00604_));
 sky130_fd_sc_hd__o22a_1 _07513_ (.A1(net119),
    .A2(net87),
    .B1(net83),
    .B2(net117),
    .X(_00605_));
 sky130_fd_sc_hd__xnor2_1 _07514_ (.A(net138),
    .B(_00605_),
    .Y(_00606_));
 sky130_fd_sc_hd__xnor2_1 _07515_ (.A(_00601_),
    .B(_00603_),
    .Y(_00607_));
 sky130_fd_sc_hd__o21ai_1 _07516_ (.A1(_00606_),
    .A2(_00607_),
    .B1(_00604_),
    .Y(_00608_));
 sky130_fd_sc_hd__nand2_1 _07517_ (.A(_00599_),
    .B(_00608_),
    .Y(_00609_));
 sky130_fd_sc_hd__xnor2_1 _07518_ (.A(_00599_),
    .B(_00608_),
    .Y(_00610_));
 sky130_fd_sc_hd__o22a_1 _07519_ (.A1(net156),
    .A2(net53),
    .B1(net51),
    .B2(net154),
    .X(_00611_));
 sky130_fd_sc_hd__xnor2_1 _07520_ (.A(net207),
    .B(_00611_),
    .Y(_00612_));
 sky130_fd_sc_hd__o22a_1 _07521_ (.A1(net133),
    .A2(net84),
    .B1(net80),
    .B2(net131),
    .X(_00613_));
 sky130_fd_sc_hd__xnor2_1 _07522_ (.A(net180),
    .B(_00613_),
    .Y(_00614_));
 sky130_fd_sc_hd__or2_1 _07523_ (.A(_00612_),
    .B(_00614_),
    .X(_00615_));
 sky130_fd_sc_hd__o22a_1 _07524_ (.A1(net148),
    .A2(net100),
    .B1(net98),
    .B2(net146),
    .X(_00616_));
 sky130_fd_sc_hd__xnor2_1 _07525_ (.A(net202),
    .B(_00616_),
    .Y(_00617_));
 sky130_fd_sc_hd__xnor2_1 _07526_ (.A(_00612_),
    .B(_00614_),
    .Y(_00618_));
 sky130_fd_sc_hd__or2_1 _07527_ (.A(_00617_),
    .B(_00618_),
    .X(_00619_));
 sky130_fd_sc_hd__a21o_1 _07528_ (.A1(_00615_),
    .A2(_00619_),
    .B1(_00610_),
    .X(_00620_));
 sky130_fd_sc_hd__nand2_1 _07529_ (.A(_00609_),
    .B(_00620_),
    .Y(_00621_));
 sky130_fd_sc_hd__and2_1 _07530_ (.A(_00542_),
    .B(_00543_),
    .X(_00622_));
 sky130_fd_sc_hd__nor2_1 _07531_ (.A(_00544_),
    .B(_00622_),
    .Y(_00623_));
 sky130_fd_sc_hd__o21bai_1 _07532_ (.A1(_00578_),
    .A2(_00579_),
    .B1_N(_00581_),
    .Y(_00624_));
 sky130_fd_sc_hd__nand3_1 _07533_ (.A(_00582_),
    .B(_00623_),
    .C(_00624_),
    .Y(_00625_));
 sky130_fd_sc_hd__nor2_1 _07534_ (.A(_00567_),
    .B(_00569_),
    .Y(_00626_));
 sky130_fd_sc_hd__nor2_1 _07535_ (.A(_00570_),
    .B(_00626_),
    .Y(_00627_));
 sky130_fd_sc_hd__a21o_1 _07536_ (.A1(_00582_),
    .A2(_00624_),
    .B1(_00623_),
    .X(_00628_));
 sky130_fd_sc_hd__nand3_1 _07537_ (.A(_00625_),
    .B(_00627_),
    .C(_00628_),
    .Y(_00629_));
 sky130_fd_sc_hd__a21boi_2 _07538_ (.A1(_00627_),
    .A2(_00628_),
    .B1_N(_00625_),
    .Y(_00630_));
 sky130_fd_sc_hd__a21o_1 _07539_ (.A1(_00609_),
    .A2(_00620_),
    .B1(_00630_),
    .X(_00631_));
 sky130_fd_sc_hd__xor2_1 _07540_ (.A(_00552_),
    .B(_00553_),
    .X(_00632_));
 sky130_fd_sc_hd__a22o_1 _07541_ (.A1(_00283_),
    .A2(_00308_),
    .B1(net113),
    .B2(_00294_),
    .X(_00633_));
 sky130_fd_sc_hd__xnor2_2 _07542_ (.A(net124),
    .B(_00633_),
    .Y(_00634_));
 sky130_fd_sc_hd__a22o_1 _07543_ (.A1(_00226_),
    .A2(net31),
    .B1(net29),
    .B2(_00258_),
    .X(_00635_));
 sky130_fd_sc_hd__xnor2_2 _07544_ (.A(net49),
    .B(_00635_),
    .Y(_00636_));
 sky130_fd_sc_hd__and2_1 _07545_ (.A(_00634_),
    .B(_00636_),
    .X(_00637_));
 sky130_fd_sc_hd__xor2_2 _07546_ (.A(_00634_),
    .B(_00636_),
    .X(_00638_));
 sky130_fd_sc_hd__o22a_1 _07547_ (.A1(net130),
    .A2(net25),
    .B1(_00375_),
    .B2(net27),
    .X(_00639_));
 sky130_fd_sc_hd__xnor2_2 _07548_ (.A(net88),
    .B(_00639_),
    .Y(_00640_));
 sky130_fd_sc_hd__and2_1 _07549_ (.A(_00638_),
    .B(_00640_),
    .X(_00641_));
 sky130_fd_sc_hd__o21a_1 _07550_ (.A1(_00637_),
    .A2(_00641_),
    .B1(_00632_),
    .X(_00642_));
 sky130_fd_sc_hd__nand2_1 _07551_ (.A(net214),
    .B(net39),
    .Y(_00643_));
 sky130_fd_sc_hd__o22a_1 _07552_ (.A1(net46),
    .A2(net144),
    .B1(_00264_),
    .B2(net48),
    .X(_00644_));
 sky130_fd_sc_hd__xor2_1 _07553_ (.A(net97),
    .B(_00644_),
    .X(_00645_));
 sky130_fd_sc_hd__and3_1 _07554_ (.A(net214),
    .B(net39),
    .C(_00645_),
    .X(_00646_));
 sky130_fd_sc_hd__a21oi_1 _07555_ (.A1(net214),
    .A2(net39),
    .B1(net91),
    .Y(_00647_));
 sky130_fd_sc_hd__nor3_1 _07556_ (.A(_00632_),
    .B(_00637_),
    .C(_00641_),
    .Y(_00648_));
 sky130_fd_sc_hd__nor4_1 _07557_ (.A(_00642_),
    .B(_00646_),
    .C(_00647_),
    .D(_00648_),
    .Y(_00649_));
 sky130_fd_sc_hd__or2_1 _07558_ (.A(_00642_),
    .B(_00649_),
    .X(_00650_));
 sky130_fd_sc_hd__xnor2_2 _07559_ (.A(_00621_),
    .B(_00630_),
    .Y(_00651_));
 sky130_fd_sc_hd__a21bo_1 _07560_ (.A1(_00650_),
    .A2(_00651_),
    .B1_N(_00631_),
    .X(_00652_));
 sky130_fd_sc_hd__xor2_2 _07561_ (.A(_00586_),
    .B(_00587_),
    .X(_00653_));
 sky130_fd_sc_hd__xnor2_2 _07562_ (.A(_00530_),
    .B(_00532_),
    .Y(_00654_));
 sky130_fd_sc_hd__xnor2_2 _07563_ (.A(_00554_),
    .B(_00556_),
    .Y(_00655_));
 sky130_fd_sc_hd__nand2_1 _07564_ (.A(_00654_),
    .B(_00655_),
    .Y(_00656_));
 sky130_fd_sc_hd__xnor2_2 _07565_ (.A(_00654_),
    .B(_00655_),
    .Y(_00657_));
 sky130_fd_sc_hd__xnor2_1 _07566_ (.A(_00583_),
    .B(_00585_),
    .Y(_00658_));
 sky130_fd_sc_hd__o21ai_2 _07567_ (.A1(_00657_),
    .A2(_00658_),
    .B1(_00656_),
    .Y(_00659_));
 sky130_fd_sc_hd__xnor2_2 _07568_ (.A(_00652_),
    .B(_00653_),
    .Y(_00660_));
 sky130_fd_sc_hd__nand2b_1 _07569_ (.A_N(_00660_),
    .B(_00659_),
    .Y(_00661_));
 sky130_fd_sc_hd__a21bo_2 _07570_ (.A1(_00652_),
    .A2(_00653_),
    .B1_N(_00661_),
    .X(_00662_));
 sky130_fd_sc_hd__xor2_4 _07571_ (.A(_00462_),
    .B(_00597_),
    .X(_00663_));
 sky130_fd_sc_hd__a21oi_4 _07572_ (.A1(_00662_),
    .A2(_00663_),
    .B1(_00598_),
    .Y(_00664_));
 sky130_fd_sc_hd__a21bo_2 _07573_ (.A1(_00588_),
    .A2(_00594_),
    .B1_N(_00596_),
    .X(_00665_));
 sky130_fd_sc_hd__o21a_2 _07574_ (.A1(_00417_),
    .A2(_00434_),
    .B1(_00433_),
    .X(_00666_));
 sky130_fd_sc_hd__o22a_1 _07575_ (.A1(net120),
    .A2(net33),
    .B1(net72),
    .B2(net35),
    .X(_00667_));
 sky130_fd_sc_hd__xnor2_1 _07576_ (.A(net125),
    .B(_00667_),
    .Y(_00668_));
 sky130_fd_sc_hd__a22o_1 _07577_ (.A1(_00308_),
    .A2(net29),
    .B1(_00330_),
    .B2(net31),
    .X(_00669_));
 sky130_fd_sc_hd__xnor2_1 _07578_ (.A(net49),
    .B(_00669_),
    .Y(_00670_));
 sky130_fd_sc_hd__and2_1 _07579_ (.A(_00668_),
    .B(_00670_),
    .X(_00671_));
 sky130_fd_sc_hd__nor2_1 _07580_ (.A(_00668_),
    .B(_00670_),
    .Y(_00672_));
 sky130_fd_sc_hd__nor2_1 _07581_ (.A(_00671_),
    .B(_00672_),
    .Y(_00673_));
 sky130_fd_sc_hd__o22a_1 _07582_ (.A1(_00290_),
    .A2(net27),
    .B1(net112),
    .B2(net25),
    .X(_00674_));
 sky130_fd_sc_hd__xnor2_1 _07583_ (.A(net88),
    .B(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hd__xor2_1 _07584_ (.A(_00673_),
    .B(_00675_),
    .X(_00676_));
 sky130_fd_sc_hd__o31a_2 _07585_ (.A1(reg1_val[28]),
    .A2(_00233_),
    .A3(_00449_),
    .B1(net261),
    .X(_00677_));
 sky130_fd_sc_hd__xor2_4 _07586_ (.A(reg1_val[29]),
    .B(_00677_),
    .X(_00678_));
 sky130_fd_sc_hd__xnor2_1 _07587_ (.A(reg1_val[29]),
    .B(_00677_),
    .Y(_00679_));
 sky130_fd_sc_hd__or2_1 _07588_ (.A(_00454_),
    .B(_00678_),
    .X(_00680_));
 sky130_fd_sc_hd__and3_1 _07589_ (.A(_00455_),
    .B(_00676_),
    .C(_00680_),
    .X(_00681_));
 sky130_fd_sc_hd__a21oi_2 _07590_ (.A1(_00455_),
    .A2(_00680_),
    .B1(_00676_),
    .Y(_00682_));
 sky130_fd_sc_hd__nor2_2 _07591_ (.A(_00681_),
    .B(_00682_),
    .Y(_00683_));
 sky130_fd_sc_hd__xnor2_4 _07592_ (.A(_00666_),
    .B(_00683_),
    .Y(_00684_));
 sky130_fd_sc_hd__a21o_1 _07593_ (.A1(_00428_),
    .A2(_00431_),
    .B1(_00427_),
    .X(_00685_));
 sky130_fd_sc_hd__a21o_1 _07594_ (.A1(net92),
    .A2(_00451_),
    .B1(_00678_),
    .X(_00686_));
 sky130_fd_sc_hd__o21ai_2 _07595_ (.A1(net92),
    .A2(_00451_),
    .B1(_00678_),
    .Y(_00687_));
 sky130_fd_sc_hd__nand2_1 _07596_ (.A(_00686_),
    .B(_00687_),
    .Y(_00688_));
 sky130_fd_sc_hd__o22a_1 _07597_ (.A1(net144),
    .A2(net24),
    .B1(net16),
    .B2(net216),
    .X(_00689_));
 sky130_fd_sc_hd__xnor2_1 _07598_ (.A(_00678_),
    .B(_00689_),
    .Y(_00690_));
 sky130_fd_sc_hd__xor2_1 _07599_ (.A(_00685_),
    .B(_00690_),
    .X(_00691_));
 sky130_fd_sc_hd__o21a_1 _07600_ (.A1(_00414_),
    .A2(_00416_),
    .B1(_00691_),
    .X(_00692_));
 sky130_fd_sc_hd__nor3_1 _07601_ (.A(_00414_),
    .B(_00416_),
    .C(_00691_),
    .Y(_00693_));
 sky130_fd_sc_hd__nor2_1 _07602_ (.A(_00692_),
    .B(_00693_),
    .Y(_00694_));
 sky130_fd_sc_hd__o22a_1 _07603_ (.A1(net68),
    .A2(net150),
    .B1(net56),
    .B2(net152),
    .X(_00695_));
 sky130_fd_sc_hd__xnor2_2 _07604_ (.A(net206),
    .B(_00695_),
    .Y(_00696_));
 sky130_fd_sc_hd__a211o_4 _07605_ (.A1(_05013_),
    .A2(_00139_),
    .B1(net183),
    .C1(_04937_),
    .X(_00697_));
 sky130_fd_sc_hd__o211ai_4 _07606_ (.A1(net183),
    .A2(_00139_),
    .B1(_00406_),
    .C1(_04937_),
    .Y(_00698_));
 sky130_fd_sc_hd__and2_4 _07607_ (.A(_00697_),
    .B(_00698_),
    .X(_00699_));
 sky130_fd_sc_hd__nand2_4 _07608_ (.A(_00697_),
    .B(_00698_),
    .Y(_00700_));
 sky130_fd_sc_hd__a22o_1 _07609_ (.A1(_06519_),
    .A2(_00408_),
    .B1(_00700_),
    .B2(net292),
    .X(_00701_));
 sky130_fd_sc_hd__xnor2_4 _07610_ (.A(_06493_),
    .B(_00701_),
    .Y(_00702_));
 sky130_fd_sc_hd__o22a_1 _07611_ (.A1(net65),
    .A2(net156),
    .B1(net154),
    .B2(net59),
    .X(_00703_));
 sky130_fd_sc_hd__xnor2_2 _07612_ (.A(net207),
    .B(_00703_),
    .Y(_00704_));
 sky130_fd_sc_hd__or2_1 _07613_ (.A(_00702_),
    .B(_00704_),
    .X(_00705_));
 sky130_fd_sc_hd__xnor2_2 _07614_ (.A(_00702_),
    .B(_00704_),
    .Y(_00706_));
 sky130_fd_sc_hd__xor2_2 _07615_ (.A(_00696_),
    .B(_00706_),
    .X(_00707_));
 sky130_fd_sc_hd__o22a_1 _07616_ (.A1(net51),
    .A2(net106),
    .B1(net104),
    .B2(net100),
    .X(_00708_));
 sky130_fd_sc_hd__xnor2_2 _07617_ (.A(net135),
    .B(_00708_),
    .Y(_00709_));
 sky130_fd_sc_hd__o22a_1 _07618_ (.A1(net57),
    .A2(net148),
    .B1(net146),
    .B2(net63),
    .X(_00710_));
 sky130_fd_sc_hd__xnor2_2 _07619_ (.A(net202),
    .B(_00710_),
    .Y(_00711_));
 sky130_fd_sc_hd__xor2_2 _07620_ (.A(_00709_),
    .B(_00711_),
    .X(_00712_));
 sky130_fd_sc_hd__o22a_1 _07621_ (.A1(net61),
    .A2(net134),
    .B1(net132),
    .B2(net53),
    .X(_00713_));
 sky130_fd_sc_hd__xnor2_2 _07622_ (.A(net181),
    .B(_00713_),
    .Y(_00714_));
 sky130_fd_sc_hd__nand2b_1 _07623_ (.A_N(_00714_),
    .B(_00712_),
    .Y(_00715_));
 sky130_fd_sc_hd__xnor2_2 _07624_ (.A(_00712_),
    .B(_00714_),
    .Y(_00716_));
 sky130_fd_sc_hd__and2_1 _07625_ (.A(_00369_),
    .B(_00716_),
    .X(_00717_));
 sky130_fd_sc_hd__xnor2_2 _07626_ (.A(_00369_),
    .B(_00716_),
    .Y(_00718_));
 sky130_fd_sc_hd__inv_2 _07627_ (.A(_00718_),
    .Y(_00719_));
 sky130_fd_sc_hd__xor2_1 _07628_ (.A(_00707_),
    .B(_00718_),
    .X(_00720_));
 sky130_fd_sc_hd__a22o_1 _07629_ (.A1(net44),
    .A2(_00258_),
    .B1(_00265_),
    .B2(net42),
    .X(_00721_));
 sky130_fd_sc_hd__xor2_1 _07630_ (.A(net94),
    .B(_00721_),
    .X(_00722_));
 sky130_fd_sc_hd__o22a_1 _07631_ (.A1(net48),
    .A2(_00313_),
    .B1(net108),
    .B2(net46),
    .X(_00723_));
 sky130_fd_sc_hd__xnor2_1 _07632_ (.A(net97),
    .B(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hd__nand2_1 _07633_ (.A(_00722_),
    .B(_00724_),
    .Y(_00725_));
 sky130_fd_sc_hd__or2_1 _07634_ (.A(_00722_),
    .B(_00724_),
    .X(_00726_));
 sky130_fd_sc_hd__and2_1 _07635_ (.A(_00725_),
    .B(_00726_),
    .X(_00727_));
 sky130_fd_sc_hd__a22o_1 _07636_ (.A1(_00213_),
    .A2(net39),
    .B1(net37),
    .B2(_00226_),
    .X(_00728_));
 sky130_fd_sc_hd__xor2_1 _07637_ (.A(net91),
    .B(_00728_),
    .X(_00729_));
 sky130_fd_sc_hd__nand2_1 _07638_ (.A(_00727_),
    .B(_00729_),
    .Y(_00730_));
 sky130_fd_sc_hd__or2_1 _07639_ (.A(_00727_),
    .B(_00729_),
    .X(_00731_));
 sky130_fd_sc_hd__and2_1 _07640_ (.A(_00730_),
    .B(_00731_),
    .X(_00732_));
 sky130_fd_sc_hd__and2b_1 _07641_ (.A_N(_00720_),
    .B(_00732_),
    .X(_00733_));
 sky130_fd_sc_hd__xnor2_1 _07642_ (.A(_00720_),
    .B(_00732_),
    .Y(_00734_));
 sky130_fd_sc_hd__nand2_1 _07643_ (.A(_00694_),
    .B(_00734_),
    .Y(_00735_));
 sky130_fd_sc_hd__or2_1 _07644_ (.A(_00694_),
    .B(_00734_),
    .X(_00736_));
 sky130_fd_sc_hd__nand2_1 _07645_ (.A(_00735_),
    .B(_00736_),
    .Y(_00737_));
 sky130_fd_sc_hd__a21oi_2 _07646_ (.A1(_00319_),
    .A2(_00332_),
    .B1(_00317_),
    .Y(_00738_));
 sky130_fd_sc_hd__o22a_1 _07647_ (.A1(net98),
    .A2(net86),
    .B1(net84),
    .B2(net82),
    .X(_00739_));
 sky130_fd_sc_hd__xnor2_1 _07648_ (.A(net137),
    .B(_00739_),
    .Y(_00740_));
 sky130_fd_sc_hd__o22a_1 _07649_ (.A1(net80),
    .A2(net78),
    .B1(net76),
    .B2(net74),
    .X(_00741_));
 sky130_fd_sc_hd__xnor2_1 _07650_ (.A(net121),
    .B(_00741_),
    .Y(_00742_));
 sky130_fd_sc_hd__nor2_1 _07651_ (.A(_00740_),
    .B(_00742_),
    .Y(_00743_));
 sky130_fd_sc_hd__and2_1 _07652_ (.A(_00740_),
    .B(_00742_),
    .X(_00744_));
 sky130_fd_sc_hd__or2_1 _07653_ (.A(_00743_),
    .B(_00744_),
    .X(_00745_));
 sky130_fd_sc_hd__a21oi_2 _07654_ (.A1(_00440_),
    .A2(_00444_),
    .B1(_00745_),
    .Y(_00746_));
 sky130_fd_sc_hd__and3_1 _07655_ (.A(_00440_),
    .B(_00444_),
    .C(_00745_),
    .X(_00747_));
 sky130_fd_sc_hd__nor2_1 _07656_ (.A(_00746_),
    .B(_00747_),
    .Y(_00748_));
 sky130_fd_sc_hd__and2b_1 _07657_ (.A_N(_00738_),
    .B(_00748_),
    .X(_00749_));
 sky130_fd_sc_hd__xnor2_2 _07658_ (.A(_00738_),
    .B(_00748_),
    .Y(_00750_));
 sky130_fd_sc_hd__xnor2_2 _07659_ (.A(_00737_),
    .B(_00750_),
    .Y(_00751_));
 sky130_fd_sc_hd__xor2_4 _07660_ (.A(_00684_),
    .B(_00751_),
    .X(_00752_));
 sky130_fd_sc_hd__a21o_1 _07661_ (.A1(_00336_),
    .A2(_00460_),
    .B1(_00459_),
    .X(_00753_));
 sky130_fd_sc_hd__o21ai_4 _07662_ (.A1(_00272_),
    .A2(_00333_),
    .B1(_00335_),
    .Y(_00754_));
 sky130_fd_sc_hd__or2_2 _07663_ (.A(_00383_),
    .B(_00401_),
    .X(_00755_));
 sky130_fd_sc_hd__a21oi_2 _07664_ (.A1(_00448_),
    .A2(_00457_),
    .B1(_00447_),
    .Y(_00756_));
 sky130_fd_sc_hd__o21ba_1 _07665_ (.A1(_00383_),
    .A2(_00401_),
    .B1_N(_00756_),
    .X(_00757_));
 sky130_fd_sc_hd__xnor2_4 _07666_ (.A(_00755_),
    .B(_00756_),
    .Y(_00758_));
 sky130_fd_sc_hd__xnor2_4 _07667_ (.A(_00754_),
    .B(_00758_),
    .Y(_00759_));
 sky130_fd_sc_hd__a21oi_4 _07668_ (.A1(_00589_),
    .A2(_00593_),
    .B1(_00592_),
    .Y(_00760_));
 sky130_fd_sc_hd__xnor2_2 _07669_ (.A(_00759_),
    .B(_00760_),
    .Y(_00761_));
 sky130_fd_sc_hd__nand2b_1 _07670_ (.A_N(_00761_),
    .B(_00753_),
    .Y(_00762_));
 sky130_fd_sc_hd__xnor2_2 _07671_ (.A(_00753_),
    .B(_00761_),
    .Y(_00763_));
 sky130_fd_sc_hd__and2_1 _07672_ (.A(_00752_),
    .B(_00763_),
    .X(_00764_));
 sky130_fd_sc_hd__xor2_4 _07673_ (.A(_00752_),
    .B(_00763_),
    .X(_00765_));
 sky130_fd_sc_hd__xnor2_4 _07674_ (.A(_00665_),
    .B(_00765_),
    .Y(_00766_));
 sky130_fd_sc_hd__or2_1 _07675_ (.A(_00664_),
    .B(_00766_),
    .X(_00767_));
 sky130_fd_sc_hd__xnor2_4 _07676_ (.A(_00664_),
    .B(_00766_),
    .Y(_00768_));
 sky130_fd_sc_hd__xnor2_4 _07677_ (.A(_00662_),
    .B(_00663_),
    .Y(_00769_));
 sky130_fd_sc_hd__xor2_4 _07678_ (.A(_00521_),
    .B(_00523_),
    .X(_00770_));
 sky130_fd_sc_hd__xnor2_2 _07679_ (.A(_00659_),
    .B(_00660_),
    .Y(_00771_));
 sky130_fd_sc_hd__and2_1 _07680_ (.A(_00770_),
    .B(_00771_),
    .X(_00772_));
 sky130_fd_sc_hd__xnor2_2 _07681_ (.A(_00650_),
    .B(_00651_),
    .Y(_00773_));
 sky130_fd_sc_hd__xor2_1 _07682_ (.A(_00573_),
    .B(_00575_),
    .X(_00774_));
 sky130_fd_sc_hd__o22a_1 _07683_ (.A1(net72),
    .A2(net107),
    .B1(net105),
    .B2(net119),
    .X(_00775_));
 sky130_fd_sc_hd__xnor2_2 _07684_ (.A(net136),
    .B(_00775_),
    .Y(_00776_));
 sky130_fd_sc_hd__o22a_1 _07685_ (.A1(net148),
    .A2(net98),
    .B1(net84),
    .B2(net145),
    .X(_00777_));
 sky130_fd_sc_hd__xnor2_2 _07686_ (.A(net201),
    .B(_00777_),
    .Y(_00778_));
 sky130_fd_sc_hd__nor2_1 _07687_ (.A(_00776_),
    .B(_00778_),
    .Y(_00779_));
 sky130_fd_sc_hd__xor2_2 _07688_ (.A(_00776_),
    .B(_00778_),
    .X(_00780_));
 sky130_fd_sc_hd__o22a_1 _07689_ (.A1(net133),
    .A2(net80),
    .B1(net76),
    .B2(net131),
    .X(_00781_));
 sky130_fd_sc_hd__xnor2_2 _07690_ (.A(net182),
    .B(_00781_),
    .Y(_00782_));
 sky130_fd_sc_hd__inv_2 _07691_ (.A(_00782_),
    .Y(_00783_));
 sky130_fd_sc_hd__a21oi_1 _07692_ (.A1(_00780_),
    .A2(_00783_),
    .B1(_00779_),
    .Y(_00784_));
 sky130_fd_sc_hd__and2b_1 _07693_ (.A_N(_00784_),
    .B(_00774_),
    .X(_00785_));
 sky130_fd_sc_hd__o22a_1 _07694_ (.A1(_06520_),
    .A2(net63),
    .B1(net57),
    .B2(net288),
    .X(_00786_));
 sky130_fd_sc_hd__xnor2_1 _07695_ (.A(net239),
    .B(_00786_),
    .Y(_00787_));
 sky130_fd_sc_hd__o22a_1 _07696_ (.A1(net156),
    .A2(net51),
    .B1(net100),
    .B2(net154),
    .X(_00788_));
 sky130_fd_sc_hd__xnor2_1 _07697_ (.A(net207),
    .B(_00788_),
    .Y(_00789_));
 sky130_fd_sc_hd__or2_1 _07698_ (.A(_00787_),
    .B(_00789_),
    .X(_00790_));
 sky130_fd_sc_hd__o22a_1 _07699_ (.A1(net61),
    .A2(net152),
    .B1(net150),
    .B2(net53),
    .X(_00791_));
 sky130_fd_sc_hd__xnor2_1 _07700_ (.A(net204),
    .B(_00791_),
    .Y(_00792_));
 sky130_fd_sc_hd__xnor2_1 _07701_ (.A(_00787_),
    .B(_00789_),
    .Y(_00793_));
 sky130_fd_sc_hd__o21ai_1 _07702_ (.A1(_00792_),
    .A2(_00793_),
    .B1(_00790_),
    .Y(_00794_));
 sky130_fd_sc_hd__xnor2_1 _07703_ (.A(_00774_),
    .B(_00784_),
    .Y(_00795_));
 sky130_fd_sc_hd__a21o_1 _07704_ (.A1(_00794_),
    .A2(_00795_),
    .B1(_00785_),
    .X(_00796_));
 sky130_fd_sc_hd__xnor2_1 _07705_ (.A(_00606_),
    .B(_00607_),
    .Y(_00797_));
 sky130_fd_sc_hd__xnor2_1 _07706_ (.A(_00643_),
    .B(_00645_),
    .Y(_00798_));
 sky130_fd_sc_hd__nor2_1 _07707_ (.A(_00797_),
    .B(_00798_),
    .Y(_00799_));
 sky130_fd_sc_hd__xor2_2 _07708_ (.A(_00638_),
    .B(_00640_),
    .X(_00800_));
 sky130_fd_sc_hd__xor2_1 _07709_ (.A(_00797_),
    .B(_00798_),
    .X(_00801_));
 sky130_fd_sc_hd__a21o_1 _07710_ (.A1(_00800_),
    .A2(_00801_),
    .B1(_00799_),
    .X(_00802_));
 sky130_fd_sc_hd__nand2_1 _07711_ (.A(_00796_),
    .B(_00802_),
    .Y(_00803_));
 sky130_fd_sc_hd__o22a_1 _07712_ (.A1(net117),
    .A2(net87),
    .B1(net83),
    .B2(net111),
    .X(_00804_));
 sky130_fd_sc_hd__xnor2_2 _07713_ (.A(net138),
    .B(_00804_),
    .Y(_00805_));
 sky130_fd_sc_hd__a22o_1 _07714_ (.A1(_00283_),
    .A2(net113),
    .B1(_00374_),
    .B2(_00294_),
    .X(_00806_));
 sky130_fd_sc_hd__xnor2_2 _07715_ (.A(net125),
    .B(_00806_),
    .Y(_00807_));
 sky130_fd_sc_hd__or2_1 _07716_ (.A(_00805_),
    .B(_00807_),
    .X(_00808_));
 sky130_fd_sc_hd__xnor2_2 _07717_ (.A(_00805_),
    .B(_00807_),
    .Y(_00809_));
 sky130_fd_sc_hd__o22a_1 _07718_ (.A1(net109),
    .A2(net79),
    .B1(net75),
    .B2(net115),
    .X(_00810_));
 sky130_fd_sc_hd__xnor2_2 _07719_ (.A(net123),
    .B(_00810_),
    .Y(_00811_));
 sky130_fd_sc_hd__o21ai_1 _07720_ (.A1(_00809_),
    .A2(_00811_),
    .B1(_00808_),
    .Y(_00812_));
 sky130_fd_sc_hd__xor2_1 _07721_ (.A(_00617_),
    .B(_00618_),
    .X(_00813_));
 sky130_fd_sc_hd__and2_1 _07722_ (.A(_00812_),
    .B(_00813_),
    .X(_00814_));
 sky130_fd_sc_hd__o22a_1 _07723_ (.A1(net129),
    .A2(net27),
    .B1(net25),
    .B2(net127),
    .X(_00815_));
 sky130_fd_sc_hd__xnor2_2 _07724_ (.A(net88),
    .B(_00815_),
    .Y(_00816_));
 sky130_fd_sc_hd__a22o_1 _07725_ (.A1(_00258_),
    .A2(net31),
    .B1(net29),
    .B2(_00265_),
    .X(_00817_));
 sky130_fd_sc_hd__xnor2_2 _07726_ (.A(net49),
    .B(_00817_),
    .Y(_00818_));
 sky130_fd_sc_hd__and2_1 _07727_ (.A(_00816_),
    .B(_00818_),
    .X(_00819_));
 sky130_fd_sc_hd__xor2_1 _07728_ (.A(_00812_),
    .B(_00813_),
    .X(_00820_));
 sky130_fd_sc_hd__a21oi_1 _07729_ (.A1(_00819_),
    .A2(_00820_),
    .B1(_00814_),
    .Y(_00821_));
 sky130_fd_sc_hd__nor2_1 _07730_ (.A(_00796_),
    .B(_00802_),
    .Y(_00822_));
 sky130_fd_sc_hd__xor2_1 _07731_ (.A(_00796_),
    .B(_00802_),
    .X(_00823_));
 sky130_fd_sc_hd__o21a_1 _07732_ (.A1(_00821_),
    .A2(_00822_),
    .B1(_00803_),
    .X(_00824_));
 sky130_fd_sc_hd__or2_1 _07733_ (.A(_00773_),
    .B(_00824_),
    .X(_00825_));
 sky130_fd_sc_hd__nand3_1 _07734_ (.A(_00610_),
    .B(_00615_),
    .C(_00619_),
    .Y(_00826_));
 sky130_fd_sc_hd__and2_1 _07735_ (.A(_00620_),
    .B(_00826_),
    .X(_00827_));
 sky130_fd_sc_hd__a21o_1 _07736_ (.A1(_00625_),
    .A2(_00628_),
    .B1(_00627_),
    .X(_00828_));
 sky130_fd_sc_hd__and3_1 _07737_ (.A(_00629_),
    .B(_00827_),
    .C(_00828_),
    .X(_00829_));
 sky130_fd_sc_hd__a21oi_1 _07738_ (.A1(_00629_),
    .A2(_00828_),
    .B1(_00827_),
    .Y(_00830_));
 sky130_fd_sc_hd__nor2_1 _07739_ (.A(_00829_),
    .B(_00830_),
    .Y(_00831_));
 sky130_fd_sc_hd__o22a_1 _07740_ (.A1(_00646_),
    .A2(_00647_),
    .B1(_00648_),
    .B2(_00642_),
    .X(_00832_));
 sky130_fd_sc_hd__or2_1 _07741_ (.A(_00649_),
    .B(_00832_),
    .X(_00833_));
 sky130_fd_sc_hd__o21ba_1 _07742_ (.A1(_00830_),
    .A2(_00833_),
    .B1_N(_00829_),
    .X(_00834_));
 sky130_fd_sc_hd__xnor2_2 _07743_ (.A(_00773_),
    .B(_00824_),
    .Y(_00835_));
 sky130_fd_sc_hd__o21ai_4 _07744_ (.A1(_00834_),
    .A2(_00835_),
    .B1(_00825_),
    .Y(_00836_));
 sky130_fd_sc_hd__xor2_4 _07745_ (.A(_00770_),
    .B(_00771_),
    .X(_00837_));
 sky130_fd_sc_hd__a21oi_4 _07746_ (.A1(_00836_),
    .A2(_00837_),
    .B1(_00772_),
    .Y(_00838_));
 sky130_fd_sc_hd__nand2_1 _07747_ (.A(_00769_),
    .B(_00838_),
    .Y(_00839_));
 sky130_fd_sc_hd__xor2_1 _07748_ (.A(_00657_),
    .B(_00658_),
    .X(_00840_));
 sky130_fd_sc_hd__xor2_1 _07749_ (.A(_00834_),
    .B(_00835_),
    .X(_00841_));
 sky130_fd_sc_hd__xnor2_1 _07750_ (.A(_00821_),
    .B(_00823_),
    .Y(_00842_));
 sky130_fd_sc_hd__xor2_2 _07751_ (.A(_00816_),
    .B(_00818_),
    .X(_00843_));
 sky130_fd_sc_hd__xnor2_2 _07752_ (.A(_00780_),
    .B(_00782_),
    .Y(_00844_));
 sky130_fd_sc_hd__nand2_1 _07753_ (.A(_00843_),
    .B(_00844_),
    .Y(_00845_));
 sky130_fd_sc_hd__xnor2_2 _07754_ (.A(_00843_),
    .B(_00844_),
    .Y(_00846_));
 sky130_fd_sc_hd__xnor2_2 _07755_ (.A(_00809_),
    .B(_00811_),
    .Y(_00847_));
 sky130_fd_sc_hd__or2_1 _07756_ (.A(_00846_),
    .B(_00847_),
    .X(_00848_));
 sky130_fd_sc_hd__o21ai_1 _07757_ (.A1(_00846_),
    .A2(_00847_),
    .B1(_00845_),
    .Y(_00849_));
 sky130_fd_sc_hd__o22a_1 _07758_ (.A1(net147),
    .A2(net84),
    .B1(net80),
    .B2(net145),
    .X(_00850_));
 sky130_fd_sc_hd__xnor2_2 _07759_ (.A(net201),
    .B(_00850_),
    .Y(_00851_));
 sky130_fd_sc_hd__o22a_1 _07760_ (.A1(net119),
    .A2(net107),
    .B1(net105),
    .B2(net117),
    .X(_00852_));
 sky130_fd_sc_hd__xnor2_2 _07761_ (.A(net136),
    .B(_00852_),
    .Y(_00853_));
 sky130_fd_sc_hd__nor2_1 _07762_ (.A(_00851_),
    .B(_00853_),
    .Y(_00854_));
 sky130_fd_sc_hd__xor2_2 _07763_ (.A(_00851_),
    .B(_00853_),
    .X(_00855_));
 sky130_fd_sc_hd__o22a_1 _07764_ (.A1(net133),
    .A2(net76),
    .B1(net72),
    .B2(net131),
    .X(_00856_));
 sky130_fd_sc_hd__xnor2_2 _07765_ (.A(net180),
    .B(_00856_),
    .Y(_00857_));
 sky130_fd_sc_hd__inv_2 _07766_ (.A(_00857_),
    .Y(_00858_));
 sky130_fd_sc_hd__a21oi_2 _07767_ (.A1(_00855_),
    .A2(_00858_),
    .B1(_00854_),
    .Y(_00859_));
 sky130_fd_sc_hd__o22a_1 _07768_ (.A1(net216),
    .A2(net46),
    .B1(net144),
    .B2(net48),
    .X(_00860_));
 sky130_fd_sc_hd__xnor2_2 _07769_ (.A(net97),
    .B(_00860_),
    .Y(_00861_));
 sky130_fd_sc_hd__and2b_1 _07770_ (.A_N(_00859_),
    .B(_00861_),
    .X(_00862_));
 sky130_fd_sc_hd__o22a_1 _07771_ (.A1(net288),
    .A2(net63),
    .B1(net61),
    .B2(_06520_),
    .X(_00863_));
 sky130_fd_sc_hd__xnor2_1 _07772_ (.A(net238),
    .B(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__o22a_1 _07773_ (.A1(net155),
    .A2(net100),
    .B1(net98),
    .B2(net153),
    .X(_00865_));
 sky130_fd_sc_hd__xnor2_1 _07774_ (.A(net208),
    .B(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__nor2_1 _07775_ (.A(_00864_),
    .B(_00866_),
    .Y(_00867_));
 sky130_fd_sc_hd__nand2_1 _07776_ (.A(_00864_),
    .B(_00866_),
    .Y(_00868_));
 sky130_fd_sc_hd__xnor2_1 _07777_ (.A(_00864_),
    .B(_00866_),
    .Y(_00869_));
 sky130_fd_sc_hd__o22a_1 _07778_ (.A1(net152),
    .A2(net53),
    .B1(net51),
    .B2(net150),
    .X(_00870_));
 sky130_fd_sc_hd__xor2_1 _07779_ (.A(net204),
    .B(_00870_),
    .X(_00871_));
 sky130_fd_sc_hd__a21o_1 _07780_ (.A1(_00868_),
    .A2(_00871_),
    .B1(_00867_),
    .X(_00872_));
 sky130_fd_sc_hd__xnor2_2 _07781_ (.A(_00859_),
    .B(_00861_),
    .Y(_00873_));
 sky130_fd_sc_hd__a21oi_2 _07782_ (.A1(_00872_),
    .A2(_00873_),
    .B1(_00862_),
    .Y(_00874_));
 sky130_fd_sc_hd__a21o_1 _07783_ (.A1(_00845_),
    .A2(_00848_),
    .B1(_00874_),
    .X(_00875_));
 sky130_fd_sc_hd__xor2_1 _07784_ (.A(_00792_),
    .B(_00793_),
    .X(_00876_));
 sky130_fd_sc_hd__o22a_1 _07785_ (.A1(net111),
    .A2(net86),
    .B1(net82),
    .B2(net109),
    .X(_00877_));
 sky130_fd_sc_hd__xnor2_1 _07786_ (.A(net138),
    .B(_00877_),
    .Y(_00878_));
 sky130_fd_sc_hd__o22a_1 _07787_ (.A1(net130),
    .A2(net33),
    .B1(_00375_),
    .B2(net35),
    .X(_00879_));
 sky130_fd_sc_hd__xnor2_1 _07788_ (.A(net124),
    .B(_00879_),
    .Y(_00880_));
 sky130_fd_sc_hd__nor2_1 _07789_ (.A(_00878_),
    .B(_00880_),
    .Y(_00881_));
 sky130_fd_sc_hd__xnor2_1 _07790_ (.A(_00878_),
    .B(_00880_),
    .Y(_00882_));
 sky130_fd_sc_hd__o22a_1 _07791_ (.A1(_00309_),
    .A2(net79),
    .B1(net75),
    .B2(_00313_),
    .X(_00883_));
 sky130_fd_sc_hd__xnor2_1 _07792_ (.A(net121),
    .B(_00883_),
    .Y(_00884_));
 sky130_fd_sc_hd__o21ba_1 _07793_ (.A1(_00882_),
    .A2(_00884_),
    .B1_N(_00881_),
    .X(_00885_));
 sky130_fd_sc_hd__and2b_1 _07794_ (.A_N(_00885_),
    .B(_00876_),
    .X(_00886_));
 sky130_fd_sc_hd__o22a_1 _07795_ (.A1(net127),
    .A2(net27),
    .B1(net25),
    .B2(net141),
    .X(_00887_));
 sky130_fd_sc_hd__xnor2_2 _07796_ (.A(net88),
    .B(_00887_),
    .Y(_00888_));
 sky130_fd_sc_hd__a22o_1 _07797_ (.A1(_00265_),
    .A2(net31),
    .B1(net29),
    .B2(_00240_),
    .X(_00889_));
 sky130_fd_sc_hd__xnor2_2 _07798_ (.A(net49),
    .B(_00889_),
    .Y(_00890_));
 sky130_fd_sc_hd__and2_1 _07799_ (.A(_00888_),
    .B(_00890_),
    .X(_00891_));
 sky130_fd_sc_hd__xnor2_1 _07800_ (.A(_00876_),
    .B(_00885_),
    .Y(_00892_));
 sky130_fd_sc_hd__a21o_1 _07801_ (.A1(_00891_),
    .A2(_00892_),
    .B1(_00886_),
    .X(_00893_));
 sky130_fd_sc_hd__xnor2_2 _07802_ (.A(_00849_),
    .B(_00874_),
    .Y(_00894_));
 sky130_fd_sc_hd__a21bo_1 _07803_ (.A1(_00893_),
    .A2(_00894_),
    .B1_N(_00875_),
    .X(_00895_));
 sky130_fd_sc_hd__xnor2_1 _07804_ (.A(_00794_),
    .B(_00795_),
    .Y(_00896_));
 sky130_fd_sc_hd__xnor2_1 _07805_ (.A(_00800_),
    .B(_00801_),
    .Y(_00897_));
 sky130_fd_sc_hd__xnor2_1 _07806_ (.A(_00819_),
    .B(_00820_),
    .Y(_00898_));
 sky130_fd_sc_hd__xnor2_1 _07807_ (.A(_00896_),
    .B(_00897_),
    .Y(_00899_));
 sky130_fd_sc_hd__nor2_1 _07808_ (.A(_00898_),
    .B(_00899_),
    .Y(_00900_));
 sky130_fd_sc_hd__o21ba_1 _07809_ (.A1(_00896_),
    .A2(_00897_),
    .B1_N(_00900_),
    .X(_00901_));
 sky130_fd_sc_hd__xor2_1 _07810_ (.A(_00842_),
    .B(_00895_),
    .X(_00902_));
 sky130_fd_sc_hd__nand2b_1 _07811_ (.A_N(_00901_),
    .B(_00902_),
    .Y(_00903_));
 sky130_fd_sc_hd__a21bo_1 _07812_ (.A1(_00842_),
    .A2(_00895_),
    .B1_N(_00903_),
    .X(_00904_));
 sky130_fd_sc_hd__xnor2_1 _07813_ (.A(_00840_),
    .B(_00841_),
    .Y(_00905_));
 sky130_fd_sc_hd__nand2b_1 _07814_ (.A_N(_00905_),
    .B(_00904_),
    .Y(_00906_));
 sky130_fd_sc_hd__a21bo_2 _07815_ (.A1(_00840_),
    .A2(_00841_),
    .B1_N(_00906_),
    .X(_00907_));
 sky130_fd_sc_hd__xor2_4 _07816_ (.A(_00836_),
    .B(_00837_),
    .X(_00908_));
 sky130_fd_sc_hd__nand2_1 _07817_ (.A(_00907_),
    .B(_00908_),
    .Y(_00909_));
 sky130_fd_sc_hd__a2bb2o_1 _07818_ (.A1_N(_00769_),
    .A2_N(_00838_),
    .B1(_00907_),
    .B2(_00908_),
    .X(_00910_));
 sky130_fd_sc_hd__xnor2_1 _07819_ (.A(_00831_),
    .B(_00833_),
    .Y(_00911_));
 sky130_fd_sc_hd__xnor2_1 _07820_ (.A(_00901_),
    .B(_00902_),
    .Y(_00912_));
 sky130_fd_sc_hd__nand2_1 _07821_ (.A(_00911_),
    .B(_00912_),
    .Y(_00913_));
 sky130_fd_sc_hd__xnor2_2 _07822_ (.A(_00893_),
    .B(_00894_),
    .Y(_00914_));
 sky130_fd_sc_hd__xor2_2 _07823_ (.A(_00888_),
    .B(_00890_),
    .X(_00915_));
 sky130_fd_sc_hd__xnor2_2 _07824_ (.A(_00855_),
    .B(_00857_),
    .Y(_00916_));
 sky130_fd_sc_hd__nand2_1 _07825_ (.A(_00915_),
    .B(_00916_),
    .Y(_00917_));
 sky130_fd_sc_hd__xnor2_1 _07826_ (.A(_00882_),
    .B(_00884_),
    .Y(_00918_));
 sky130_fd_sc_hd__nor2_1 _07827_ (.A(_00915_),
    .B(_00916_),
    .Y(_00919_));
 sky130_fd_sc_hd__xor2_1 _07828_ (.A(_00915_),
    .B(_00916_),
    .X(_00920_));
 sky130_fd_sc_hd__o21a_2 _07829_ (.A1(_00918_),
    .A2(_00919_),
    .B1(_00917_),
    .X(_00921_));
 sky130_fd_sc_hd__nor2_1 _07830_ (.A(net216),
    .B(net48),
    .Y(_00922_));
 sky130_fd_sc_hd__a21oi_1 _07831_ (.A1(_06544_),
    .A2(_06545_),
    .B1(net288),
    .Y(_00923_));
 sky130_fd_sc_hd__and3_1 _07832_ (.A(_06519_),
    .B(_00161_),
    .C(_00162_),
    .X(_00924_));
 sky130_fd_sc_hd__o21a_1 _07833_ (.A1(_00923_),
    .A2(_00924_),
    .B1(net240),
    .X(_00925_));
 sky130_fd_sc_hd__nor3_1 _07834_ (.A(net240),
    .B(_00923_),
    .C(_00924_),
    .Y(_00926_));
 sky130_fd_sc_hd__o22a_1 _07835_ (.A1(net156),
    .A2(net98),
    .B1(net84),
    .B2(net154),
    .X(_00927_));
 sky130_fd_sc_hd__xnor2_1 _07836_ (.A(net207),
    .B(_00927_),
    .Y(_00928_));
 sky130_fd_sc_hd__or3_1 _07837_ (.A(_00925_),
    .B(_00926_),
    .C(_00928_),
    .X(_00929_));
 sky130_fd_sc_hd__o21ai_1 _07838_ (.A1(_00925_),
    .A2(_00926_),
    .B1(_00928_),
    .Y(_00930_));
 sky130_fd_sc_hd__o22a_1 _07839_ (.A1(net152),
    .A2(net51),
    .B1(net100),
    .B2(net150),
    .X(_00931_));
 sky130_fd_sc_hd__xor2_1 _07840_ (.A(net205),
    .B(_00931_),
    .X(_00932_));
 sky130_fd_sc_hd__nand3_1 _07841_ (.A(_00929_),
    .B(_00930_),
    .C(_00932_),
    .Y(_00933_));
 sky130_fd_sc_hd__nand2_1 _07842_ (.A(_00929_),
    .B(_00933_),
    .Y(_00934_));
 sky130_fd_sc_hd__mux2_2 _07843_ (.A0(net97),
    .A1(_00934_),
    .S(_00922_),
    .X(_00935_));
 sky130_fd_sc_hd__nand2b_1 _07844_ (.A_N(_00921_),
    .B(_00935_),
    .Y(_00936_));
 sky130_fd_sc_hd__xnor2_1 _07845_ (.A(_00869_),
    .B(_00871_),
    .Y(_00937_));
 sky130_fd_sc_hd__o22a_1 _07846_ (.A1(net117),
    .A2(net107),
    .B1(net105),
    .B2(net111),
    .X(_00938_));
 sky130_fd_sc_hd__xnor2_1 _07847_ (.A(net136),
    .B(_00938_),
    .Y(_00939_));
 sky130_fd_sc_hd__o22a_1 _07848_ (.A1(net148),
    .A2(net80),
    .B1(net76),
    .B2(net145),
    .X(_00940_));
 sky130_fd_sc_hd__xnor2_1 _07849_ (.A(net201),
    .B(_00940_),
    .Y(_00941_));
 sky130_fd_sc_hd__xor2_1 _07850_ (.A(_00939_),
    .B(_00941_),
    .X(_00942_));
 sky130_fd_sc_hd__o22a_1 _07851_ (.A1(net131),
    .A2(net119),
    .B1(net72),
    .B2(net133),
    .X(_00943_));
 sky130_fd_sc_hd__xnor2_1 _07852_ (.A(net182),
    .B(_00943_),
    .Y(_00944_));
 sky130_fd_sc_hd__and2b_1 _07853_ (.A_N(_00944_),
    .B(_00942_),
    .X(_00945_));
 sky130_fd_sc_hd__o21ba_1 _07854_ (.A1(_00939_),
    .A2(_00941_),
    .B1_N(_00945_),
    .X(_00946_));
 sky130_fd_sc_hd__and2b_1 _07855_ (.A_N(_00946_),
    .B(_00937_),
    .X(_00947_));
 sky130_fd_sc_hd__o22a_1 _07856_ (.A1(net109),
    .A2(net87),
    .B1(net83),
    .B2(net115),
    .X(_00948_));
 sky130_fd_sc_hd__xnor2_1 _07857_ (.A(net138),
    .B(_00948_),
    .Y(_00949_));
 sky130_fd_sc_hd__o22a_1 _07858_ (.A1(net114),
    .A2(net79),
    .B1(net75),
    .B2(net108),
    .X(_00950_));
 sky130_fd_sc_hd__xnor2_1 _07859_ (.A(net123),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__nor2_1 _07860_ (.A(_00949_),
    .B(_00951_),
    .Y(_00952_));
 sky130_fd_sc_hd__xnor2_1 _07861_ (.A(_00937_),
    .B(_00946_),
    .Y(_00953_));
 sky130_fd_sc_hd__a21o_2 _07862_ (.A1(_00952_),
    .A2(_00953_),
    .B1(_00947_),
    .X(_00954_));
 sky130_fd_sc_hd__xnor2_4 _07863_ (.A(_00921_),
    .B(_00935_),
    .Y(_00955_));
 sky130_fd_sc_hd__a21bo_1 _07864_ (.A1(_00954_),
    .A2(_00955_),
    .B1_N(_00936_),
    .X(_00956_));
 sky130_fd_sc_hd__and2b_1 _07865_ (.A_N(_00914_),
    .B(_00956_),
    .X(_00957_));
 sky130_fd_sc_hd__xor2_2 _07866_ (.A(_00846_),
    .B(_00847_),
    .X(_00958_));
 sky130_fd_sc_hd__xor2_2 _07867_ (.A(_00872_),
    .B(_00873_),
    .X(_00959_));
 sky130_fd_sc_hd__xnor2_1 _07868_ (.A(_00958_),
    .B(_00959_),
    .Y(_00960_));
 sky130_fd_sc_hd__xnor2_1 _07869_ (.A(_00891_),
    .B(_00892_),
    .Y(_00961_));
 sky130_fd_sc_hd__nor2_1 _07870_ (.A(_00960_),
    .B(_00961_),
    .Y(_00962_));
 sky130_fd_sc_hd__a21oi_2 _07871_ (.A1(_00958_),
    .A2(_00959_),
    .B1(_00962_),
    .Y(_00963_));
 sky130_fd_sc_hd__xnor2_2 _07872_ (.A(_00914_),
    .B(_00956_),
    .Y(_00964_));
 sky130_fd_sc_hd__and2b_1 _07873_ (.A_N(_00963_),
    .B(_00964_),
    .X(_00965_));
 sky130_fd_sc_hd__xor2_1 _07874_ (.A(_00911_),
    .B(_00912_),
    .X(_00966_));
 sky130_fd_sc_hd__o21ai_1 _07875_ (.A1(_00957_),
    .A2(_00965_),
    .B1(_00966_),
    .Y(_00967_));
 sky130_fd_sc_hd__xor2_1 _07876_ (.A(_00904_),
    .B(_00905_),
    .X(_00968_));
 sky130_fd_sc_hd__and3_1 _07877_ (.A(_00913_),
    .B(_00967_),
    .C(_00968_),
    .X(_00969_));
 sky130_fd_sc_hd__and2_1 _07878_ (.A(_00898_),
    .B(_00899_),
    .X(_00970_));
 sky130_fd_sc_hd__nor2_1 _07879_ (.A(_00900_),
    .B(_00970_),
    .Y(_00971_));
 sky130_fd_sc_hd__xnor2_2 _07880_ (.A(_00963_),
    .B(_00964_),
    .Y(_00972_));
 sky130_fd_sc_hd__nand2_1 _07881_ (.A(_00971_),
    .B(_00972_),
    .Y(_00973_));
 sky130_fd_sc_hd__a21o_1 _07882_ (.A1(_00929_),
    .A2(_00930_),
    .B1(_00932_),
    .X(_00974_));
 sky130_fd_sc_hd__and2_1 _07883_ (.A(_00949_),
    .B(_00951_),
    .X(_00975_));
 sky130_fd_sc_hd__nor2_1 _07884_ (.A(_00952_),
    .B(_00975_),
    .Y(_00976_));
 sky130_fd_sc_hd__and3_1 _07885_ (.A(_00933_),
    .B(_00974_),
    .C(_00976_),
    .X(_00977_));
 sky130_fd_sc_hd__a21oi_1 _07886_ (.A1(_00933_),
    .A2(_00974_),
    .B1(_00976_),
    .Y(_00978_));
 sky130_fd_sc_hd__and2b_1 _07887_ (.A_N(_00942_),
    .B(_00944_),
    .X(_00979_));
 sky130_fd_sc_hd__or2_1 _07888_ (.A(_00945_),
    .B(_00979_),
    .X(_00980_));
 sky130_fd_sc_hd__or3_1 _07889_ (.A(_00977_),
    .B(_00978_),
    .C(_00980_),
    .X(_00981_));
 sky130_fd_sc_hd__o21ba_1 _07890_ (.A1(_00978_),
    .A2(_00980_),
    .B1_N(_00977_),
    .X(_00982_));
 sky130_fd_sc_hd__o22a_1 _07891_ (.A1(net130),
    .A2(net35),
    .B1(net33),
    .B2(net128),
    .X(_00983_));
 sky130_fd_sc_hd__xnor2_1 _07892_ (.A(net125),
    .B(_00983_),
    .Y(_00984_));
 sky130_fd_sc_hd__a22o_1 _07893_ (.A1(_00240_),
    .A2(net31),
    .B1(net29),
    .B2(net214),
    .X(_00985_));
 sky130_fd_sc_hd__xnor2_1 _07894_ (.A(net49),
    .B(_00985_),
    .Y(_00986_));
 sky130_fd_sc_hd__and2_1 _07895_ (.A(_00984_),
    .B(_00986_),
    .X(_00987_));
 sky130_fd_sc_hd__nor2_1 _07896_ (.A(_00984_),
    .B(_00986_),
    .Y(_00988_));
 sky130_fd_sc_hd__nor2_1 _07897_ (.A(_00987_),
    .B(_00988_),
    .Y(_00989_));
 sky130_fd_sc_hd__o22a_1 _07898_ (.A1(net142),
    .A2(net27),
    .B1(net25),
    .B2(_00264_),
    .X(_00990_));
 sky130_fd_sc_hd__xnor2_2 _07899_ (.A(net88),
    .B(_00990_),
    .Y(_00991_));
 sky130_fd_sc_hd__a21oi_2 _07900_ (.A1(_00989_),
    .A2(_00991_),
    .B1(_00987_),
    .Y(_00992_));
 sky130_fd_sc_hd__nor2_1 _07901_ (.A(_00982_),
    .B(_00992_),
    .Y(_00993_));
 sky130_fd_sc_hd__o22a_1 _07902_ (.A1(net115),
    .A2(net87),
    .B1(net83),
    .B2(net114),
    .X(_00994_));
 sky130_fd_sc_hd__xnor2_2 _07903_ (.A(net138),
    .B(_00994_),
    .Y(_00995_));
 sky130_fd_sc_hd__o22a_1 _07904_ (.A1(net129),
    .A2(net75),
    .B1(net108),
    .B2(net79),
    .X(_00996_));
 sky130_fd_sc_hd__xnor2_2 _07905_ (.A(net123),
    .B(_00996_),
    .Y(_00997_));
 sky130_fd_sc_hd__nor2_1 _07906_ (.A(_00995_),
    .B(_00997_),
    .Y(_00998_));
 sky130_fd_sc_hd__and3_1 _07907_ (.A(net292),
    .B(_00161_),
    .C(_00162_),
    .X(_00999_));
 sky130_fd_sc_hd__a21oi_1 _07908_ (.A1(_00169_),
    .A2(_00170_),
    .B1(net237),
    .Y(_01000_));
 sky130_fd_sc_hd__o21ai_1 _07909_ (.A1(_00999_),
    .A2(_01000_),
    .B1(net240),
    .Y(_01001_));
 sky130_fd_sc_hd__or3_1 _07910_ (.A(net240),
    .B(_00999_),
    .C(_01000_),
    .X(_01002_));
 sky130_fd_sc_hd__o22a_1 _07911_ (.A1(net156),
    .A2(net84),
    .B1(net80),
    .B2(net154),
    .X(_01003_));
 sky130_fd_sc_hd__xnor2_1 _07912_ (.A(_06532_),
    .B(_01003_),
    .Y(_01004_));
 sky130_fd_sc_hd__and3_1 _07913_ (.A(_01001_),
    .B(_01002_),
    .C(_01004_),
    .X(_01005_));
 sky130_fd_sc_hd__a22o_1 _07914_ (.A1(_06557_),
    .A2(_00179_),
    .B1(_00189_),
    .B2(_06565_),
    .X(_01006_));
 sky130_fd_sc_hd__xnor2_1 _07915_ (.A(net205),
    .B(_01006_),
    .Y(_01007_));
 sky130_fd_sc_hd__a21oi_1 _07916_ (.A1(_01001_),
    .A2(_01002_),
    .B1(_01004_),
    .Y(_01008_));
 sky130_fd_sc_hd__a21o_1 _07917_ (.A1(_01001_),
    .A2(_01002_),
    .B1(_01004_),
    .X(_01009_));
 sky130_fd_sc_hd__or3b_1 _07918_ (.A(_01005_),
    .B(_01008_),
    .C_N(_01007_),
    .X(_01010_));
 sky130_fd_sc_hd__a21oi_2 _07919_ (.A1(_01007_),
    .A2(_01009_),
    .B1(_01005_),
    .Y(_01011_));
 sky130_fd_sc_hd__o22a_1 _07920_ (.A1(net147),
    .A2(net76),
    .B1(net72),
    .B2(net145),
    .X(_01012_));
 sky130_fd_sc_hd__xnor2_1 _07921_ (.A(net203),
    .B(_01012_),
    .Y(_01013_));
 sky130_fd_sc_hd__o22a_1 _07922_ (.A1(net111),
    .A2(net107),
    .B1(net105),
    .B2(net109),
    .X(_01014_));
 sky130_fd_sc_hd__xnor2_1 _07923_ (.A(net136),
    .B(_01014_),
    .Y(_01015_));
 sky130_fd_sc_hd__xor2_1 _07924_ (.A(_01013_),
    .B(_01015_),
    .X(_01016_));
 sky130_fd_sc_hd__o22a_1 _07925_ (.A1(net133),
    .A2(net119),
    .B1(net117),
    .B2(net131),
    .X(_01017_));
 sky130_fd_sc_hd__xnor2_1 _07926_ (.A(net182),
    .B(_01017_),
    .Y(_01018_));
 sky130_fd_sc_hd__and2b_1 _07927_ (.A_N(_01018_),
    .B(_01016_),
    .X(_01019_));
 sky130_fd_sc_hd__o21bai_2 _07928_ (.A1(_01013_),
    .A2(_01015_),
    .B1_N(_01019_),
    .Y(_01020_));
 sky130_fd_sc_hd__xnor2_1 _07929_ (.A(_00998_),
    .B(_01011_),
    .Y(_01021_));
 sky130_fd_sc_hd__nand2_1 _07930_ (.A(_01020_),
    .B(_01021_),
    .Y(_01022_));
 sky130_fd_sc_hd__o31ai_4 _07931_ (.A1(_00995_),
    .A2(_00997_),
    .A3(_01011_),
    .B1(_01022_),
    .Y(_01023_));
 sky130_fd_sc_hd__xor2_2 _07932_ (.A(_00982_),
    .B(_00992_),
    .X(_01024_));
 sky130_fd_sc_hd__a21o_2 _07933_ (.A1(_01023_),
    .A2(_01024_),
    .B1(_00993_),
    .X(_01025_));
 sky130_fd_sc_hd__xor2_4 _07934_ (.A(_00954_),
    .B(_00955_),
    .X(_01026_));
 sky130_fd_sc_hd__xnor2_1 _07935_ (.A(_00918_),
    .B(_00920_),
    .Y(_01027_));
 sky130_fd_sc_hd__xor2_1 _07936_ (.A(_00922_),
    .B(_00934_),
    .X(_01028_));
 sky130_fd_sc_hd__xnor2_1 _07937_ (.A(_00952_),
    .B(_00953_),
    .Y(_01029_));
 sky130_fd_sc_hd__xnor2_1 _07938_ (.A(_01027_),
    .B(_01028_),
    .Y(_01030_));
 sky130_fd_sc_hd__or2_1 _07939_ (.A(_01029_),
    .B(_01030_),
    .X(_01031_));
 sky130_fd_sc_hd__a21bo_2 _07940_ (.A1(_01027_),
    .A2(_01028_),
    .B1_N(_01031_),
    .X(_01032_));
 sky130_fd_sc_hd__xnor2_4 _07941_ (.A(_01025_),
    .B(_01026_),
    .Y(_01033_));
 sky130_fd_sc_hd__and2b_1 _07942_ (.A_N(_01033_),
    .B(_01032_),
    .X(_01034_));
 sky130_fd_sc_hd__a21o_2 _07943_ (.A1(_01025_),
    .A2(_01026_),
    .B1(_01034_),
    .X(_01035_));
 sky130_fd_sc_hd__xnor2_2 _07944_ (.A(_00971_),
    .B(_00972_),
    .Y(_01036_));
 sky130_fd_sc_hd__nand2b_1 _07945_ (.A_N(_01036_),
    .B(_01035_),
    .Y(_01037_));
 sky130_fd_sc_hd__or3_1 _07946_ (.A(_00957_),
    .B(_00965_),
    .C(_00966_),
    .X(_01038_));
 sky130_fd_sc_hd__nand2_1 _07947_ (.A(_00967_),
    .B(_01038_),
    .Y(_01039_));
 sky130_fd_sc_hd__and3_1 _07948_ (.A(_00973_),
    .B(_01037_),
    .C(_01039_),
    .X(_01040_));
 sky130_fd_sc_hd__a21o_1 _07949_ (.A1(_00973_),
    .A2(_01037_),
    .B1(_01039_),
    .X(_01041_));
 sky130_fd_sc_hd__nand2b_2 _07950_ (.A_N(_01040_),
    .B(_01041_),
    .Y(_01042_));
 sky130_fd_sc_hd__and2_1 _07951_ (.A(_00960_),
    .B(_00961_),
    .X(_01043_));
 sky130_fd_sc_hd__nor2_2 _07952_ (.A(_00962_),
    .B(_01043_),
    .Y(_01044_));
 sky130_fd_sc_hd__xnor2_4 _07953_ (.A(_01032_),
    .B(_01033_),
    .Y(_01045_));
 sky130_fd_sc_hd__nand2_1 _07954_ (.A(_01044_),
    .B(_01045_),
    .Y(_01046_));
 sky130_fd_sc_hd__xnor2_4 _07955_ (.A(_01044_),
    .B(_01045_),
    .Y(_01047_));
 sky130_fd_sc_hd__xnor2_2 _07956_ (.A(_01023_),
    .B(_01024_),
    .Y(_01048_));
 sky130_fd_sc_hd__o22a_1 _07957_ (.A1(net127),
    .A2(net35),
    .B1(net33),
    .B2(net141),
    .X(_01049_));
 sky130_fd_sc_hd__xnor2_1 _07958_ (.A(net125),
    .B(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__nand2_1 _07959_ (.A(net214),
    .B(net31),
    .Y(_01051_));
 sky130_fd_sc_hd__xnor2_2 _07960_ (.A(net49),
    .B(_01051_),
    .Y(_01052_));
 sky130_fd_sc_hd__and2b_1 _07961_ (.A_N(_01052_),
    .B(_01050_),
    .X(_01053_));
 sky130_fd_sc_hd__xor2_1 _07962_ (.A(_01050_),
    .B(_01052_),
    .X(_01054_));
 sky130_fd_sc_hd__o22a_1 _07963_ (.A1(net140),
    .A2(net27),
    .B1(net25),
    .B2(net143),
    .X(_01055_));
 sky130_fd_sc_hd__xnor2_1 _07964_ (.A(net88),
    .B(_01055_),
    .Y(_01056_));
 sky130_fd_sc_hd__and2b_1 _07965_ (.A_N(_01054_),
    .B(_01056_),
    .X(_01057_));
 sky130_fd_sc_hd__or2_1 _07966_ (.A(_01053_),
    .B(_01057_),
    .X(_01058_));
 sky130_fd_sc_hd__o21bai_1 _07967_ (.A1(_01005_),
    .A2(_01008_),
    .B1_N(_01007_),
    .Y(_01059_));
 sky130_fd_sc_hd__and2_1 _07968_ (.A(_00995_),
    .B(_00997_),
    .X(_01060_));
 sky130_fd_sc_hd__nor2_1 _07969_ (.A(_00998_),
    .B(_01060_),
    .Y(_01061_));
 sky130_fd_sc_hd__and3_1 _07970_ (.A(_01010_),
    .B(_01059_),
    .C(_01061_),
    .X(_01062_));
 sky130_fd_sc_hd__and2b_1 _07971_ (.A_N(_01016_),
    .B(_01018_),
    .X(_01063_));
 sky130_fd_sc_hd__or2_1 _07972_ (.A(_01019_),
    .B(_01063_),
    .X(_01064_));
 sky130_fd_sc_hd__a21oi_2 _07973_ (.A1(_01010_),
    .A2(_01059_),
    .B1(_01061_),
    .Y(_01065_));
 sky130_fd_sc_hd__or3_1 _07974_ (.A(_01062_),
    .B(_01064_),
    .C(_01065_),
    .X(_01066_));
 sky130_fd_sc_hd__o21ba_1 _07975_ (.A1(_01064_),
    .A2(_01065_),
    .B1_N(_01062_),
    .X(_01067_));
 sky130_fd_sc_hd__o21ba_1 _07976_ (.A1(_01053_),
    .A2(_01057_),
    .B1_N(_01067_),
    .X(_01068_));
 sky130_fd_sc_hd__o22a_1 _07977_ (.A1(net145),
    .A2(net119),
    .B1(net72),
    .B2(net147),
    .X(_01069_));
 sky130_fd_sc_hd__xnor2_1 _07978_ (.A(net201),
    .B(_01069_),
    .Y(_01070_));
 sky130_fd_sc_hd__o22a_1 _07979_ (.A1(net133),
    .A2(net117),
    .B1(net111),
    .B2(net131),
    .X(_01071_));
 sky130_fd_sc_hd__xnor2_1 _07980_ (.A(net180),
    .B(_01071_),
    .Y(_01072_));
 sky130_fd_sc_hd__or2_1 _07981_ (.A(_01070_),
    .B(_01072_),
    .X(_01073_));
 sky130_fd_sc_hd__a21o_1 _07982_ (.A1(_00169_),
    .A2(_00170_),
    .B1(net288),
    .X(_01074_));
 sky130_fd_sc_hd__nand2_1 _07983_ (.A(_06519_),
    .B(_00179_),
    .Y(_01075_));
 sky130_fd_sc_hd__a21oi_1 _07984_ (.A1(_01074_),
    .A2(_01075_),
    .B1(net238),
    .Y(_01076_));
 sky130_fd_sc_hd__and3_1 _07985_ (.A(net238),
    .B(_01074_),
    .C(_01075_),
    .X(_01077_));
 sky130_fd_sc_hd__o22a_1 _07986_ (.A1(net155),
    .A2(net80),
    .B1(net76),
    .B2(net153),
    .X(_01078_));
 sky130_fd_sc_hd__xnor2_1 _07987_ (.A(net208),
    .B(_01078_),
    .Y(_01079_));
 sky130_fd_sc_hd__or3_2 _07988_ (.A(_01076_),
    .B(_01077_),
    .C(_01079_),
    .X(_01080_));
 sky130_fd_sc_hd__a22o_1 _07989_ (.A1(_06557_),
    .A2(_00189_),
    .B1(_00348_),
    .B2(_06565_),
    .X(_01081_));
 sky130_fd_sc_hd__xnor2_1 _07990_ (.A(net204),
    .B(_01081_),
    .Y(_01082_));
 sky130_fd_sc_hd__o21ai_1 _07991_ (.A1(_01076_),
    .A2(_01077_),
    .B1(_01079_),
    .Y(_01083_));
 sky130_fd_sc_hd__nand3_2 _07992_ (.A(_01080_),
    .B(_01082_),
    .C(_01083_),
    .Y(_01084_));
 sky130_fd_sc_hd__xnor2_1 _07993_ (.A(net49),
    .B(_01073_),
    .Y(_01085_));
 sky130_fd_sc_hd__a21o_1 _07994_ (.A1(_01080_),
    .A2(_01084_),
    .B1(_01085_),
    .X(_01086_));
 sky130_fd_sc_hd__o21ai_2 _07995_ (.A1(net49),
    .A2(_01073_),
    .B1(_01086_),
    .Y(_01087_));
 sky130_fd_sc_hd__xnor2_2 _07996_ (.A(_01058_),
    .B(_01067_),
    .Y(_01088_));
 sky130_fd_sc_hd__a21o_1 _07997_ (.A1(_01087_),
    .A2(_01088_),
    .B1(_01068_),
    .X(_01089_));
 sky130_fd_sc_hd__nand2b_1 _07998_ (.A_N(_01048_),
    .B(_01089_),
    .Y(_01090_));
 sky130_fd_sc_hd__o21ai_1 _07999_ (.A1(_00977_),
    .A2(_00978_),
    .B1(_00980_),
    .Y(_01091_));
 sky130_fd_sc_hd__xor2_1 _08000_ (.A(_00989_),
    .B(_00991_),
    .X(_01092_));
 sky130_fd_sc_hd__and3_1 _08001_ (.A(_00981_),
    .B(_01091_),
    .C(_01092_),
    .X(_01093_));
 sky130_fd_sc_hd__a21oi_1 _08002_ (.A1(_00981_),
    .A2(_01091_),
    .B1(_01092_),
    .Y(_01094_));
 sky130_fd_sc_hd__xnor2_1 _08003_ (.A(_01020_),
    .B(_01021_),
    .Y(_01095_));
 sky130_fd_sc_hd__nor3_1 _08004_ (.A(_01093_),
    .B(_01094_),
    .C(_01095_),
    .Y(_01096_));
 sky130_fd_sc_hd__nor2_1 _08005_ (.A(_01093_),
    .B(_01096_),
    .Y(_01097_));
 sky130_fd_sc_hd__xnor2_2 _08006_ (.A(_01048_),
    .B(_01089_),
    .Y(_01098_));
 sky130_fd_sc_hd__nand2b_1 _08007_ (.A_N(_01097_),
    .B(_01098_),
    .Y(_01099_));
 sky130_fd_sc_hd__and2_1 _08008_ (.A(_01090_),
    .B(_01099_),
    .X(_01100_));
 sky130_fd_sc_hd__nand2_2 _08009_ (.A(_01090_),
    .B(_01099_),
    .Y(_01101_));
 sky130_fd_sc_hd__o21ai_4 _08010_ (.A1(_01047_),
    .A2(_01100_),
    .B1(_01046_),
    .Y(_01102_));
 sky130_fd_sc_hd__xnor2_4 _08011_ (.A(_01035_),
    .B(_01036_),
    .Y(_01103_));
 sky130_fd_sc_hd__nand2_1 _08012_ (.A(_01102_),
    .B(_01103_),
    .Y(_01104_));
 sky130_fd_sc_hd__xnor2_4 _08013_ (.A(_01102_),
    .B(_01103_),
    .Y(_01105_));
 sky130_fd_sc_hd__nand2_1 _08014_ (.A(_01029_),
    .B(_01030_),
    .Y(_01106_));
 sky130_fd_sc_hd__and2_1 _08015_ (.A(_01031_),
    .B(_01106_),
    .X(_01107_));
 sky130_fd_sc_hd__xnor2_2 _08016_ (.A(_01097_),
    .B(_01098_),
    .Y(_01108_));
 sky130_fd_sc_hd__and2_1 _08017_ (.A(_01107_),
    .B(_01108_),
    .X(_01109_));
 sky130_fd_sc_hd__o22a_1 _08018_ (.A1(net147),
    .A2(net119),
    .B1(net117),
    .B2(net145),
    .X(_01110_));
 sky130_fd_sc_hd__xnor2_1 _08019_ (.A(net201),
    .B(_01110_),
    .Y(_01111_));
 sky130_fd_sc_hd__o22a_1 _08020_ (.A1(net133),
    .A2(net111),
    .B1(net109),
    .B2(net131),
    .X(_01112_));
 sky130_fd_sc_hd__xnor2_1 _08021_ (.A(net180),
    .B(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__or2_1 _08022_ (.A(_01111_),
    .B(_01113_),
    .X(_01114_));
 sky130_fd_sc_hd__xnor2_1 _08023_ (.A(_01070_),
    .B(_01072_),
    .Y(_01115_));
 sky130_fd_sc_hd__nor2_1 _08024_ (.A(_01114_),
    .B(_01115_),
    .Y(_01116_));
 sky130_fd_sc_hd__xor2_1 _08025_ (.A(_01114_),
    .B(_01115_),
    .X(_01117_));
 sky130_fd_sc_hd__a21o_1 _08026_ (.A1(_01080_),
    .A2(_01083_),
    .B1(_01082_),
    .X(_01118_));
 sky130_fd_sc_hd__nand3_1 _08027_ (.A(_01084_),
    .B(_01117_),
    .C(_01118_),
    .Y(_01119_));
 sky130_fd_sc_hd__and2b_1 _08028_ (.A_N(_01116_),
    .B(_01119_),
    .X(_01120_));
 sky130_fd_sc_hd__a31o_1 _08029_ (.A1(_01084_),
    .A2(_01117_),
    .A3(_01118_),
    .B1(_01116_),
    .X(_01121_));
 sky130_fd_sc_hd__o22a_1 _08030_ (.A1(net109),
    .A2(net107),
    .B1(net105),
    .B2(net115),
    .X(_01122_));
 sky130_fd_sc_hd__xnor2_1 _08031_ (.A(net136),
    .B(_01122_),
    .Y(_01123_));
 sky130_fd_sc_hd__o22a_1 _08032_ (.A1(net129),
    .A2(net79),
    .B1(net75),
    .B2(net127),
    .X(_01124_));
 sky130_fd_sc_hd__xnor2_1 _08033_ (.A(net123),
    .B(_01124_),
    .Y(_01125_));
 sky130_fd_sc_hd__o22a_1 _08034_ (.A1(net114),
    .A2(net87),
    .B1(net83),
    .B2(net108),
    .X(_01126_));
 sky130_fd_sc_hd__xnor2_1 _08035_ (.A(net138),
    .B(_01126_),
    .Y(_01127_));
 sky130_fd_sc_hd__xnor2_1 _08036_ (.A(_01123_),
    .B(_01125_),
    .Y(_01128_));
 sky130_fd_sc_hd__or2_1 _08037_ (.A(_01127_),
    .B(_01128_),
    .X(_01129_));
 sky130_fd_sc_hd__o21a_1 _08038_ (.A1(_01123_),
    .A2(_01125_),
    .B1(_01129_),
    .X(_01130_));
 sky130_fd_sc_hd__o22a_1 _08039_ (.A1(net287),
    .A2(net100),
    .B1(net98),
    .B2(net237),
    .X(_01131_));
 sky130_fd_sc_hd__xnor2_2 _08040_ (.A(net238),
    .B(_01131_),
    .Y(_01132_));
 sky130_fd_sc_hd__o22a_1 _08041_ (.A1(net155),
    .A2(net76),
    .B1(net72),
    .B2(net153),
    .X(_01133_));
 sky130_fd_sc_hd__xnor2_2 _08042_ (.A(net208),
    .B(_01133_),
    .Y(_01134_));
 sky130_fd_sc_hd__or2_1 _08043_ (.A(_01132_),
    .B(_01134_),
    .X(_01135_));
 sky130_fd_sc_hd__o22a_1 _08044_ (.A1(net151),
    .A2(net84),
    .B1(net80),
    .B2(net149),
    .X(_01136_));
 sky130_fd_sc_hd__xnor2_2 _08045_ (.A(net204),
    .B(_01136_),
    .Y(_01137_));
 sky130_fd_sc_hd__xnor2_2 _08046_ (.A(_01132_),
    .B(_01134_),
    .Y(_01138_));
 sky130_fd_sc_hd__o21ai_2 _08047_ (.A1(_01137_),
    .A2(_01138_),
    .B1(_01135_),
    .Y(_01139_));
 sky130_fd_sc_hd__o22a_1 _08048_ (.A1(net141),
    .A2(net35),
    .B1(net33),
    .B2(net140),
    .X(_01140_));
 sky130_fd_sc_hd__xnor2_1 _08049_ (.A(net125),
    .B(_01140_),
    .Y(_01141_));
 sky130_fd_sc_hd__nand2_1 _08050_ (.A(_01139_),
    .B(_01141_),
    .Y(_01142_));
 sky130_fd_sc_hd__xnor2_1 _08051_ (.A(_01139_),
    .B(_01141_),
    .Y(_01143_));
 sky130_fd_sc_hd__o22a_1 _08052_ (.A1(net143),
    .A2(net27),
    .B1(net25),
    .B2(net215),
    .X(_01144_));
 sky130_fd_sc_hd__xnor2_1 _08053_ (.A(net88),
    .B(_01144_),
    .Y(_01145_));
 sky130_fd_sc_hd__inv_2 _08054_ (.A(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hd__o21a_1 _08055_ (.A1(_01143_),
    .A2(_01146_),
    .B1(_01142_),
    .X(_01147_));
 sky130_fd_sc_hd__xnor2_2 _08056_ (.A(_01121_),
    .B(_01130_),
    .Y(_01148_));
 sky130_fd_sc_hd__nand2b_1 _08057_ (.A_N(_01147_),
    .B(_01148_),
    .Y(_01149_));
 sky130_fd_sc_hd__o21ai_2 _08058_ (.A1(_01120_),
    .A2(_01130_),
    .B1(_01149_),
    .Y(_01150_));
 sky130_fd_sc_hd__xnor2_2 _08059_ (.A(_01087_),
    .B(_01088_),
    .Y(_01151_));
 sky130_fd_sc_hd__nand2b_1 _08060_ (.A_N(_01151_),
    .B(_01150_),
    .Y(_01152_));
 sky130_fd_sc_hd__and2b_1 _08061_ (.A_N(_01056_),
    .B(_01054_),
    .X(_01153_));
 sky130_fd_sc_hd__nor2_1 _08062_ (.A(_01057_),
    .B(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__o21ai_1 _08063_ (.A1(_01062_),
    .A2(_01065_),
    .B1(_01064_),
    .Y(_01155_));
 sky130_fd_sc_hd__and3_1 _08064_ (.A(_01066_),
    .B(_01154_),
    .C(_01155_),
    .X(_01156_));
 sky130_fd_sc_hd__nand3_1 _08065_ (.A(_01080_),
    .B(_01084_),
    .C(_01085_),
    .Y(_01157_));
 sky130_fd_sc_hd__nand2_1 _08066_ (.A(_01086_),
    .B(_01157_),
    .Y(_01158_));
 sky130_fd_sc_hd__a21oi_1 _08067_ (.A1(_01066_),
    .A2(_01155_),
    .B1(_01154_),
    .Y(_01159_));
 sky130_fd_sc_hd__or3_1 _08068_ (.A(_01156_),
    .B(_01158_),
    .C(_01159_),
    .X(_01160_));
 sky130_fd_sc_hd__and2b_1 _08069_ (.A_N(_01156_),
    .B(_01160_),
    .X(_01161_));
 sky130_fd_sc_hd__xnor2_2 _08070_ (.A(_01150_),
    .B(_01151_),
    .Y(_01162_));
 sky130_fd_sc_hd__nand2b_1 _08071_ (.A_N(_01161_),
    .B(_01162_),
    .Y(_01163_));
 sky130_fd_sc_hd__nand2_1 _08072_ (.A(_01152_),
    .B(_01163_),
    .Y(_01164_));
 sky130_fd_sc_hd__xor2_2 _08073_ (.A(_01107_),
    .B(_01108_),
    .X(_01165_));
 sky130_fd_sc_hd__a21o_1 _08074_ (.A1(_01164_),
    .A2(_01165_),
    .B1(_01109_),
    .X(_01166_));
 sky130_fd_sc_hd__xnor2_4 _08075_ (.A(_01047_),
    .B(_01101_),
    .Y(_01167_));
 sky130_fd_sc_hd__xnor2_2 _08076_ (.A(_01166_),
    .B(_01167_),
    .Y(_01168_));
 sky130_fd_sc_hd__or2_1 _08077_ (.A(_01105_),
    .B(_01168_),
    .X(_01169_));
 sky130_fd_sc_hd__o21ai_1 _08078_ (.A1(_01156_),
    .A2(_01159_),
    .B1(_01158_),
    .Y(_01170_));
 sky130_fd_sc_hd__nand2_2 _08079_ (.A(_01160_),
    .B(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hd__a21o_1 _08080_ (.A1(_01084_),
    .A2(_01118_),
    .B1(_01117_),
    .X(_01172_));
 sky130_fd_sc_hd__nand2_1 _08081_ (.A(_01127_),
    .B(_01128_),
    .Y(_01173_));
 sky130_fd_sc_hd__and2_1 _08082_ (.A(_01129_),
    .B(_01173_),
    .X(_01174_));
 sky130_fd_sc_hd__and3_1 _08083_ (.A(_01119_),
    .B(_01172_),
    .C(_01174_),
    .X(_01175_));
 sky130_fd_sc_hd__a21oi_1 _08084_ (.A1(_01119_),
    .A2(_01172_),
    .B1(_01174_),
    .Y(_01176_));
 sky130_fd_sc_hd__xnor2_1 _08085_ (.A(_01143_),
    .B(_01146_),
    .Y(_01177_));
 sky130_fd_sc_hd__nor3_1 _08086_ (.A(_01175_),
    .B(_01176_),
    .C(_01177_),
    .Y(_01178_));
 sky130_fd_sc_hd__or2_1 _08087_ (.A(_01175_),
    .B(_01178_),
    .X(_01179_));
 sky130_fd_sc_hd__xnor2_2 _08088_ (.A(_01147_),
    .B(_01148_),
    .Y(_01180_));
 sky130_fd_sc_hd__o22a_1 _08089_ (.A1(net287),
    .A2(net98),
    .B1(net84),
    .B2(net237),
    .X(_01181_));
 sky130_fd_sc_hd__xnor2_1 _08090_ (.A(net238),
    .B(_01181_),
    .Y(_01182_));
 sky130_fd_sc_hd__o22a_1 _08091_ (.A1(net151),
    .A2(net80),
    .B1(net76),
    .B2(net149),
    .X(_01183_));
 sky130_fd_sc_hd__xnor2_1 _08092_ (.A(net204),
    .B(_01183_),
    .Y(_01184_));
 sky130_fd_sc_hd__or2_1 _08093_ (.A(_01182_),
    .B(_01184_),
    .X(_01185_));
 sky130_fd_sc_hd__nand2_1 _08094_ (.A(_01111_),
    .B(_01113_),
    .Y(_01186_));
 sky130_fd_sc_hd__nand2_1 _08095_ (.A(_01114_),
    .B(_01186_),
    .Y(_01187_));
 sky130_fd_sc_hd__nor2_1 _08096_ (.A(_01185_),
    .B(_01187_),
    .Y(_01188_));
 sky130_fd_sc_hd__nand2_1 _08097_ (.A(_01185_),
    .B(_01187_),
    .Y(_01189_));
 sky130_fd_sc_hd__xnor2_1 _08098_ (.A(_01185_),
    .B(_01187_),
    .Y(_01190_));
 sky130_fd_sc_hd__xor2_2 _08099_ (.A(_01137_),
    .B(_01138_),
    .X(_01191_));
 sky130_fd_sc_hd__a21o_1 _08100_ (.A1(_01189_),
    .A2(_01191_),
    .B1(_01188_),
    .X(_01192_));
 sky130_fd_sc_hd__o22a_1 _08101_ (.A1(net115),
    .A2(net107),
    .B1(net105),
    .B2(net114),
    .X(_01193_));
 sky130_fd_sc_hd__xnor2_1 _08102_ (.A(net136),
    .B(_01193_),
    .Y(_01194_));
 sky130_fd_sc_hd__o22a_1 _08103_ (.A1(net127),
    .A2(net79),
    .B1(net75),
    .B2(net141),
    .X(_01195_));
 sky130_fd_sc_hd__xnor2_1 _08104_ (.A(net123),
    .B(_01195_),
    .Y(_01196_));
 sky130_fd_sc_hd__nor2_1 _08105_ (.A(_01194_),
    .B(_01196_),
    .Y(_01197_));
 sky130_fd_sc_hd__o22a_1 _08106_ (.A1(net129),
    .A2(net83),
    .B1(net108),
    .B2(net87),
    .X(_01198_));
 sky130_fd_sc_hd__xnor2_1 _08107_ (.A(net138),
    .B(_01198_),
    .Y(_01199_));
 sky130_fd_sc_hd__xnor2_1 _08108_ (.A(_01194_),
    .B(_01196_),
    .Y(_01200_));
 sky130_fd_sc_hd__nor2_1 _08109_ (.A(_01199_),
    .B(_01200_),
    .Y(_01201_));
 sky130_fd_sc_hd__nor2_1 _08110_ (.A(_01197_),
    .B(_01201_),
    .Y(_01202_));
 sky130_fd_sc_hd__o21a_1 _08111_ (.A1(_01197_),
    .A2(_01201_),
    .B1(_01192_),
    .X(_01203_));
 sky130_fd_sc_hd__nor2_1 _08112_ (.A(net215),
    .B(net27),
    .Y(_01204_));
 sky130_fd_sc_hd__o22a_1 _08113_ (.A1(net140),
    .A2(net35),
    .B1(net33),
    .B2(net143),
    .X(_01205_));
 sky130_fd_sc_hd__xnor2_1 _08114_ (.A(net125),
    .B(_01205_),
    .Y(_01206_));
 sky130_fd_sc_hd__mux2_2 _08115_ (.A0(net88),
    .A1(_01206_),
    .S(_01204_),
    .X(_01207_));
 sky130_fd_sc_hd__xnor2_2 _08116_ (.A(_01192_),
    .B(_01202_),
    .Y(_01208_));
 sky130_fd_sc_hd__a21oi_2 _08117_ (.A1(_01207_),
    .A2(_01208_),
    .B1(_01203_),
    .Y(_01209_));
 sky130_fd_sc_hd__and2b_1 _08118_ (.A_N(_01209_),
    .B(_01180_),
    .X(_01210_));
 sky130_fd_sc_hd__xnor2_2 _08119_ (.A(_01180_),
    .B(_01209_),
    .Y(_01211_));
 sky130_fd_sc_hd__xnor2_2 _08120_ (.A(_01179_),
    .B(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hd__xor2_2 _08121_ (.A(_01207_),
    .B(_01208_),
    .X(_01213_));
 sky130_fd_sc_hd__xor2_1 _08122_ (.A(_01182_),
    .B(_01184_),
    .X(_01214_));
 sky130_fd_sc_hd__o22a_1 _08123_ (.A1(net143),
    .A2(net35),
    .B1(net33),
    .B2(net215),
    .X(_01215_));
 sky130_fd_sc_hd__xnor2_1 _08124_ (.A(net125),
    .B(_01215_),
    .Y(_01216_));
 sky130_fd_sc_hd__and2_1 _08125_ (.A(_01214_),
    .B(_01216_),
    .X(_01217_));
 sky130_fd_sc_hd__o22a_1 _08126_ (.A1(net287),
    .A2(net84),
    .B1(net80),
    .B2(net237),
    .X(_01218_));
 sky130_fd_sc_hd__xnor2_1 _08127_ (.A(net238),
    .B(_01218_),
    .Y(_01219_));
 sky130_fd_sc_hd__o22a_1 _08128_ (.A1(net151),
    .A2(net76),
    .B1(net72),
    .B2(net149),
    .X(_01220_));
 sky130_fd_sc_hd__xnor2_1 _08129_ (.A(net204),
    .B(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__nor2_1 _08130_ (.A(_01219_),
    .B(_01221_),
    .Y(_01222_));
 sky130_fd_sc_hd__xor2_1 _08131_ (.A(_01214_),
    .B(_01216_),
    .X(_01223_));
 sky130_fd_sc_hd__and2_1 _08132_ (.A(_01222_),
    .B(_01223_),
    .X(_01224_));
 sky130_fd_sc_hd__a21o_1 _08133_ (.A1(_01222_),
    .A2(_01223_),
    .B1(_01217_),
    .X(_01225_));
 sky130_fd_sc_hd__o22a_1 _08134_ (.A1(net131),
    .A2(net115),
    .B1(net109),
    .B2(net133),
    .X(_01226_));
 sky130_fd_sc_hd__xnor2_1 _08135_ (.A(net180),
    .B(_01226_),
    .Y(_01227_));
 sky130_fd_sc_hd__o22a_1 _08136_ (.A1(net153),
    .A2(net119),
    .B1(net72),
    .B2(net155),
    .X(_01228_));
 sky130_fd_sc_hd__xnor2_1 _08137_ (.A(net208),
    .B(_01228_),
    .Y(_01229_));
 sky130_fd_sc_hd__o22a_1 _08138_ (.A1(net147),
    .A2(net117),
    .B1(net111),
    .B2(net145),
    .X(_01230_));
 sky130_fd_sc_hd__xnor2_1 _08139_ (.A(net201),
    .B(_01230_),
    .Y(_01231_));
 sky130_fd_sc_hd__xnor2_1 _08140_ (.A(_01227_),
    .B(_01229_),
    .Y(_01232_));
 sky130_fd_sc_hd__or2_1 _08141_ (.A(_01231_),
    .B(_01232_),
    .X(_01233_));
 sky130_fd_sc_hd__o21a_2 _08142_ (.A1(_01227_),
    .A2(_01229_),
    .B1(_01233_),
    .X(_01234_));
 sky130_fd_sc_hd__o21ba_1 _08143_ (.A1(_01217_),
    .A2(_01224_),
    .B1_N(_01234_),
    .X(_01235_));
 sky130_fd_sc_hd__o22a_1 _08144_ (.A1(net114),
    .A2(net107),
    .B1(net105),
    .B2(net108),
    .X(_01236_));
 sky130_fd_sc_hd__xnor2_2 _08145_ (.A(net136),
    .B(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__o22a_1 _08146_ (.A1(net141),
    .A2(net79),
    .B1(net75),
    .B2(net140),
    .X(_01238_));
 sky130_fd_sc_hd__xnor2_2 _08147_ (.A(net123),
    .B(_01238_),
    .Y(_01239_));
 sky130_fd_sc_hd__o22a_1 _08148_ (.A1(net129),
    .A2(net87),
    .B1(net83),
    .B2(net127),
    .X(_01240_));
 sky130_fd_sc_hd__xnor2_1 _08149_ (.A(net138),
    .B(_01240_),
    .Y(_01241_));
 sky130_fd_sc_hd__xnor2_1 _08150_ (.A(_01237_),
    .B(_01239_),
    .Y(_01242_));
 sky130_fd_sc_hd__or2_1 _08151_ (.A(_01241_),
    .B(_01242_),
    .X(_01243_));
 sky130_fd_sc_hd__o21ai_4 _08152_ (.A1(_01237_),
    .A2(_01239_),
    .B1(_01243_),
    .Y(_01244_));
 sky130_fd_sc_hd__xnor2_4 _08153_ (.A(_01225_),
    .B(_01234_),
    .Y(_01245_));
 sky130_fd_sc_hd__a21o_1 _08154_ (.A1(_01244_),
    .A2(_01245_),
    .B1(_01235_),
    .X(_01246_));
 sky130_fd_sc_hd__xnor2_2 _08155_ (.A(_01190_),
    .B(_01191_),
    .Y(_01247_));
 sky130_fd_sc_hd__and2_1 _08156_ (.A(_01199_),
    .B(_01200_),
    .X(_01248_));
 sky130_fd_sc_hd__nor2_1 _08157_ (.A(_01201_),
    .B(_01248_),
    .Y(_01249_));
 sky130_fd_sc_hd__xnor2_1 _08158_ (.A(_01247_),
    .B(_01249_),
    .Y(_01250_));
 sky130_fd_sc_hd__xnor2_1 _08159_ (.A(_01204_),
    .B(_01206_),
    .Y(_01251_));
 sky130_fd_sc_hd__nor2_1 _08160_ (.A(_01250_),
    .B(_01251_),
    .Y(_01252_));
 sky130_fd_sc_hd__a21oi_2 _08161_ (.A1(_01247_),
    .A2(_01249_),
    .B1(_01252_),
    .Y(_01253_));
 sky130_fd_sc_hd__xor2_2 _08162_ (.A(_01213_),
    .B(_01246_),
    .X(_01254_));
 sky130_fd_sc_hd__nand2b_1 _08163_ (.A_N(_01253_),
    .B(_01254_),
    .Y(_01255_));
 sky130_fd_sc_hd__a21bo_1 _08164_ (.A1(_01213_),
    .A2(_01246_),
    .B1_N(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__xnor2_2 _08165_ (.A(_01171_),
    .B(_01212_),
    .Y(_01257_));
 sky130_fd_sc_hd__nand2b_1 _08166_ (.A_N(_01257_),
    .B(_01256_),
    .Y(_01258_));
 sky130_fd_sc_hd__o21ai_2 _08167_ (.A1(_01171_),
    .A2(_01212_),
    .B1(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hd__o21a_1 _08168_ (.A1(_01093_),
    .A2(_01094_),
    .B1(_01095_),
    .X(_01260_));
 sky130_fd_sc_hd__nor2_2 _08169_ (.A(_01096_),
    .B(_01260_),
    .Y(_01261_));
 sky130_fd_sc_hd__xnor2_2 _08170_ (.A(_01161_),
    .B(_01162_),
    .Y(_01262_));
 sky130_fd_sc_hd__and2_1 _08171_ (.A(_01261_),
    .B(_01262_),
    .X(_01263_));
 sky130_fd_sc_hd__xor2_2 _08172_ (.A(_01261_),
    .B(_01262_),
    .X(_01264_));
 sky130_fd_sc_hd__a21o_1 _08173_ (.A1(_01179_),
    .A2(_01211_),
    .B1(_01210_),
    .X(_01265_));
 sky130_fd_sc_hd__xor2_2 _08174_ (.A(_01264_),
    .B(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__nor2_1 _08175_ (.A(_01259_),
    .B(_01266_),
    .Y(_01267_));
 sky130_fd_sc_hd__nand2_1 _08176_ (.A(_01259_),
    .B(_01266_),
    .Y(_01268_));
 sky130_fd_sc_hd__xnor2_2 _08177_ (.A(_01259_),
    .B(_01266_),
    .Y(_01269_));
 sky130_fd_sc_hd__a21o_1 _08178_ (.A1(_01264_),
    .A2(_01265_),
    .B1(_01263_),
    .X(_01270_));
 sky130_fd_sc_hd__xnor2_2 _08179_ (.A(_01164_),
    .B(_01165_),
    .Y(_01271_));
 sky130_fd_sc_hd__nand2b_1 _08180_ (.A_N(_01271_),
    .B(_01270_),
    .Y(_01272_));
 sky130_fd_sc_hd__and2b_1 _08181_ (.A_N(_01270_),
    .B(_01271_),
    .X(_01273_));
 sky130_fd_sc_hd__xor2_1 _08182_ (.A(_01270_),
    .B(_01271_),
    .X(_01274_));
 sky130_fd_sc_hd__or2_1 _08183_ (.A(_01269_),
    .B(_01274_),
    .X(_01275_));
 sky130_fd_sc_hd__o21a_1 _08184_ (.A1(_01175_),
    .A2(_01176_),
    .B1(_01177_),
    .X(_01276_));
 sky130_fd_sc_hd__nor2_1 _08185_ (.A(_01178_),
    .B(_01276_),
    .Y(_01277_));
 sky130_fd_sc_hd__xnor2_2 _08186_ (.A(_01253_),
    .B(_01254_),
    .Y(_01278_));
 sky130_fd_sc_hd__and2_1 _08187_ (.A(_01277_),
    .B(_01278_),
    .X(_01279_));
 sky130_fd_sc_hd__xor2_2 _08188_ (.A(_01277_),
    .B(_01278_),
    .X(_01280_));
 sky130_fd_sc_hd__o22a_1 _08189_ (.A1(net133),
    .A2(net115),
    .B1(net114),
    .B2(net131),
    .X(_01281_));
 sky130_fd_sc_hd__xnor2_1 _08190_ (.A(net180),
    .B(_01281_),
    .Y(_01282_));
 sky130_fd_sc_hd__o22a_1 _08191_ (.A1(net155),
    .A2(net119),
    .B1(net117),
    .B2(net153),
    .X(_01283_));
 sky130_fd_sc_hd__xnor2_1 _08192_ (.A(net208),
    .B(_01283_),
    .Y(_01284_));
 sky130_fd_sc_hd__xnor2_1 _08193_ (.A(_01282_),
    .B(_01284_),
    .Y(_01285_));
 sky130_fd_sc_hd__o22a_1 _08194_ (.A1(net147),
    .A2(net111),
    .B1(net109),
    .B2(net145),
    .X(_01286_));
 sky130_fd_sc_hd__xnor2_1 _08195_ (.A(net201),
    .B(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__nor2_1 _08196_ (.A(_01285_),
    .B(_01287_),
    .Y(_01288_));
 sky130_fd_sc_hd__o21ba_1 _08197_ (.A1(_01282_),
    .A2(_01284_),
    .B1_N(_01288_),
    .X(_01289_));
 sky130_fd_sc_hd__xor2_1 _08198_ (.A(_01219_),
    .B(_01221_),
    .X(_01290_));
 sky130_fd_sc_hd__nor2_1 _08199_ (.A(net215),
    .B(net35),
    .Y(_01291_));
 sky130_fd_sc_hd__mux2_1 _08200_ (.A0(net125),
    .A1(_01290_),
    .S(_01291_),
    .X(_01292_));
 sky130_fd_sc_hd__and2b_1 _08201_ (.A_N(_01289_),
    .B(_01292_),
    .X(_01293_));
 sky130_fd_sc_hd__o22a_1 _08202_ (.A1(net108),
    .A2(net107),
    .B1(net105),
    .B2(net129),
    .X(_01294_));
 sky130_fd_sc_hd__xnor2_1 _08203_ (.A(net136),
    .B(_01294_),
    .Y(_01295_));
 sky130_fd_sc_hd__o22a_1 _08204_ (.A1(net140),
    .A2(net79),
    .B1(net75),
    .B2(net143),
    .X(_01296_));
 sky130_fd_sc_hd__xnor2_2 _08205_ (.A(net123),
    .B(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__o22a_1 _08206_ (.A1(net127),
    .A2(net87),
    .B1(net83),
    .B2(net141),
    .X(_01298_));
 sky130_fd_sc_hd__xnor2_1 _08207_ (.A(net138),
    .B(_01298_),
    .Y(_01299_));
 sky130_fd_sc_hd__xnor2_1 _08208_ (.A(_01295_),
    .B(_01297_),
    .Y(_01300_));
 sky130_fd_sc_hd__or2_1 _08209_ (.A(_01299_),
    .B(_01300_),
    .X(_01301_));
 sky130_fd_sc_hd__o21ai_2 _08210_ (.A1(_01295_),
    .A2(_01297_),
    .B1(_01301_),
    .Y(_01302_));
 sky130_fd_sc_hd__xnor2_2 _08211_ (.A(_01289_),
    .B(_01292_),
    .Y(_01303_));
 sky130_fd_sc_hd__a21oi_4 _08212_ (.A1(_01302_),
    .A2(_01303_),
    .B1(_01293_),
    .Y(_01304_));
 sky130_fd_sc_hd__xor2_4 _08213_ (.A(_01244_),
    .B(_01245_),
    .X(_01305_));
 sky130_fd_sc_hd__and2b_1 _08214_ (.A_N(_01304_),
    .B(_01305_),
    .X(_01306_));
 sky130_fd_sc_hd__nor2_1 _08215_ (.A(_01222_),
    .B(_01223_),
    .Y(_01307_));
 sky130_fd_sc_hd__or2_1 _08216_ (.A(_01224_),
    .B(_01307_),
    .X(_01308_));
 sky130_fd_sc_hd__nand2_1 _08217_ (.A(_01231_),
    .B(_01232_),
    .Y(_01309_));
 sky130_fd_sc_hd__and2_1 _08218_ (.A(_01233_),
    .B(_01309_),
    .X(_01310_));
 sky130_fd_sc_hd__and2b_1 _08219_ (.A_N(_01308_),
    .B(_01310_),
    .X(_01311_));
 sky130_fd_sc_hd__nand2_1 _08220_ (.A(_01241_),
    .B(_01242_),
    .Y(_01312_));
 sky130_fd_sc_hd__and2_1 _08221_ (.A(_01243_),
    .B(_01312_),
    .X(_01313_));
 sky130_fd_sc_hd__xnor2_1 _08222_ (.A(_01308_),
    .B(_01310_),
    .Y(_01314_));
 sky130_fd_sc_hd__a21o_2 _08223_ (.A1(_01313_),
    .A2(_01314_),
    .B1(_01311_),
    .X(_01315_));
 sky130_fd_sc_hd__xnor2_4 _08224_ (.A(_01304_),
    .B(_01305_),
    .Y(_01316_));
 sky130_fd_sc_hd__a21o_1 _08225_ (.A1(_01315_),
    .A2(_01316_),
    .B1(_01306_),
    .X(_01317_));
 sky130_fd_sc_hd__a21oi_2 _08226_ (.A1(_01280_),
    .A2(_01317_),
    .B1(_01279_),
    .Y(_01318_));
 sky130_fd_sc_hd__xor2_2 _08227_ (.A(_01256_),
    .B(_01257_),
    .X(_01319_));
 sky130_fd_sc_hd__and2_1 _08228_ (.A(_01318_),
    .B(_01319_),
    .X(_01320_));
 sky130_fd_sc_hd__or2_1 _08229_ (.A(_01318_),
    .B(_01319_),
    .X(_01321_));
 sky130_fd_sc_hd__and2_1 _08230_ (.A(_01250_),
    .B(_01251_),
    .X(_01322_));
 sky130_fd_sc_hd__or2_2 _08231_ (.A(_01252_),
    .B(_01322_),
    .X(_01323_));
 sky130_fd_sc_hd__xnor2_4 _08232_ (.A(_01315_),
    .B(_01316_),
    .Y(_01324_));
 sky130_fd_sc_hd__nor2_1 _08233_ (.A(_01323_),
    .B(_01324_),
    .Y(_01325_));
 sky130_fd_sc_hd__xor2_4 _08234_ (.A(_01323_),
    .B(_01324_),
    .X(_01326_));
 sky130_fd_sc_hd__xnor2_1 _08235_ (.A(_01302_),
    .B(_01303_),
    .Y(_01327_));
 sky130_fd_sc_hd__o22a_1 _08236_ (.A1(net141),
    .A2(net87),
    .B1(net83),
    .B2(net140),
    .X(_01328_));
 sky130_fd_sc_hd__xnor2_1 _08237_ (.A(net138),
    .B(_01328_),
    .Y(_01329_));
 sky130_fd_sc_hd__o22a_1 _08238_ (.A1(net143),
    .A2(net79),
    .B1(net75),
    .B2(net215),
    .X(_01330_));
 sky130_fd_sc_hd__xnor2_1 _08239_ (.A(net123),
    .B(_01330_),
    .Y(_01331_));
 sky130_fd_sc_hd__nor2_1 _08240_ (.A(_01329_),
    .B(_01331_),
    .Y(_01332_));
 sky130_fd_sc_hd__o22a_1 _08241_ (.A1(net287),
    .A2(net80),
    .B1(net76),
    .B2(net237),
    .X(_01333_));
 sky130_fd_sc_hd__xnor2_2 _08242_ (.A(net238),
    .B(_01333_),
    .Y(_01334_));
 sky130_fd_sc_hd__o22a_1 _08243_ (.A1(net155),
    .A2(net117),
    .B1(net111),
    .B2(net153),
    .X(_01335_));
 sky130_fd_sc_hd__xnor2_2 _08244_ (.A(net208),
    .B(_01335_),
    .Y(_01336_));
 sky130_fd_sc_hd__or2_1 _08245_ (.A(_01334_),
    .B(_01336_),
    .X(_01337_));
 sky130_fd_sc_hd__xnor2_2 _08246_ (.A(_01334_),
    .B(_01336_),
    .Y(_01338_));
 sky130_fd_sc_hd__o22a_1 _08247_ (.A1(net149),
    .A2(net119),
    .B1(net72),
    .B2(net151),
    .X(_01339_));
 sky130_fd_sc_hd__xnor2_2 _08248_ (.A(net204),
    .B(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__o21ai_1 _08249_ (.A1(_01338_),
    .A2(_01340_),
    .B1(_01337_),
    .Y(_01341_));
 sky130_fd_sc_hd__nand2_1 _08250_ (.A(_01332_),
    .B(_01341_),
    .Y(_01342_));
 sky130_fd_sc_hd__o22a_1 _08251_ (.A1(net129),
    .A2(net107),
    .B1(net105),
    .B2(net127),
    .X(_01343_));
 sky130_fd_sc_hd__xnor2_2 _08252_ (.A(net136),
    .B(_01343_),
    .Y(_01344_));
 sky130_fd_sc_hd__o22a_1 _08253_ (.A1(net145),
    .A2(net115),
    .B1(net109),
    .B2(net147),
    .X(_01345_));
 sky130_fd_sc_hd__xnor2_2 _08254_ (.A(net201),
    .B(_01345_),
    .Y(_01346_));
 sky130_fd_sc_hd__xor2_2 _08255_ (.A(_01344_),
    .B(_01346_),
    .X(_01347_));
 sky130_fd_sc_hd__o22a_1 _08256_ (.A1(net133),
    .A2(net114),
    .B1(net108),
    .B2(net131),
    .X(_01348_));
 sky130_fd_sc_hd__xnor2_2 _08257_ (.A(net180),
    .B(_01348_),
    .Y(_01349_));
 sky130_fd_sc_hd__nand2b_1 _08258_ (.A_N(_01349_),
    .B(_01347_),
    .Y(_01350_));
 sky130_fd_sc_hd__o21ai_2 _08259_ (.A1(_01344_),
    .A2(_01346_),
    .B1(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__xor2_1 _08260_ (.A(_01332_),
    .B(_01341_),
    .X(_01352_));
 sky130_fd_sc_hd__a21boi_1 _08261_ (.A1(_01351_),
    .A2(_01352_),
    .B1_N(_01342_),
    .Y(_01353_));
 sky130_fd_sc_hd__nor2_1 _08262_ (.A(_01327_),
    .B(_01353_),
    .Y(_01354_));
 sky130_fd_sc_hd__and2_1 _08263_ (.A(_01285_),
    .B(_01287_),
    .X(_01355_));
 sky130_fd_sc_hd__nor2_1 _08264_ (.A(_01288_),
    .B(_01355_),
    .Y(_01356_));
 sky130_fd_sc_hd__xnor2_1 _08265_ (.A(_01290_),
    .B(_01291_),
    .Y(_01357_));
 sky130_fd_sc_hd__and2b_1 _08266_ (.A_N(_01357_),
    .B(_01356_),
    .X(_01358_));
 sky130_fd_sc_hd__and2b_1 _08267_ (.A_N(_01356_),
    .B(_01357_),
    .X(_01359_));
 sky130_fd_sc_hd__nor2_1 _08268_ (.A(_01358_),
    .B(_01359_),
    .Y(_01360_));
 sky130_fd_sc_hd__nand2_1 _08269_ (.A(_01299_),
    .B(_01300_),
    .Y(_01361_));
 sky130_fd_sc_hd__and2_1 _08270_ (.A(_01301_),
    .B(_01361_),
    .X(_01362_));
 sky130_fd_sc_hd__a21o_1 _08271_ (.A1(_01360_),
    .A2(_01362_),
    .B1(_01358_),
    .X(_01363_));
 sky130_fd_sc_hd__xor2_1 _08272_ (.A(_01327_),
    .B(_01353_),
    .X(_01364_));
 sky130_fd_sc_hd__a21o_1 _08273_ (.A1(_01363_),
    .A2(_01364_),
    .B1(_01354_),
    .X(_01365_));
 sky130_fd_sc_hd__a21o_1 _08274_ (.A1(_01326_),
    .A2(_01365_),
    .B1(_01325_),
    .X(_01366_));
 sky130_fd_sc_hd__xor2_2 _08275_ (.A(_01280_),
    .B(_01317_),
    .X(_01367_));
 sky130_fd_sc_hd__nand2_1 _08276_ (.A(_01366_),
    .B(_01367_),
    .Y(_01368_));
 sky130_fd_sc_hd__a21o_1 _08277_ (.A1(_01321_),
    .A2(_01368_),
    .B1(_01320_),
    .X(_01369_));
 sky130_fd_sc_hd__xnor2_2 _08278_ (.A(_01318_),
    .B(_01319_),
    .Y(_01370_));
 sky130_fd_sc_hd__nor2_1 _08279_ (.A(_01366_),
    .B(_01367_),
    .Y(_01371_));
 sky130_fd_sc_hd__xnor2_2 _08280_ (.A(_01366_),
    .B(_01367_),
    .Y(_01372_));
 sky130_fd_sc_hd__or2_1 _08281_ (.A(_01370_),
    .B(_01372_),
    .X(_01373_));
 sky130_fd_sc_hd__xor2_4 _08282_ (.A(_01326_),
    .B(_01365_),
    .X(_01374_));
 sky130_fd_sc_hd__xnor2_1 _08283_ (.A(_01313_),
    .B(_01314_),
    .Y(_01375_));
 sky130_fd_sc_hd__xnor2_1 _08284_ (.A(_01363_),
    .B(_01364_),
    .Y(_01376_));
 sky130_fd_sc_hd__nor2_1 _08285_ (.A(_01375_),
    .B(_01376_),
    .Y(_01377_));
 sky130_fd_sc_hd__xnor2_1 _08286_ (.A(_01351_),
    .B(_01352_),
    .Y(_01378_));
 sky130_fd_sc_hd__o22a_2 _08287_ (.A1(net140),
    .A2(net87),
    .B1(net83),
    .B2(net143),
    .X(_01379_));
 sky130_fd_sc_hd__xnor2_4 _08288_ (.A(net138),
    .B(_01379_),
    .Y(_01380_));
 sky130_fd_sc_hd__nor2_2 _08289_ (.A(net215),
    .B(net79),
    .Y(_01381_));
 sky130_fd_sc_hd__xnor2_4 _08290_ (.A(net123),
    .B(_01381_),
    .Y(_01382_));
 sky130_fd_sc_hd__nand2b_1 _08291_ (.A_N(_01380_),
    .B(_01382_),
    .Y(_01383_));
 sky130_fd_sc_hd__o22a_2 _08292_ (.A1(net287),
    .A2(net76),
    .B1(net72),
    .B2(net237),
    .X(_01384_));
 sky130_fd_sc_hd__xnor2_4 _08293_ (.A(net238),
    .B(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__o22a_1 _08294_ (.A1(net155),
    .A2(net111),
    .B1(net109),
    .B2(net153),
    .X(_01386_));
 sky130_fd_sc_hd__xnor2_2 _08295_ (.A(net208),
    .B(_01386_),
    .Y(_01387_));
 sky130_fd_sc_hd__or2_1 _08296_ (.A(_01385_),
    .B(_01387_),
    .X(_01388_));
 sky130_fd_sc_hd__xnor2_4 _08297_ (.A(_01385_),
    .B(_01387_),
    .Y(_01389_));
 sky130_fd_sc_hd__o22a_2 _08298_ (.A1(net151),
    .A2(net119),
    .B1(net117),
    .B2(net149),
    .X(_01390_));
 sky130_fd_sc_hd__xnor2_4 _08299_ (.A(net204),
    .B(_01390_),
    .Y(_01391_));
 sky130_fd_sc_hd__o21a_1 _08300_ (.A1(_01389_),
    .A2(_01391_),
    .B1(_01388_),
    .X(_01392_));
 sky130_fd_sc_hd__nor2_1 _08301_ (.A(_01383_),
    .B(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__o22a_1 _08302_ (.A1(net127),
    .A2(net107),
    .B1(net105),
    .B2(net141),
    .X(_01394_));
 sky130_fd_sc_hd__xnor2_2 _08303_ (.A(net136),
    .B(_01394_),
    .Y(_01395_));
 sky130_fd_sc_hd__o22a_1 _08304_ (.A1(net147),
    .A2(net115),
    .B1(net114),
    .B2(net145),
    .X(_01396_));
 sky130_fd_sc_hd__xnor2_2 _08305_ (.A(net201),
    .B(_01396_),
    .Y(_01397_));
 sky130_fd_sc_hd__xor2_2 _08306_ (.A(_01395_),
    .B(_01397_),
    .X(_01398_));
 sky130_fd_sc_hd__o22a_1 _08307_ (.A1(net131),
    .A2(net129),
    .B1(net108),
    .B2(net133),
    .X(_01399_));
 sky130_fd_sc_hd__xnor2_2 _08308_ (.A(net180),
    .B(_01399_),
    .Y(_01400_));
 sky130_fd_sc_hd__nand2b_1 _08309_ (.A_N(_01400_),
    .B(_01398_),
    .Y(_01401_));
 sky130_fd_sc_hd__o21ai_2 _08310_ (.A1(_01395_),
    .A2(_01397_),
    .B1(_01401_),
    .Y(_01402_));
 sky130_fd_sc_hd__xor2_2 _08311_ (.A(_01383_),
    .B(_01392_),
    .X(_01403_));
 sky130_fd_sc_hd__a21oi_2 _08312_ (.A1(_01402_),
    .A2(_01403_),
    .B1(_01393_),
    .Y(_01404_));
 sky130_fd_sc_hd__xnor2_2 _08313_ (.A(_01338_),
    .B(_01340_),
    .Y(_01405_));
 sky130_fd_sc_hd__and2_1 _08314_ (.A(_01329_),
    .B(_01331_),
    .X(_01406_));
 sky130_fd_sc_hd__or2_1 _08315_ (.A(_01332_),
    .B(_01406_),
    .X(_01407_));
 sky130_fd_sc_hd__xnor2_2 _08316_ (.A(_01405_),
    .B(_01407_),
    .Y(_01408_));
 sky130_fd_sc_hd__xnor2_2 _08317_ (.A(_01347_),
    .B(_01349_),
    .Y(_01409_));
 sky130_fd_sc_hd__nand2b_1 _08318_ (.A_N(_01408_),
    .B(_01409_),
    .Y(_01410_));
 sky130_fd_sc_hd__o21ai_1 _08319_ (.A1(_01405_),
    .A2(_01407_),
    .B1(_01410_),
    .Y(_01411_));
 sky130_fd_sc_hd__xnor2_1 _08320_ (.A(_01378_),
    .B(_01404_),
    .Y(_01412_));
 sky130_fd_sc_hd__and2b_1 _08321_ (.A_N(_01412_),
    .B(_01411_),
    .X(_01413_));
 sky130_fd_sc_hd__o21bai_2 _08322_ (.A1(_01378_),
    .A2(_01404_),
    .B1_N(_01413_),
    .Y(_01414_));
 sky130_fd_sc_hd__xor2_1 _08323_ (.A(_01375_),
    .B(_01376_),
    .X(_01415_));
 sky130_fd_sc_hd__a21o_2 _08324_ (.A1(_01414_),
    .A2(_01415_),
    .B1(_01377_),
    .X(_01416_));
 sky130_fd_sc_hd__nor2_1 _08325_ (.A(_01374_),
    .B(_01416_),
    .Y(_01417_));
 sky130_fd_sc_hd__nand2_1 _08326_ (.A(_01374_),
    .B(_01416_),
    .Y(_01418_));
 sky130_fd_sc_hd__xnor2_1 _08327_ (.A(_01360_),
    .B(_01362_),
    .Y(_01419_));
 sky130_fd_sc_hd__xor2_1 _08328_ (.A(_01411_),
    .B(_01412_),
    .X(_01420_));
 sky130_fd_sc_hd__or2_1 _08329_ (.A(_01419_),
    .B(_01420_),
    .X(_01421_));
 sky130_fd_sc_hd__o22a_1 _08330_ (.A1(net147),
    .A2(net114),
    .B1(net108),
    .B2(net145),
    .X(_01422_));
 sky130_fd_sc_hd__xnor2_2 _08331_ (.A(net201),
    .B(_01422_),
    .Y(_01423_));
 sky130_fd_sc_hd__o22a_1 _08332_ (.A1(net133),
    .A2(net129),
    .B1(net127),
    .B2(net131),
    .X(_01424_));
 sky130_fd_sc_hd__xnor2_2 _08333_ (.A(net180),
    .B(_01424_),
    .Y(_01425_));
 sky130_fd_sc_hd__or3_1 _08334_ (.A(net123),
    .B(_01423_),
    .C(_01425_),
    .X(_01426_));
 sky130_fd_sc_hd__a22o_1 _08335_ (.A1(_06519_),
    .A2(_00287_),
    .B1(_00366_),
    .B2(net292),
    .X(_01427_));
 sky130_fd_sc_hd__xnor2_4 _08336_ (.A(net240),
    .B(_01427_),
    .Y(_01428_));
 sky130_fd_sc_hd__o22a_1 _08337_ (.A1(net153),
    .A2(net115),
    .B1(net109),
    .B2(net155),
    .X(_01429_));
 sky130_fd_sc_hd__xnor2_1 _08338_ (.A(net208),
    .B(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__or2_1 _08339_ (.A(_01428_),
    .B(_01430_),
    .X(_01431_));
 sky130_fd_sc_hd__o22a_1 _08340_ (.A1(net151),
    .A2(net117),
    .B1(net111),
    .B2(net149),
    .X(_01432_));
 sky130_fd_sc_hd__xnor2_1 _08341_ (.A(net204),
    .B(_01432_),
    .Y(_01433_));
 sky130_fd_sc_hd__xnor2_1 _08342_ (.A(_01428_),
    .B(_01430_),
    .Y(_01434_));
 sky130_fd_sc_hd__o21a_1 _08343_ (.A1(_01433_),
    .A2(_01434_),
    .B1(_01431_),
    .X(_01435_));
 sky130_fd_sc_hd__o21ai_1 _08344_ (.A1(_01423_),
    .A2(_01425_),
    .B1(net123),
    .Y(_01436_));
 sky130_fd_sc_hd__nand2_1 _08345_ (.A(_01426_),
    .B(_01436_),
    .Y(_01437_));
 sky130_fd_sc_hd__o21ai_2 _08346_ (.A1(_01435_),
    .A2(_01437_),
    .B1(_01426_),
    .Y(_01438_));
 sky130_fd_sc_hd__xnor2_2 _08347_ (.A(_01402_),
    .B(_01403_),
    .Y(_01439_));
 sky130_fd_sc_hd__nand2b_1 _08348_ (.A_N(_01439_),
    .B(_01438_),
    .Y(_01440_));
 sky130_fd_sc_hd__xor2_4 _08349_ (.A(_01389_),
    .B(_01391_),
    .X(_01441_));
 sky130_fd_sc_hd__xnor2_4 _08350_ (.A(_01380_),
    .B(_01382_),
    .Y(_01442_));
 sky130_fd_sc_hd__xnor2_4 _08351_ (.A(_01441_),
    .B(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__xnor2_2 _08352_ (.A(_01398_),
    .B(_01400_),
    .Y(_01444_));
 sky130_fd_sc_hd__and2b_1 _08353_ (.A_N(_01443_),
    .B(_01444_),
    .X(_01445_));
 sky130_fd_sc_hd__a21o_1 _08354_ (.A1(_01441_),
    .A2(_01442_),
    .B1(_01445_),
    .X(_01446_));
 sky130_fd_sc_hd__xor2_2 _08355_ (.A(_01438_),
    .B(_01439_),
    .X(_01447_));
 sky130_fd_sc_hd__nand2b_1 _08356_ (.A_N(_01447_),
    .B(_01446_),
    .Y(_01448_));
 sky130_fd_sc_hd__nand2_1 _08357_ (.A(_01440_),
    .B(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hd__xor2_1 _08358_ (.A(_01419_),
    .B(_01420_),
    .X(_01450_));
 sky130_fd_sc_hd__nand2_1 _08359_ (.A(_01449_),
    .B(_01450_),
    .Y(_01451_));
 sky130_fd_sc_hd__xnor2_1 _08360_ (.A(_01414_),
    .B(_01415_),
    .Y(_01452_));
 sky130_fd_sc_hd__a21oi_1 _08361_ (.A1(_01421_),
    .A2(_01451_),
    .B1(_01452_),
    .Y(_01453_));
 sky130_fd_sc_hd__inv_2 _08362_ (.A(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__a21o_1 _08363_ (.A1(_01418_),
    .A2(_01454_),
    .B1(_01417_),
    .X(_01455_));
 sky130_fd_sc_hd__xnor2_2 _08364_ (.A(_01408_),
    .B(_01409_),
    .Y(_01456_));
 sky130_fd_sc_hd__xnor2_2 _08365_ (.A(_01446_),
    .B(_01447_),
    .Y(_01457_));
 sky130_fd_sc_hd__nand2_1 _08366_ (.A(_01456_),
    .B(_01457_),
    .Y(_01458_));
 sky130_fd_sc_hd__xor2_2 _08367_ (.A(_01435_),
    .B(_01437_),
    .X(_01459_));
 sky130_fd_sc_hd__o22a_1 _08368_ (.A1(net287),
    .A2(net119),
    .B1(net117),
    .B2(net237),
    .X(_01460_));
 sky130_fd_sc_hd__xnor2_2 _08369_ (.A(net238),
    .B(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__o22a_1 _08370_ (.A1(net155),
    .A2(net115),
    .B1(net114),
    .B2(net153),
    .X(_01462_));
 sky130_fd_sc_hd__xnor2_2 _08371_ (.A(net208),
    .B(_01462_),
    .Y(_01463_));
 sky130_fd_sc_hd__or2_1 _08372_ (.A(_01461_),
    .B(_01463_),
    .X(_01464_));
 sky130_fd_sc_hd__o22a_1 _08373_ (.A1(net151),
    .A2(net111),
    .B1(net109),
    .B2(net149),
    .X(_01465_));
 sky130_fd_sc_hd__xnor2_2 _08374_ (.A(net204),
    .B(_01465_),
    .Y(_01466_));
 sky130_fd_sc_hd__xnor2_2 _08375_ (.A(_01461_),
    .B(_01463_),
    .Y(_01467_));
 sky130_fd_sc_hd__nor2_1 _08376_ (.A(_01466_),
    .B(_01467_),
    .Y(_01468_));
 sky130_fd_sc_hd__o21ai_2 _08377_ (.A1(_01466_),
    .A2(_01467_),
    .B1(_01464_),
    .Y(_01469_));
 sky130_fd_sc_hd__o22a_2 _08378_ (.A1(net141),
    .A2(net106),
    .B1(net105),
    .B2(_00264_),
    .X(_01470_));
 sky130_fd_sc_hd__xnor2_4 _08379_ (.A(_00342_),
    .B(_01470_),
    .Y(_01471_));
 sky130_fd_sc_hd__and2_1 _08380_ (.A(_01469_),
    .B(_01471_),
    .X(_01472_));
 sky130_fd_sc_hd__o22a_1 _08381_ (.A1(net143),
    .A2(net87),
    .B1(net83),
    .B2(net215),
    .X(_01473_));
 sky130_fd_sc_hd__xnor2_2 _08382_ (.A(net138),
    .B(_01473_),
    .Y(_01474_));
 sky130_fd_sc_hd__inv_2 _08383_ (.A(_01474_),
    .Y(_01475_));
 sky130_fd_sc_hd__xor2_2 _08384_ (.A(_01469_),
    .B(_01471_),
    .X(_01476_));
 sky130_fd_sc_hd__a21oi_2 _08385_ (.A1(_01475_),
    .A2(_01476_),
    .B1(_01472_),
    .Y(_01477_));
 sky130_fd_sc_hd__nand2b_1 _08386_ (.A_N(_01477_),
    .B(_01459_),
    .Y(_01478_));
 sky130_fd_sc_hd__o22a_1 _08387_ (.A1(net145),
    .A2(net129),
    .B1(net108),
    .B2(net147),
    .X(_01479_));
 sky130_fd_sc_hd__xnor2_1 _08388_ (.A(net201),
    .B(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__o22a_1 _08389_ (.A1(net133),
    .A2(net127),
    .B1(net141),
    .B2(net131),
    .X(_01481_));
 sky130_fd_sc_hd__xnor2_1 _08390_ (.A(net180),
    .B(_01481_),
    .Y(_01482_));
 sky130_fd_sc_hd__or2_1 _08391_ (.A(_01480_),
    .B(_01482_),
    .X(_01483_));
 sky130_fd_sc_hd__xnor2_2 _08392_ (.A(_01423_),
    .B(_01425_),
    .Y(_01484_));
 sky130_fd_sc_hd__xnor2_1 _08393_ (.A(_01433_),
    .B(_01434_),
    .Y(_01485_));
 sky130_fd_sc_hd__xnor2_1 _08394_ (.A(_01483_),
    .B(_01484_),
    .Y(_01486_));
 sky130_fd_sc_hd__or2_1 _08395_ (.A(_01485_),
    .B(_01486_),
    .X(_01487_));
 sky130_fd_sc_hd__o21ai_2 _08396_ (.A1(_01483_),
    .A2(_01484_),
    .B1(_01487_),
    .Y(_01488_));
 sky130_fd_sc_hd__xor2_2 _08397_ (.A(_01459_),
    .B(_01477_),
    .X(_01489_));
 sky130_fd_sc_hd__nand2b_1 _08398_ (.A_N(_01489_),
    .B(_01488_),
    .Y(_01490_));
 sky130_fd_sc_hd__nand2_1 _08399_ (.A(_01478_),
    .B(_01490_),
    .Y(_01491_));
 sky130_fd_sc_hd__xnor2_2 _08400_ (.A(_01456_),
    .B(_01457_),
    .Y(_01492_));
 sky130_fd_sc_hd__nand2b_1 _08401_ (.A_N(_01492_),
    .B(_01491_),
    .Y(_01493_));
 sky130_fd_sc_hd__xnor2_1 _08402_ (.A(_01449_),
    .B(_01450_),
    .Y(_01494_));
 sky130_fd_sc_hd__and3_1 _08403_ (.A(_01458_),
    .B(_01493_),
    .C(_01494_),
    .X(_01495_));
 sky130_fd_sc_hd__a21o_1 _08404_ (.A1(_01458_),
    .A2(_01493_),
    .B1(_01494_),
    .X(_01496_));
 sky130_fd_sc_hd__xor2_4 _08405_ (.A(_01443_),
    .B(_01444_),
    .X(_01497_));
 sky130_fd_sc_hd__xor2_2 _08406_ (.A(_01488_),
    .B(_01489_),
    .X(_01498_));
 sky130_fd_sc_hd__xor2_1 _08407_ (.A(_01497_),
    .B(_01498_),
    .X(_01499_));
 sky130_fd_sc_hd__xnor2_2 _08408_ (.A(_01474_),
    .B(_01476_),
    .Y(_01500_));
 sky130_fd_sc_hd__o22a_1 _08409_ (.A1(net140),
    .A2(net107),
    .B1(net105),
    .B2(net143),
    .X(_01501_));
 sky130_fd_sc_hd__xnor2_1 _08410_ (.A(net136),
    .B(_01501_),
    .Y(_01502_));
 sky130_fd_sc_hd__nor2_1 _08411_ (.A(net215),
    .B(net87),
    .Y(_01503_));
 sky130_fd_sc_hd__nand2_1 _08412_ (.A(_01502_),
    .B(_01503_),
    .Y(_01504_));
 sky130_fd_sc_hd__o21a_1 _08413_ (.A1(_00339_),
    .A2(_01503_),
    .B1(_01504_),
    .X(_01505_));
 sky130_fd_sc_hd__nand2_1 _08414_ (.A(_01500_),
    .B(_01505_),
    .Y(_01506_));
 sky130_fd_sc_hd__o22a_1 _08415_ (.A1(net287),
    .A2(net117),
    .B1(net111),
    .B2(net237),
    .X(_01507_));
 sky130_fd_sc_hd__xnor2_1 _08416_ (.A(net238),
    .B(_01507_),
    .Y(_01508_));
 sky130_fd_sc_hd__o22a_1 _08417_ (.A1(net149),
    .A2(net115),
    .B1(net109),
    .B2(net151),
    .X(_01509_));
 sky130_fd_sc_hd__xnor2_1 _08418_ (.A(net204),
    .B(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hd__or2_2 _08419_ (.A(_01508_),
    .B(_01510_),
    .X(_01511_));
 sky130_fd_sc_hd__nand2_1 _08420_ (.A(_01480_),
    .B(_01482_),
    .Y(_01512_));
 sky130_fd_sc_hd__nand2_1 _08421_ (.A(_01483_),
    .B(_01512_),
    .Y(_01513_));
 sky130_fd_sc_hd__or2_1 _08422_ (.A(_01511_),
    .B(_01513_),
    .X(_01514_));
 sky130_fd_sc_hd__xnor2_2 _08423_ (.A(_01511_),
    .B(_01513_),
    .Y(_01515_));
 sky130_fd_sc_hd__and2_1 _08424_ (.A(_01466_),
    .B(_01467_),
    .X(_01516_));
 sky130_fd_sc_hd__nor2_1 _08425_ (.A(_01468_),
    .B(_01516_),
    .Y(_01517_));
 sky130_fd_sc_hd__o31a_1 _08426_ (.A1(_01468_),
    .A2(_01515_),
    .A3(_01516_),
    .B1(_01514_),
    .X(_01518_));
 sky130_fd_sc_hd__xnor2_2 _08427_ (.A(_01500_),
    .B(_01505_),
    .Y(_01519_));
 sky130_fd_sc_hd__o21a_1 _08428_ (.A1(_01518_),
    .A2(_01519_),
    .B1(_01506_),
    .X(_01520_));
 sky130_fd_sc_hd__and2b_1 _08429_ (.A_N(_01520_),
    .B(_01499_),
    .X(_01521_));
 sky130_fd_sc_hd__o21bai_4 _08430_ (.A1(_01497_),
    .A2(_01498_),
    .B1_N(_01521_),
    .Y(_01522_));
 sky130_fd_sc_hd__xnor2_2 _08431_ (.A(_01491_),
    .B(_01492_),
    .Y(_01523_));
 sky130_fd_sc_hd__nand2_1 _08432_ (.A(_01522_),
    .B(_01523_),
    .Y(_01524_));
 sky130_fd_sc_hd__nand2b_1 _08433_ (.A_N(_01495_),
    .B(_01496_),
    .Y(_01525_));
 sky130_fd_sc_hd__xnor2_1 _08434_ (.A(_01522_),
    .B(_01523_),
    .Y(_01526_));
 sky130_fd_sc_hd__xor2_1 _08435_ (.A(_01499_),
    .B(_01520_),
    .X(_01527_));
 sky130_fd_sc_hd__nand2_1 _08436_ (.A(_01485_),
    .B(_01486_),
    .Y(_01528_));
 sky130_fd_sc_hd__nand2_1 _08437_ (.A(_01487_),
    .B(_01528_),
    .Y(_01529_));
 sky130_fd_sc_hd__xnor2_2 _08438_ (.A(_01518_),
    .B(_01519_),
    .Y(_01530_));
 sky130_fd_sc_hd__or2_1 _08439_ (.A(_01529_),
    .B(_01530_),
    .X(_01531_));
 sky130_fd_sc_hd__o22a_1 _08440_ (.A1(net133),
    .A2(net141),
    .B1(net140),
    .B2(net131),
    .X(_01532_));
 sky130_fd_sc_hd__xnor2_1 _08441_ (.A(net180),
    .B(_01532_),
    .Y(_01533_));
 sky130_fd_sc_hd__o22a_1 _08442_ (.A1(net156),
    .A2(net114),
    .B1(net108),
    .B2(net153),
    .X(_01534_));
 sky130_fd_sc_hd__xnor2_1 _08443_ (.A(net208),
    .B(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hd__or2_1 _08444_ (.A(_01533_),
    .B(_01535_),
    .X(_01536_));
 sky130_fd_sc_hd__o22a_1 _08445_ (.A1(net147),
    .A2(net129),
    .B1(net127),
    .B2(net145),
    .X(_01537_));
 sky130_fd_sc_hd__xnor2_1 _08446_ (.A(net201),
    .B(_01537_),
    .Y(_01538_));
 sky130_fd_sc_hd__xnor2_1 _08447_ (.A(_01533_),
    .B(_01535_),
    .Y(_01539_));
 sky130_fd_sc_hd__o21a_1 _08448_ (.A1(_01538_),
    .A2(_01539_),
    .B1(_01536_),
    .X(_01540_));
 sky130_fd_sc_hd__or2_1 _08449_ (.A(_01502_),
    .B(_01503_),
    .X(_01541_));
 sky130_fd_sc_hd__nand2_1 _08450_ (.A(_01504_),
    .B(_01541_),
    .Y(_01542_));
 sky130_fd_sc_hd__nand2b_1 _08451_ (.A_N(_01540_),
    .B(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__xnor2_1 _08452_ (.A(_01508_),
    .B(_01510_),
    .Y(_01544_));
 sky130_fd_sc_hd__o22a_1 _08453_ (.A1(net143),
    .A2(net107),
    .B1(net105),
    .B2(net215),
    .X(_01545_));
 sky130_fd_sc_hd__xnor2_1 _08454_ (.A(net136),
    .B(_01545_),
    .Y(_01546_));
 sky130_fd_sc_hd__o22a_1 _08455_ (.A1(net151),
    .A2(net115),
    .B1(net114),
    .B2(net149),
    .X(_01547_));
 sky130_fd_sc_hd__xnor2_1 _08456_ (.A(net204),
    .B(_01547_),
    .Y(_01548_));
 sky130_fd_sc_hd__o22a_1 _08457_ (.A1(net287),
    .A2(net111),
    .B1(net109),
    .B2(net237),
    .X(_01549_));
 sky130_fd_sc_hd__xnor2_1 _08458_ (.A(_06494_),
    .B(_01549_),
    .Y(_01550_));
 sky130_fd_sc_hd__or2_1 _08459_ (.A(_01548_),
    .B(_01550_),
    .X(_01551_));
 sky130_fd_sc_hd__xnor2_1 _08460_ (.A(_01544_),
    .B(_01546_),
    .Y(_01552_));
 sky130_fd_sc_hd__o32a_1 _08461_ (.A1(_01548_),
    .A2(_01550_),
    .A3(_01552_),
    .B1(_01546_),
    .B2(_01544_),
    .X(_01553_));
 sky130_fd_sc_hd__xnor2_1 _08462_ (.A(_01540_),
    .B(_01542_),
    .Y(_01554_));
 sky130_fd_sc_hd__nand2b_1 _08463_ (.A_N(_01553_),
    .B(_01554_),
    .Y(_01555_));
 sky130_fd_sc_hd__nand2_1 _08464_ (.A(_01543_),
    .B(_01555_),
    .Y(_01556_));
 sky130_fd_sc_hd__xor2_2 _08465_ (.A(_01529_),
    .B(_01530_),
    .X(_01557_));
 sky130_fd_sc_hd__nand2_1 _08466_ (.A(_01556_),
    .B(_01557_),
    .Y(_01558_));
 sky130_fd_sc_hd__and3_1 _08467_ (.A(_01527_),
    .B(_01531_),
    .C(_01558_),
    .X(_01559_));
 sky130_fd_sc_hd__xnor2_2 _08468_ (.A(_01515_),
    .B(_01517_),
    .Y(_01560_));
 sky130_fd_sc_hd__xnor2_1 _08469_ (.A(_01553_),
    .B(_01554_),
    .Y(_01561_));
 sky130_fd_sc_hd__xnor2_1 _08470_ (.A(_01560_),
    .B(_01561_),
    .Y(_01562_));
 sky130_fd_sc_hd__xor2_1 _08471_ (.A(_01538_),
    .B(_01539_),
    .X(_01563_));
 sky130_fd_sc_hd__o22a_1 _08472_ (.A1(net131),
    .A2(net143),
    .B1(net140),
    .B2(net133),
    .X(_01564_));
 sky130_fd_sc_hd__xnor2_2 _08473_ (.A(net180),
    .B(_01564_),
    .Y(_01565_));
 sky130_fd_sc_hd__o22a_1 _08474_ (.A1(net153),
    .A2(net129),
    .B1(net108),
    .B2(net155),
    .X(_01566_));
 sky130_fd_sc_hd__xnor2_2 _08475_ (.A(net208),
    .B(_01566_),
    .Y(_01567_));
 sky130_fd_sc_hd__or2_1 _08476_ (.A(_01565_),
    .B(_01567_),
    .X(_01568_));
 sky130_fd_sc_hd__o22a_1 _08477_ (.A1(net147),
    .A2(net127),
    .B1(net141),
    .B2(net145),
    .X(_01569_));
 sky130_fd_sc_hd__xor2_2 _08478_ (.A(net201),
    .B(_01569_),
    .X(_01570_));
 sky130_fd_sc_hd__inv_2 _08479_ (.A(_01570_),
    .Y(_01571_));
 sky130_fd_sc_hd__xnor2_2 _08480_ (.A(_01565_),
    .B(_01567_),
    .Y(_01572_));
 sky130_fd_sc_hd__o21a_1 _08481_ (.A1(_01571_),
    .A2(_01572_),
    .B1(_01568_),
    .X(_01573_));
 sky130_fd_sc_hd__nand2b_1 _08482_ (.A_N(_01573_),
    .B(_01563_),
    .Y(_01574_));
 sky130_fd_sc_hd__xnor2_1 _08483_ (.A(_01563_),
    .B(_01573_),
    .Y(_01575_));
 sky130_fd_sc_hd__or2_1 _08484_ (.A(net215),
    .B(net107),
    .X(_01576_));
 sky130_fd_sc_hd__xor2_1 _08485_ (.A(_01548_),
    .B(_01550_),
    .X(_01577_));
 sky130_fd_sc_hd__nor2_1 _08486_ (.A(_01576_),
    .B(_01577_),
    .Y(_01578_));
 sky130_fd_sc_hd__a21oi_1 _08487_ (.A1(net136),
    .A2(_01576_),
    .B1(_01578_),
    .Y(_01579_));
 sky130_fd_sc_hd__a21bo_1 _08488_ (.A1(_01575_),
    .A2(_01579_),
    .B1_N(_01574_),
    .X(_01580_));
 sky130_fd_sc_hd__nand2b_1 _08489_ (.A_N(_01562_),
    .B(_01580_),
    .Y(_01581_));
 sky130_fd_sc_hd__a21bo_1 _08490_ (.A1(_01560_),
    .A2(_01561_),
    .B1_N(_01581_),
    .X(_01582_));
 sky130_fd_sc_hd__xor2_2 _08491_ (.A(_01556_),
    .B(_01557_),
    .X(_01583_));
 sky130_fd_sc_hd__and2_1 _08492_ (.A(_01582_),
    .B(_01583_),
    .X(_01584_));
 sky130_fd_sc_hd__a21oi_2 _08493_ (.A1(_01531_),
    .A2(_01558_),
    .B1(_01527_),
    .Y(_01585_));
 sky130_fd_sc_hd__or2_1 _08494_ (.A(_01582_),
    .B(_01583_),
    .X(_01586_));
 sky130_fd_sc_hd__xor2_1 _08495_ (.A(_01582_),
    .B(_01583_),
    .X(_01587_));
 sky130_fd_sc_hd__xor2_1 _08496_ (.A(_01562_),
    .B(_01580_),
    .X(_01588_));
 sky130_fd_sc_hd__xnor2_1 _08497_ (.A(_01551_),
    .B(_01552_),
    .Y(_01589_));
 sky130_fd_sc_hd__xnor2_1 _08498_ (.A(_01575_),
    .B(_01579_),
    .Y(_01590_));
 sky130_fd_sc_hd__or2_1 _08499_ (.A(_01589_),
    .B(_01590_),
    .X(_01591_));
 sky130_fd_sc_hd__xnor2_1 _08500_ (.A(_01589_),
    .B(_01590_),
    .Y(_01592_));
 sky130_fd_sc_hd__o22a_1 _08501_ (.A1(net237),
    .A2(net115),
    .B1(net109),
    .B2(net287),
    .X(_01593_));
 sky130_fd_sc_hd__xnor2_1 _08502_ (.A(_06494_),
    .B(_01593_),
    .Y(_01594_));
 sky130_fd_sc_hd__o22a_1 _08503_ (.A1(net155),
    .A2(net129),
    .B1(net127),
    .B2(net153),
    .X(_01595_));
 sky130_fd_sc_hd__xnor2_1 _08504_ (.A(net208),
    .B(_01595_),
    .Y(_01596_));
 sky130_fd_sc_hd__or2_1 _08505_ (.A(_01594_),
    .B(_01596_),
    .X(_01597_));
 sky130_fd_sc_hd__xnor2_1 _08506_ (.A(_01594_),
    .B(_01596_),
    .Y(_01598_));
 sky130_fd_sc_hd__a22o_1 _08507_ (.A1(_06557_),
    .A2(net113),
    .B1(_00374_),
    .B2(_06565_),
    .X(_01599_));
 sky130_fd_sc_hd__xnor2_2 _08508_ (.A(_06534_),
    .B(_01599_),
    .Y(_01600_));
 sky130_fd_sc_hd__inv_2 _08509_ (.A(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__o21a_1 _08510_ (.A1(_01598_),
    .A2(_01601_),
    .B1(_01597_),
    .X(_01602_));
 sky130_fd_sc_hd__xnor2_2 _08511_ (.A(_01570_),
    .B(_01572_),
    .Y(_01603_));
 sky130_fd_sc_hd__nand2b_1 _08512_ (.A_N(_01602_),
    .B(_01603_),
    .Y(_01604_));
 sky130_fd_sc_hd__o22a_1 _08513_ (.A1(net147),
    .A2(net141),
    .B1(net140),
    .B2(net145),
    .X(_01605_));
 sky130_fd_sc_hd__xnor2_1 _08514_ (.A(net203),
    .B(_01605_),
    .Y(_01606_));
 sky130_fd_sc_hd__o22a_1 _08515_ (.A1(net215),
    .A2(net131),
    .B1(net143),
    .B2(net134),
    .X(_01607_));
 sky130_fd_sc_hd__xnor2_1 _08516_ (.A(net180),
    .B(_01607_),
    .Y(_01608_));
 sky130_fd_sc_hd__nor2_1 _08517_ (.A(_01606_),
    .B(_01608_),
    .Y(_01609_));
 sky130_fd_sc_hd__xnor2_2 _08518_ (.A(_01602_),
    .B(_01603_),
    .Y(_01610_));
 sky130_fd_sc_hd__a21bo_1 _08519_ (.A1(_01609_),
    .A2(_01610_),
    .B1_N(_01604_),
    .X(_01611_));
 sky130_fd_sc_hd__nand2b_1 _08520_ (.A_N(_01592_),
    .B(_01611_),
    .Y(_01612_));
 sky130_fd_sc_hd__and3_1 _08521_ (.A(_01588_),
    .B(_01591_),
    .C(_01612_),
    .X(_01613_));
 sky130_fd_sc_hd__xnor2_1 _08522_ (.A(_01592_),
    .B(_01611_),
    .Y(_01614_));
 sky130_fd_sc_hd__xnor2_2 _08523_ (.A(_01609_),
    .B(_01610_),
    .Y(_01615_));
 sky130_fd_sc_hd__and2_1 _08524_ (.A(_01576_),
    .B(_01577_),
    .X(_01616_));
 sky130_fd_sc_hd__nor2_1 _08525_ (.A(_01578_),
    .B(_01616_),
    .Y(_01617_));
 sky130_fd_sc_hd__nor2_1 _08526_ (.A(_01615_),
    .B(_01617_),
    .Y(_01618_));
 sky130_fd_sc_hd__xnor2_1 _08527_ (.A(_01598_),
    .B(_01600_),
    .Y(_01619_));
 sky130_fd_sc_hd__o22a_1 _08528_ (.A1(net287),
    .A2(net115),
    .B1(net114),
    .B2(net237),
    .X(_01620_));
 sky130_fd_sc_hd__xnor2_2 _08529_ (.A(net238),
    .B(_01620_),
    .Y(_01621_));
 sky130_fd_sc_hd__o22a_1 _08530_ (.A1(net155),
    .A2(net127),
    .B1(net141),
    .B2(net153),
    .X(_01622_));
 sky130_fd_sc_hd__xnor2_2 _08531_ (.A(net208),
    .B(_01622_),
    .Y(_01623_));
 sky130_fd_sc_hd__or2_1 _08532_ (.A(_01621_),
    .B(_01623_),
    .X(_01624_));
 sky130_fd_sc_hd__o22a_1 _08533_ (.A1(net149),
    .A2(net129),
    .B1(net108),
    .B2(net151),
    .X(_01625_));
 sky130_fd_sc_hd__xnor2_2 _08534_ (.A(net204),
    .B(_01625_),
    .Y(_01626_));
 sky130_fd_sc_hd__xnor2_2 _08535_ (.A(_01621_),
    .B(_01623_),
    .Y(_01627_));
 sky130_fd_sc_hd__o21a_1 _08536_ (.A1(_01626_),
    .A2(_01627_),
    .B1(_01624_),
    .X(_01628_));
 sky130_fd_sc_hd__nand2b_1 _08537_ (.A_N(_01628_),
    .B(_01619_),
    .Y(_01629_));
 sky130_fd_sc_hd__o22a_1 _08538_ (.A1(net145),
    .A2(net143),
    .B1(net140),
    .B2(net147),
    .X(_01630_));
 sky130_fd_sc_hd__xnor2_2 _08539_ (.A(net201),
    .B(_01630_),
    .Y(_01631_));
 sky130_fd_sc_hd__nor2_1 _08540_ (.A(net215),
    .B(net133),
    .Y(_01632_));
 sky130_fd_sc_hd__xnor2_1 _08541_ (.A(net180),
    .B(_01632_),
    .Y(_01633_));
 sky130_fd_sc_hd__and2b_1 _08542_ (.A_N(_01631_),
    .B(_01633_),
    .X(_01634_));
 sky130_fd_sc_hd__xnor2_1 _08543_ (.A(_01619_),
    .B(_01628_),
    .Y(_01635_));
 sky130_fd_sc_hd__a21bo_1 _08544_ (.A1(_01634_),
    .A2(_01635_),
    .B1_N(_01629_),
    .X(_01636_));
 sky130_fd_sc_hd__xnor2_2 _08545_ (.A(_01615_),
    .B(_01617_),
    .Y(_01637_));
 sky130_fd_sc_hd__and2b_1 _08546_ (.A_N(_01637_),
    .B(_01636_),
    .X(_01638_));
 sky130_fd_sc_hd__o21ai_1 _08547_ (.A1(_01618_),
    .A2(_01638_),
    .B1(_01614_),
    .Y(_01639_));
 sky130_fd_sc_hd__a21oi_1 _08548_ (.A1(_01591_),
    .A2(_01612_),
    .B1(_01588_),
    .Y(_01640_));
 sky130_fd_sc_hd__a21o_1 _08549_ (.A1(_01591_),
    .A2(_01612_),
    .B1(_01588_),
    .X(_01641_));
 sky130_fd_sc_hd__or3_2 _08550_ (.A(_01614_),
    .B(_01618_),
    .C(_01638_),
    .X(_01642_));
 sky130_fd_sc_hd__and2_1 _08551_ (.A(_01639_),
    .B(_01642_),
    .X(_01643_));
 sky130_fd_sc_hd__and2_1 _08552_ (.A(_01606_),
    .B(_01608_),
    .X(_01644_));
 sky130_fd_sc_hd__or2_1 _08553_ (.A(_01609_),
    .B(_01644_),
    .X(_01645_));
 sky130_fd_sc_hd__xnor2_1 _08554_ (.A(_01634_),
    .B(_01635_),
    .Y(_01646_));
 sky130_fd_sc_hd__or2_1 _08555_ (.A(_01645_),
    .B(_01646_),
    .X(_01647_));
 sky130_fd_sc_hd__xor2_1 _08556_ (.A(_01645_),
    .B(_01646_),
    .X(_01648_));
 sky130_fd_sc_hd__xor2_2 _08557_ (.A(_01626_),
    .B(_01627_),
    .X(_01649_));
 sky130_fd_sc_hd__and2b_1 _08558_ (.A_N(net180),
    .B(_01649_),
    .X(_01650_));
 sky130_fd_sc_hd__o22a_1 _08559_ (.A1(net287),
    .A2(net114),
    .B1(net108),
    .B2(net237),
    .X(_01651_));
 sky130_fd_sc_hd__xnor2_1 _08560_ (.A(net238),
    .B(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__o22a_1 _08561_ (.A1(net151),
    .A2(net129),
    .B1(net127),
    .B2(net149),
    .X(_01653_));
 sky130_fd_sc_hd__xnor2_1 _08562_ (.A(net204),
    .B(_01653_),
    .Y(_01654_));
 sky130_fd_sc_hd__nor2_2 _08563_ (.A(_01652_),
    .B(_01654_),
    .Y(_01655_));
 sky130_fd_sc_hd__xnor2_2 _08564_ (.A(net180),
    .B(_01649_),
    .Y(_01656_));
 sky130_fd_sc_hd__a21o_1 _08565_ (.A1(_01655_),
    .A2(_01656_),
    .B1(_01650_),
    .X(_01657_));
 sky130_fd_sc_hd__nand2_1 _08566_ (.A(_01648_),
    .B(_01657_),
    .Y(_01658_));
 sky130_fd_sc_hd__xor2_2 _08567_ (.A(_01636_),
    .B(_01637_),
    .X(_01659_));
 sky130_fd_sc_hd__nand3_2 _08568_ (.A(_01647_),
    .B(_01658_),
    .C(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__xnor2_2 _08569_ (.A(_01631_),
    .B(_01633_),
    .Y(_01661_));
 sky130_fd_sc_hd__xor2_2 _08570_ (.A(_01655_),
    .B(_01656_),
    .X(_01662_));
 sky130_fd_sc_hd__nand2_1 _08571_ (.A(_01661_),
    .B(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__a22o_1 _08572_ (.A1(_06519_),
    .A2(_00213_),
    .B1(_00374_),
    .B2(net292),
    .X(_01664_));
 sky130_fd_sc_hd__xnor2_2 _08573_ (.A(net238),
    .B(_01664_),
    .Y(_01665_));
 sky130_fd_sc_hd__a22o_1 _08574_ (.A1(_06557_),
    .A2(_00226_),
    .B1(_00258_),
    .B2(_06565_),
    .X(_01666_));
 sky130_fd_sc_hd__xnor2_2 _08575_ (.A(net204),
    .B(_01666_),
    .Y(_01667_));
 sky130_fd_sc_hd__o22a_1 _08576_ (.A1(net155),
    .A2(net141),
    .B1(net140),
    .B2(net153),
    .X(_01668_));
 sky130_fd_sc_hd__xnor2_1 _08577_ (.A(_06532_),
    .B(_01668_),
    .Y(_01669_));
 sky130_fd_sc_hd__nand3_2 _08578_ (.A(_01665_),
    .B(_01667_),
    .C(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__o22a_1 _08579_ (.A1(net216),
    .A2(net146),
    .B1(net144),
    .B2(net148),
    .X(_01671_));
 sky130_fd_sc_hd__xor2_1 _08580_ (.A(net201),
    .B(_01671_),
    .X(_01672_));
 sky130_fd_sc_hd__a21o_1 _08581_ (.A1(_01665_),
    .A2(_01667_),
    .B1(_01669_),
    .X(_01673_));
 sky130_fd_sc_hd__nand3_2 _08582_ (.A(_01670_),
    .B(_01672_),
    .C(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__nand2_2 _08583_ (.A(_01670_),
    .B(_01674_),
    .Y(_01675_));
 sky130_fd_sc_hd__inv_2 _08584_ (.A(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__xnor2_2 _08585_ (.A(_01661_),
    .B(_01662_),
    .Y(_01677_));
 sky130_fd_sc_hd__o21ai_1 _08586_ (.A1(_01676_),
    .A2(_01677_),
    .B1(_01663_),
    .Y(_01678_));
 sky130_fd_sc_hd__xor2_1 _08587_ (.A(_01648_),
    .B(_01657_),
    .X(_01679_));
 sky130_fd_sc_hd__and2_1 _08588_ (.A(_01678_),
    .B(_01679_),
    .X(_01680_));
 sky130_fd_sc_hd__a21oi_1 _08589_ (.A1(_01647_),
    .A2(_01658_),
    .B1(_01659_),
    .Y(_01681_));
 sky130_fd_sc_hd__a21o_1 _08590_ (.A1(_01647_),
    .A2(_01658_),
    .B1(_01659_),
    .X(_01682_));
 sky130_fd_sc_hd__or2_1 _08591_ (.A(_01678_),
    .B(_01679_),
    .X(_01683_));
 sky130_fd_sc_hd__xor2_1 _08592_ (.A(_01678_),
    .B(_01679_),
    .X(_01684_));
 sky130_fd_sc_hd__and2_1 _08593_ (.A(_01652_),
    .B(_01654_),
    .X(_01685_));
 sky130_fd_sc_hd__nor2_1 _08594_ (.A(_01655_),
    .B(_01685_),
    .Y(_01686_));
 sky130_fd_sc_hd__a21o_1 _08595_ (.A1(_01670_),
    .A2(_01673_),
    .B1(_01672_),
    .X(_01687_));
 sky130_fd_sc_hd__nand3_1 _08596_ (.A(_01674_),
    .B(_01686_),
    .C(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__a21o_1 _08597_ (.A1(_01674_),
    .A2(_01687_),
    .B1(_01686_),
    .X(_01689_));
 sky130_fd_sc_hd__nor2_1 _08598_ (.A(net215),
    .B(net147),
    .Y(_01690_));
 sky130_fd_sc_hd__o22a_1 _08599_ (.A1(net153),
    .A2(net143),
    .B1(net140),
    .B2(net155),
    .X(_01691_));
 sky130_fd_sc_hd__xnor2_1 _08600_ (.A(net208),
    .B(_01691_),
    .Y(_01692_));
 sky130_fd_sc_hd__nand2_1 _08601_ (.A(_01690_),
    .B(_01692_),
    .Y(_01693_));
 sky130_fd_sc_hd__o21ai_1 _08602_ (.A1(net216),
    .A2(net147),
    .B1(net201),
    .Y(_01694_));
 sky130_fd_sc_hd__and4_1 _08603_ (.A(_01688_),
    .B(_01689_),
    .C(_01693_),
    .D(_01694_),
    .X(_01695_));
 sky130_fd_sc_hd__a31o_1 _08604_ (.A1(_01674_),
    .A2(_01686_),
    .A3(_01687_),
    .B1(_01695_),
    .X(_01696_));
 sky130_fd_sc_hd__xnor2_2 _08605_ (.A(_01675_),
    .B(_01677_),
    .Y(_01697_));
 sky130_fd_sc_hd__or2_1 _08606_ (.A(_01696_),
    .B(_01697_),
    .X(_01698_));
 sky130_fd_sc_hd__and2_1 _08607_ (.A(_01696_),
    .B(_01697_),
    .X(_01699_));
 sky130_fd_sc_hd__xor2_1 _08608_ (.A(_01665_),
    .B(_01667_),
    .X(_01700_));
 sky130_fd_sc_hd__or2_1 _08609_ (.A(_01690_),
    .B(_01692_),
    .X(_01701_));
 sky130_fd_sc_hd__nand2_1 _08610_ (.A(_01693_),
    .B(_01701_),
    .Y(_01702_));
 sky130_fd_sc_hd__nand2_1 _08611_ (.A(_01700_),
    .B(_01702_),
    .Y(_01703_));
 sky130_fd_sc_hd__a21o_1 _08612_ (.A1(_00210_),
    .A2(_00211_),
    .B1(net287),
    .X(_01704_));
 sky130_fd_sc_hd__or3_1 _08613_ (.A(net237),
    .B(_00224_),
    .C(_00225_),
    .X(_01705_));
 sky130_fd_sc_hd__a21o_1 _08614_ (.A1(_01704_),
    .A2(_01705_),
    .B1(net239),
    .X(_01706_));
 sky130_fd_sc_hd__nand3_1 _08615_ (.A(net239),
    .B(_01704_),
    .C(_01705_),
    .Y(_01707_));
 sky130_fd_sc_hd__a22o_1 _08616_ (.A1(_06557_),
    .A2(_00258_),
    .B1(_00265_),
    .B2(_06565_),
    .X(_01708_));
 sky130_fd_sc_hd__xnor2_1 _08617_ (.A(net205),
    .B(_01708_),
    .Y(_01709_));
 sky130_fd_sc_hd__and3_2 _08618_ (.A(_01706_),
    .B(_01707_),
    .C(_01709_),
    .X(_01710_));
 sky130_fd_sc_hd__xor2_1 _08619_ (.A(_01700_),
    .B(_01702_),
    .X(_01711_));
 sky130_fd_sc_hd__nand2_1 _08620_ (.A(_01710_),
    .B(_01711_),
    .Y(_01712_));
 sky130_fd_sc_hd__a22oi_2 _08621_ (.A1(_01688_),
    .A2(_01689_),
    .B1(_01693_),
    .B2(_01694_),
    .Y(_01713_));
 sky130_fd_sc_hd__a211oi_1 _08622_ (.A1(_01703_),
    .A2(_01712_),
    .B1(_01713_),
    .C1(_01695_),
    .Y(_01714_));
 sky130_fd_sc_hd__o211a_1 _08623_ (.A1(_01695_),
    .A2(_01713_),
    .B1(_01712_),
    .C1(_01703_),
    .X(_01715_));
 sky130_fd_sc_hd__nor2_1 _08624_ (.A(_01714_),
    .B(_01715_),
    .Y(_01716_));
 sky130_fd_sc_hd__xnor2_1 _08625_ (.A(_01710_),
    .B(_01711_),
    .Y(_01717_));
 sky130_fd_sc_hd__a21oi_2 _08626_ (.A1(_01706_),
    .A2(_01707_),
    .B1(_01709_),
    .Y(_01718_));
 sky130_fd_sc_hd__o22a_1 _08627_ (.A1(net215),
    .A2(net153),
    .B1(net143),
    .B2(net155),
    .X(_01719_));
 sky130_fd_sc_hd__xnor2_1 _08628_ (.A(_06532_),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__nor3b_1 _08629_ (.A(_01710_),
    .B(_01718_),
    .C_N(_01720_),
    .Y(_01721_));
 sky130_fd_sc_hd__or3b_1 _08630_ (.A(_01710_),
    .B(_01718_),
    .C_N(_01720_),
    .X(_01722_));
 sky130_fd_sc_hd__a22o_1 _08631_ (.A1(_06565_),
    .A2(_00240_),
    .B1(_00265_),
    .B2(_06557_),
    .X(_01723_));
 sky130_fd_sc_hd__xor2_2 _08632_ (.A(net205),
    .B(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__o32ai_4 _08633_ (.A1(net287),
    .A2(_00224_),
    .A3(_00225_),
    .B1(net142),
    .B2(_06520_),
    .Y(_01725_));
 sky130_fd_sc_hd__xnor2_2 _08634_ (.A(net240),
    .B(_01725_),
    .Y(_01726_));
 sky130_fd_sc_hd__or2_1 _08635_ (.A(_01724_),
    .B(_01726_),
    .X(_01727_));
 sky130_fd_sc_hd__o21ba_1 _08636_ (.A1(_01710_),
    .A2(_01718_),
    .B1_N(_01720_),
    .X(_01728_));
 sky130_fd_sc_hd__or3_2 _08637_ (.A(_01721_),
    .B(_01727_),
    .C(_01728_),
    .X(_01729_));
 sky130_fd_sc_hd__and3_1 _08638_ (.A(_01717_),
    .B(_01722_),
    .C(_01729_),
    .X(_01730_));
 sky130_fd_sc_hd__a21oi_1 _08639_ (.A1(_01722_),
    .A2(_01729_),
    .B1(_01717_),
    .Y(_01731_));
 sky130_fd_sc_hd__xor2_2 _08640_ (.A(_01724_),
    .B(_01726_),
    .X(_01732_));
 sky130_fd_sc_hd__nor2_1 _08641_ (.A(net216),
    .B(net155),
    .Y(_01733_));
 sky130_fd_sc_hd__mux2_1 _08642_ (.A0(_06532_),
    .A1(_01732_),
    .S(_01733_),
    .X(_01734_));
 sky130_fd_sc_hd__o21ai_1 _08643_ (.A1(_01721_),
    .A2(_01728_),
    .B1(_01727_),
    .Y(_01735_));
 sky130_fd_sc_hd__a21oi_1 _08644_ (.A1(_01729_),
    .A2(_01735_),
    .B1(_01734_),
    .Y(_01736_));
 sky130_fd_sc_hd__a21o_1 _08645_ (.A1(_01729_),
    .A2(_01735_),
    .B1(_01734_),
    .X(_01737_));
 sky130_fd_sc_hd__and3_1 _08646_ (.A(_01729_),
    .B(_01734_),
    .C(_01735_),
    .X(_01738_));
 sky130_fd_sc_hd__a22o_1 _08647_ (.A1(net292),
    .A2(_00258_),
    .B1(_00265_),
    .B2(_06519_),
    .X(_01739_));
 sky130_fd_sc_hd__xnor2_1 _08648_ (.A(net240),
    .B(_01739_),
    .Y(_01740_));
 sky130_fd_sc_hd__o22a_1 _08649_ (.A1(net215),
    .A2(net149),
    .B1(net143),
    .B2(net151),
    .X(_01741_));
 sky130_fd_sc_hd__xnor2_1 _08650_ (.A(_06534_),
    .B(_01741_),
    .Y(_01742_));
 sky130_fd_sc_hd__nor2_1 _08651_ (.A(_01740_),
    .B(_01742_),
    .Y(_01743_));
 sky130_fd_sc_hd__xnor2_2 _08652_ (.A(_01732_),
    .B(_01733_),
    .Y(_01744_));
 sky130_fd_sc_hd__and2b_1 _08653_ (.A_N(_01744_),
    .B(_01743_),
    .X(_01745_));
 sky130_fd_sc_hd__xnor2_2 _08654_ (.A(_01743_),
    .B(_01744_),
    .Y(_01746_));
 sky130_fd_sc_hd__a22o_1 _08655_ (.A1(_06519_),
    .A2(_00240_),
    .B1(_00265_),
    .B2(net293),
    .X(_01747_));
 sky130_fd_sc_hd__xnor2_2 _08656_ (.A(net240),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__nor2_1 _08657_ (.A(net216),
    .B(net151),
    .Y(_01749_));
 sky130_fd_sc_hd__xnor2_1 _08658_ (.A(_06534_),
    .B(_01749_),
    .Y(_01750_));
 sky130_fd_sc_hd__and2b_1 _08659_ (.A_N(_01748_),
    .B(_01750_),
    .X(_01751_));
 sky130_fd_sc_hd__and2b_1 _08660_ (.A_N(_01750_),
    .B(_01748_),
    .X(_01752_));
 sky130_fd_sc_hd__xor2_1 _08661_ (.A(_01748_),
    .B(_01749_),
    .X(_01753_));
 sky130_fd_sc_hd__a22o_1 _08662_ (.A1(net214),
    .A2(_06519_),
    .B1(_00240_),
    .B2(net292),
    .X(_01754_));
 sky130_fd_sc_hd__or2_1 _08663_ (.A(_06441_),
    .B(_01754_),
    .X(_01755_));
 sky130_fd_sc_hd__or3_1 _08664_ (.A(net238),
    .B(_01753_),
    .C(_01755_),
    .X(_01756_));
 sky130_fd_sc_hd__xor2_1 _08665_ (.A(_01740_),
    .B(_01742_),
    .X(_01757_));
 sky130_fd_sc_hd__xnor2_1 _08666_ (.A(_01751_),
    .B(_01757_),
    .Y(_01758_));
 sky130_fd_sc_hd__mux2_1 _08667_ (.A0(_06534_),
    .A1(_01748_),
    .S(_01749_),
    .X(_01759_));
 sky130_fd_sc_hd__inv_2 _08668_ (.A(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__a2bb2o_1 _08669_ (.A1_N(_01756_),
    .A2_N(_01758_),
    .B1(_01760_),
    .B2(_01757_),
    .X(_01761_));
 sky130_fd_sc_hd__a21o_1 _08670_ (.A1(_01746_),
    .A2(_01761_),
    .B1(_01745_),
    .X(_01762_));
 sky130_fd_sc_hd__nor2_1 _08671_ (.A(_01736_),
    .B(_01738_),
    .Y(_01763_));
 sky130_fd_sc_hd__a21o_1 _08672_ (.A1(_01737_),
    .A2(_01762_),
    .B1(_01738_),
    .X(_01764_));
 sky130_fd_sc_hd__o21ba_1 _08673_ (.A1(_01731_),
    .A2(_01764_),
    .B1_N(_01730_),
    .X(_01765_));
 sky130_fd_sc_hd__or2_1 _08674_ (.A(_01730_),
    .B(_01731_),
    .X(_01766_));
 sky130_fd_sc_hd__o21ba_1 _08675_ (.A1(_01714_),
    .A2(_01765_),
    .B1_N(_01715_),
    .X(_01767_));
 sky130_fd_sc_hd__a21o_1 _08676_ (.A1(_01696_),
    .A2(_01697_),
    .B1(_01767_),
    .X(_01768_));
 sky130_fd_sc_hd__xor2_2 _08677_ (.A(_01696_),
    .B(_01697_),
    .X(_01769_));
 sky130_fd_sc_hd__and3_1 _08678_ (.A(_01684_),
    .B(_01698_),
    .C(_01768_),
    .X(_01770_));
 sky130_fd_sc_hd__a311o_1 _08679_ (.A1(_01684_),
    .A2(_01698_),
    .A3(_01768_),
    .B1(_01681_),
    .C1(_01680_),
    .X(_01771_));
 sky130_fd_sc_hd__and2_1 _08680_ (.A(_01660_),
    .B(_01682_),
    .X(_01772_));
 sky130_fd_sc_hd__nand3_1 _08681_ (.A(_01643_),
    .B(_01660_),
    .C(_01771_),
    .Y(_01773_));
 sky130_fd_sc_hd__a21oi_1 _08682_ (.A1(_01639_),
    .A2(_01641_),
    .B1(_01613_),
    .Y(_01774_));
 sky130_fd_sc_hd__nor2_1 _08683_ (.A(_01613_),
    .B(_01640_),
    .Y(_01775_));
 sky130_fd_sc_hd__a41o_1 _08684_ (.A1(_01643_),
    .A2(_01660_),
    .A3(_01771_),
    .A4(_01775_),
    .B1(_01774_),
    .X(_01776_));
 sky130_fd_sc_hd__a211oi_1 _08685_ (.A1(_01587_),
    .A2(_01776_),
    .B1(_01584_),
    .C1(_01585_),
    .Y(_01777_));
 sky130_fd_sc_hd__or2_1 _08686_ (.A(_01559_),
    .B(_01585_),
    .X(_01778_));
 sky130_fd_sc_hd__or3_2 _08687_ (.A(_01526_),
    .B(_01559_),
    .C(_01777_),
    .X(_01779_));
 sky130_fd_sc_hd__a31o_2 _08688_ (.A1(_01496_),
    .A2(_01524_),
    .A3(_01779_),
    .B1(_01495_),
    .X(_01780_));
 sky130_fd_sc_hd__xnor2_4 _08689_ (.A(_01374_),
    .B(_01416_),
    .Y(_01781_));
 sky130_fd_sc_hd__and3_1 _08690_ (.A(_01421_),
    .B(_01451_),
    .C(_01452_),
    .X(_01782_));
 sky130_fd_sc_hd__or2_2 _08691_ (.A(_01453_),
    .B(_01782_),
    .X(_01783_));
 sky130_fd_sc_hd__o31ai_2 _08692_ (.A1(_01780_),
    .A2(_01781_),
    .A3(_01783_),
    .B1(_01455_),
    .Y(_01784_));
 sky130_fd_sc_hd__or4_1 _08693_ (.A(_01370_),
    .B(_01372_),
    .C(_01781_),
    .D(_01783_),
    .X(_01785_));
 sky130_fd_sc_hd__o221a_2 _08694_ (.A1(_01373_),
    .A2(_01455_),
    .B1(_01780_),
    .B2(_01785_),
    .C1(_01369_),
    .X(_01786_));
 sky130_fd_sc_hd__a22o_1 _08695_ (.A1(_01102_),
    .A2(_01103_),
    .B1(_01166_),
    .B2(_01167_),
    .X(_01787_));
 sky130_fd_sc_hd__o21ai_1 _08696_ (.A1(_01102_),
    .A2(_01103_),
    .B1(_01787_),
    .Y(_01788_));
 sky130_fd_sc_hd__a21o_1 _08697_ (.A1(_01268_),
    .A2(_01272_),
    .B1(_01273_),
    .X(_01789_));
 sky130_fd_sc_hd__a2111o_1 _08698_ (.A1(_01268_),
    .A2(_01272_),
    .B1(_01273_),
    .C1(_01168_),
    .D1(_01105_),
    .X(_01790_));
 sky130_fd_sc_hd__o311a_2 _08699_ (.A1(_01169_),
    .A2(_01275_),
    .A3(_01786_),
    .B1(_01788_),
    .C1(_01790_),
    .X(_01791_));
 sky130_fd_sc_hd__a21o_1 _08700_ (.A1(_00913_),
    .A2(_00967_),
    .B1(_00968_),
    .X(_01792_));
 sky130_fd_sc_hd__a21o_1 _08701_ (.A1(_01041_),
    .A2(_01792_),
    .B1(_00969_),
    .X(_01793_));
 sky130_fd_sc_hd__nand2b_2 _08702_ (.A_N(_00969_),
    .B(_01792_),
    .Y(_01794_));
 sky130_fd_sc_hd__o31ai_4 _08703_ (.A1(_01042_),
    .A2(_01791_),
    .A3(_01794_),
    .B1(_01793_),
    .Y(_01795_));
 sky130_fd_sc_hd__nor2_1 _08704_ (.A(_00907_),
    .B(_00908_),
    .Y(_01796_));
 sky130_fd_sc_hd__xor2_2 _08705_ (.A(_00907_),
    .B(_00908_),
    .X(_01797_));
 sky130_fd_sc_hd__xnor2_1 _08706_ (.A(_00907_),
    .B(_00908_),
    .Y(_01798_));
 sky130_fd_sc_hd__xor2_1 _08707_ (.A(_00769_),
    .B(_00838_),
    .X(_01799_));
 sky130_fd_sc_hd__xnor2_1 _08708_ (.A(_00769_),
    .B(_00838_),
    .Y(_01800_));
 sky130_fd_sc_hd__a32o_2 _08709_ (.A1(_01795_),
    .A2(_01797_),
    .A3(_01799_),
    .B1(_00910_),
    .B2(_00839_),
    .X(_01801_));
 sky130_fd_sc_hd__xor2_2 _08710_ (.A(_00768_),
    .B(_01801_),
    .X(_01802_));
 sky130_fd_sc_hd__xnor2_2 _08711_ (.A(_01042_),
    .B(_01791_),
    .Y(_01803_));
 sky130_fd_sc_hd__inv_2 _08712_ (.A(_01803_),
    .Y(_01804_));
 sky130_fd_sc_hd__o21ai_1 _08713_ (.A1(net238),
    .A2(_01755_),
    .B1(_01753_),
    .Y(_01805_));
 sky130_fd_sc_hd__and2_1 _08714_ (.A(_01756_),
    .B(_01805_),
    .X(_01806_));
 sky130_fd_sc_hd__nor2_1 _08715_ (.A(_01755_),
    .B(_01806_),
    .Y(_01807_));
 sky130_fd_sc_hd__o31ai_1 _08716_ (.A1(net204),
    .A2(_01751_),
    .A3(_01752_),
    .B1(_01756_),
    .Y(_01808_));
 sky130_fd_sc_hd__xor2_1 _08717_ (.A(_01758_),
    .B(_01808_),
    .X(_01809_));
 sky130_fd_sc_hd__nand2_1 _08718_ (.A(_01807_),
    .B(_01809_),
    .Y(_01810_));
 sky130_fd_sc_hd__xor2_2 _08719_ (.A(_01746_),
    .B(_01761_),
    .X(_01811_));
 sky130_fd_sc_hd__nor2_1 _08720_ (.A(_01810_),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__xnor2_1 _08721_ (.A(_01762_),
    .B(_01763_),
    .Y(_01813_));
 sky130_fd_sc_hd__and2_1 _08722_ (.A(_01812_),
    .B(_01813_),
    .X(_01814_));
 sky130_fd_sc_hd__xor2_1 _08723_ (.A(_01764_),
    .B(_01766_),
    .X(_01815_));
 sky130_fd_sc_hd__and2_1 _08724_ (.A(_01814_),
    .B(_01815_),
    .X(_01816_));
 sky130_fd_sc_hd__xnor2_1 _08725_ (.A(_01716_),
    .B(_01765_),
    .Y(_01817_));
 sky130_fd_sc_hd__and2_2 _08726_ (.A(_01816_),
    .B(_01817_),
    .X(_01818_));
 sky130_fd_sc_hd__xnor2_2 _08727_ (.A(_01767_),
    .B(_01769_),
    .Y(_01819_));
 sky130_fd_sc_hd__and2_1 _08728_ (.A(_01818_),
    .B(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__a21oi_2 _08729_ (.A1(_01698_),
    .A2(_01768_),
    .B1(_01684_),
    .Y(_01821_));
 sky130_fd_sc_hd__or2_1 _08730_ (.A(_01770_),
    .B(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__o211ai_4 _08731_ (.A1(_01770_),
    .A2(_01821_),
    .B1(_01819_),
    .C1(_01818_),
    .Y(_01823_));
 sky130_fd_sc_hd__a211o_1 _08732_ (.A1(_01767_),
    .A2(_01769_),
    .B1(_01680_),
    .C1(_01699_),
    .X(_01824_));
 sky130_fd_sc_hd__nand3_2 _08733_ (.A(_01683_),
    .B(_01772_),
    .C(_01824_),
    .Y(_01825_));
 sky130_fd_sc_hd__a21o_1 _08734_ (.A1(_01683_),
    .A2(_01824_),
    .B1(_01772_),
    .X(_01826_));
 sky130_fd_sc_hd__a21oi_1 _08735_ (.A1(_01825_),
    .A2(_01826_),
    .B1(_01823_),
    .Y(_01827_));
 sky130_fd_sc_hd__a21o_1 _08736_ (.A1(_01660_),
    .A2(_01771_),
    .B1(_01643_),
    .X(_01828_));
 sky130_fd_sc_hd__nand2_1 _08737_ (.A(_01773_),
    .B(_01828_),
    .Y(_01829_));
 sky130_fd_sc_hd__a221o_1 _08738_ (.A1(_01825_),
    .A2(_01826_),
    .B1(_01828_),
    .B2(_01773_),
    .C1(_01823_),
    .X(_01830_));
 sky130_fd_sc_hd__nand2_1 _08739_ (.A(_01639_),
    .B(_01682_),
    .Y(_01831_));
 sky130_fd_sc_hd__a31o_1 _08740_ (.A1(_01683_),
    .A2(_01772_),
    .A3(_01824_),
    .B1(_01831_),
    .X(_01832_));
 sky130_fd_sc_hd__nand3_1 _08741_ (.A(_01642_),
    .B(_01775_),
    .C(_01832_),
    .Y(_01833_));
 sky130_fd_sc_hd__a21o_1 _08742_ (.A1(_01642_),
    .A2(_01832_),
    .B1(_01775_),
    .X(_01834_));
 sky130_fd_sc_hd__and2_1 _08743_ (.A(_01833_),
    .B(_01834_),
    .X(_01835_));
 sky130_fd_sc_hd__or2_1 _08744_ (.A(_01830_),
    .B(_01835_),
    .X(_01836_));
 sky130_fd_sc_hd__xor2_1 _08745_ (.A(_01587_),
    .B(_01776_),
    .X(_01837_));
 sky130_fd_sc_hd__a211o_1 _08746_ (.A1(_01833_),
    .A2(_01834_),
    .B1(_01837_),
    .C1(_01830_),
    .X(_01838_));
 sky130_fd_sc_hd__a311o_1 _08747_ (.A1(_01642_),
    .A2(_01775_),
    .A3(_01832_),
    .B1(_01640_),
    .C1(_01584_),
    .X(_01839_));
 sky130_fd_sc_hd__a21oi_2 _08748_ (.A1(_01586_),
    .A2(_01839_),
    .B1(_01778_),
    .Y(_01840_));
 sky130_fd_sc_hd__and3_1 _08749_ (.A(_01586_),
    .B(_01778_),
    .C(_01839_),
    .X(_01841_));
 sky130_fd_sc_hd__nor2_1 _08750_ (.A(_01840_),
    .B(_01841_),
    .Y(_01842_));
 sky130_fd_sc_hd__or3_1 _08751_ (.A(_01838_),
    .B(_01840_),
    .C(_01841_),
    .X(_01843_));
 sky130_fd_sc_hd__o21ai_1 _08752_ (.A1(_01559_),
    .A2(_01777_),
    .B1(_01526_),
    .Y(_01844_));
 sky130_fd_sc_hd__and2_1 _08753_ (.A(_01779_),
    .B(_01844_),
    .X(_01845_));
 sky130_fd_sc_hd__a2111o_1 _08754_ (.A1(_01779_),
    .A2(_01844_),
    .B1(_01841_),
    .C1(_01840_),
    .D1(_01838_),
    .X(_01846_));
 sky130_fd_sc_hd__a21o_1 _08755_ (.A1(_01522_),
    .A2(_01523_),
    .B1(_01585_),
    .X(_01847_));
 sky130_fd_sc_hd__o21ai_2 _08756_ (.A1(_01522_),
    .A2(_01523_),
    .B1(_01847_),
    .Y(_01848_));
 sky130_fd_sc_hd__or4bb_2 _08757_ (.A(_01526_),
    .B(_01778_),
    .C_N(_01839_),
    .D_N(_01586_),
    .X(_01849_));
 sky130_fd_sc_hd__a21o_1 _08758_ (.A1(_01848_),
    .A2(_01849_),
    .B1(_01525_),
    .X(_01850_));
 sky130_fd_sc_hd__nand3_2 _08759_ (.A(_01525_),
    .B(_01848_),
    .C(_01849_),
    .Y(_01851_));
 sky130_fd_sc_hd__a21oi_1 _08760_ (.A1(_01850_),
    .A2(_01851_),
    .B1(_01846_),
    .Y(_01852_));
 sky130_fd_sc_hd__xnor2_2 _08761_ (.A(_01780_),
    .B(_01783_),
    .Y(_01853_));
 sky130_fd_sc_hd__nand2_1 _08762_ (.A(_01852_),
    .B(_01853_),
    .Y(_01854_));
 sky130_fd_sc_hd__a21o_1 _08763_ (.A1(_01454_),
    .A2(_01496_),
    .B1(_01782_),
    .X(_01855_));
 sky130_fd_sc_hd__a211o_1 _08764_ (.A1(_01848_),
    .A2(_01849_),
    .B1(_01525_),
    .C1(_01783_),
    .X(_01856_));
 sky130_fd_sc_hd__nand2_1 _08765_ (.A(_01855_),
    .B(_01856_),
    .Y(_01857_));
 sky130_fd_sc_hd__xnor2_2 _08766_ (.A(_01781_),
    .B(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__nor2_1 _08767_ (.A(_01854_),
    .B(_01858_),
    .Y(_01859_));
 sky130_fd_sc_hd__xnor2_1 _08768_ (.A(_01372_),
    .B(_01784_),
    .Y(_01860_));
 sky130_fd_sc_hd__xor2_1 _08769_ (.A(_01372_),
    .B(_01784_),
    .X(_01861_));
 sky130_fd_sc_hd__a21o_1 _08770_ (.A1(_01368_),
    .A2(_01418_),
    .B1(_01371_),
    .X(_01862_));
 sky130_fd_sc_hd__a211o_1 _08771_ (.A1(_01855_),
    .A2(_01856_),
    .B1(_01372_),
    .C1(_01781_),
    .X(_01863_));
 sky130_fd_sc_hd__nand3_1 _08772_ (.A(_01370_),
    .B(_01862_),
    .C(_01863_),
    .Y(_01864_));
 sky130_fd_sc_hd__a21o_1 _08773_ (.A1(_01862_),
    .A2(_01863_),
    .B1(_01370_),
    .X(_01865_));
 sky130_fd_sc_hd__and2_1 _08774_ (.A(_01864_),
    .B(_01865_),
    .X(_01866_));
 sky130_fd_sc_hd__a2111o_1 _08775_ (.A1(_01864_),
    .A2(_01865_),
    .B1(_01854_),
    .C1(_01858_),
    .D1(_01860_),
    .X(_01867_));
 sky130_fd_sc_hd__xor2_2 _08776_ (.A(_01269_),
    .B(_01786_),
    .X(_01868_));
 sky130_fd_sc_hd__nor2_1 _08777_ (.A(_01867_),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__a21o_1 _08778_ (.A1(_01268_),
    .A2(_01321_),
    .B1(_01267_),
    .X(_01870_));
 sky130_fd_sc_hd__or2_1 _08779_ (.A(_01269_),
    .B(_01370_),
    .X(_01871_));
 sky130_fd_sc_hd__a21o_1 _08780_ (.A1(_01862_),
    .A2(_01863_),
    .B1(_01871_),
    .X(_01872_));
 sky130_fd_sc_hd__nand3_1 _08781_ (.A(_01274_),
    .B(_01870_),
    .C(_01872_),
    .Y(_01873_));
 sky130_fd_sc_hd__a21o_1 _08782_ (.A1(_01870_),
    .A2(_01872_),
    .B1(_01274_),
    .X(_01874_));
 sky130_fd_sc_hd__nand2_1 _08783_ (.A(_01873_),
    .B(_01874_),
    .Y(_01875_));
 sky130_fd_sc_hd__nand2_1 _08784_ (.A(_01869_),
    .B(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__o21ai_1 _08785_ (.A1(_01275_),
    .A2(_01786_),
    .B1(_01789_),
    .Y(_01877_));
 sky130_fd_sc_hd__xnor2_1 _08786_ (.A(_01168_),
    .B(_01877_),
    .Y(_01878_));
 sky130_fd_sc_hd__a2111o_2 _08787_ (.A1(_01873_),
    .A2(_01874_),
    .B1(_01878_),
    .C1(_01868_),
    .D1(_01867_),
    .X(_01879_));
 sky130_fd_sc_hd__a21bo_1 _08788_ (.A1(_01166_),
    .A2(_01167_),
    .B1_N(_01272_),
    .X(_01880_));
 sky130_fd_sc_hd__o21ai_1 _08789_ (.A1(_01166_),
    .A2(_01167_),
    .B1(_01880_),
    .Y(_01881_));
 sky130_fd_sc_hd__or2_1 _08790_ (.A(_01168_),
    .B(_01274_),
    .X(_01882_));
 sky130_fd_sc_hd__or2_1 _08791_ (.A(_01870_),
    .B(_01882_),
    .X(_01883_));
 sky130_fd_sc_hd__a211o_1 _08792_ (.A1(_01862_),
    .A2(_01863_),
    .B1(_01871_),
    .C1(_01882_),
    .X(_01884_));
 sky130_fd_sc_hd__and3_1 _08793_ (.A(_01881_),
    .B(_01883_),
    .C(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__xor2_4 _08794_ (.A(_01105_),
    .B(_01885_),
    .X(_01886_));
 sky130_fd_sc_hd__nor2_1 _08795_ (.A(_01879_),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__a21o_1 _08796_ (.A1(_01041_),
    .A2(_01104_),
    .B1(_01040_),
    .X(_01888_));
 sky130_fd_sc_hd__a311o_2 _08797_ (.A1(_01881_),
    .A2(_01883_),
    .A3(_01884_),
    .B1(_01105_),
    .C1(_01042_),
    .X(_01889_));
 sky130_fd_sc_hd__a21o_1 _08798_ (.A1(_01888_),
    .A2(_01889_),
    .B1(_01794_),
    .X(_01890_));
 sky130_fd_sc_hd__nand3_1 _08799_ (.A(_01794_),
    .B(_01888_),
    .C(_01889_),
    .Y(_01891_));
 sky130_fd_sc_hd__nand2_1 _08800_ (.A(_01890_),
    .B(_01891_),
    .Y(_01892_));
 sky130_fd_sc_hd__a2111oi_2 _08801_ (.A1(_01890_),
    .A2(_01891_),
    .B1(_01804_),
    .C1(_01879_),
    .D1(_01886_),
    .Y(_01893_));
 sky130_fd_sc_hd__xnor2_2 _08802_ (.A(_01795_),
    .B(_01797_),
    .Y(_01894_));
 sky130_fd_sc_hd__and2_2 _08803_ (.A(_01893_),
    .B(_01894_),
    .X(_01895_));
 sky130_fd_sc_hd__a21o_1 _08804_ (.A1(_00909_),
    .A2(_01792_),
    .B1(_01796_),
    .X(_01896_));
 sky130_fd_sc_hd__or2_1 _08805_ (.A(_01794_),
    .B(_01798_),
    .X(_01897_));
 sky130_fd_sc_hd__a211o_1 _08806_ (.A1(_01888_),
    .A2(_01889_),
    .B1(_01794_),
    .C1(_01798_),
    .X(_01898_));
 sky130_fd_sc_hd__and3_1 _08807_ (.A(_01800_),
    .B(_01896_),
    .C(_01898_),
    .X(_01899_));
 sky130_fd_sc_hd__a21oi_1 _08808_ (.A1(_01896_),
    .A2(_01898_),
    .B1(_01800_),
    .Y(_01900_));
 sky130_fd_sc_hd__or2_1 _08809_ (.A(_01899_),
    .B(_01900_),
    .X(_01901_));
 sky130_fd_sc_hd__nand2_1 _08810_ (.A(_01895_),
    .B(_01901_),
    .Y(_01902_));
 sky130_fd_sc_hd__o21a_1 _08811_ (.A1(_01899_),
    .A2(_01900_),
    .B1(_01802_),
    .X(_01903_));
 sky130_fd_sc_hd__a21oi_4 _08812_ (.A1(_00665_),
    .A2(_00765_),
    .B1(_00764_),
    .Y(_01904_));
 sky130_fd_sc_hd__o21ai_4 _08813_ (.A1(_00759_),
    .A2(_00760_),
    .B1(_00762_),
    .Y(_01905_));
 sky130_fd_sc_hd__a21o_1 _08814_ (.A1(_00707_),
    .A2(_00719_),
    .B1(_00717_),
    .X(_01906_));
 sky130_fd_sc_hd__a21o_1 _08815_ (.A1(_00685_),
    .A2(_00690_),
    .B1(_00692_),
    .X(_01907_));
 sky130_fd_sc_hd__o22a_1 _08816_ (.A1(net48),
    .A2(_00309_),
    .B1(_00313_),
    .B2(net46),
    .X(_01908_));
 sky130_fd_sc_hd__xnor2_1 _08817_ (.A(net97),
    .B(_01908_),
    .Y(_01909_));
 sky130_fd_sc_hd__a22o_1 _08818_ (.A1(_00226_),
    .A2(net44),
    .B1(net42),
    .B2(_00258_),
    .X(_01910_));
 sky130_fd_sc_hd__xor2_1 _08819_ (.A(net94),
    .B(_01910_),
    .X(_01911_));
 sky130_fd_sc_hd__and2_1 _08820_ (.A(_01909_),
    .B(_01911_),
    .X(_01912_));
 sky130_fd_sc_hd__nor2_1 _08821_ (.A(_01909_),
    .B(_01911_),
    .Y(_01913_));
 sky130_fd_sc_hd__nor2_1 _08822_ (.A(_01912_),
    .B(_01913_),
    .Y(_01914_));
 sky130_fd_sc_hd__a22o_1 _08823_ (.A1(_00213_),
    .A2(net37),
    .B1(_00374_),
    .B2(net39),
    .X(_01915_));
 sky130_fd_sc_hd__xor2_1 _08824_ (.A(net91),
    .B(_01915_),
    .X(_01916_));
 sky130_fd_sc_hd__xor2_1 _08825_ (.A(_01914_),
    .B(_01916_),
    .X(_01917_));
 sky130_fd_sc_hd__xnor2_1 _08826_ (.A(_01907_),
    .B(_01917_),
    .Y(_01918_));
 sky130_fd_sc_hd__and2b_1 _08827_ (.A_N(_01918_),
    .B(_01906_),
    .X(_01919_));
 sky130_fd_sc_hd__and2b_1 _08828_ (.A_N(_01906_),
    .B(_01918_),
    .X(_01920_));
 sky130_fd_sc_hd__nor2_2 _08829_ (.A(_01919_),
    .B(_01920_),
    .Y(_01921_));
 sky130_fd_sc_hd__o21ai_1 _08830_ (.A1(_00709_),
    .A2(_00711_),
    .B1(_00715_),
    .Y(_01922_));
 sky130_fd_sc_hd__o21ai_2 _08831_ (.A1(_00696_),
    .A2(_00706_),
    .B1(_00705_),
    .Y(_01923_));
 sky130_fd_sc_hd__nand2_1 _08832_ (.A(_00743_),
    .B(_01923_),
    .Y(_01924_));
 sky130_fd_sc_hd__xor2_1 _08833_ (.A(_00743_),
    .B(_01923_),
    .X(_01925_));
 sky130_fd_sc_hd__xnor2_1 _08834_ (.A(_01922_),
    .B(_01925_),
    .Y(_01926_));
 sky130_fd_sc_hd__o22a_1 _08835_ (.A1(net53),
    .A2(net106),
    .B1(net104),
    .B2(net51),
    .X(_01927_));
 sky130_fd_sc_hd__xnor2_2 _08836_ (.A(net135),
    .B(_01927_),
    .Y(_01928_));
 sky130_fd_sc_hd__o22a_1 _08837_ (.A1(net59),
    .A2(net148),
    .B1(net146),
    .B2(net57),
    .X(_01929_));
 sky130_fd_sc_hd__xnor2_2 _08838_ (.A(net202),
    .B(_01929_),
    .Y(_01930_));
 sky130_fd_sc_hd__nor2_1 _08839_ (.A(_01928_),
    .B(_01930_),
    .Y(_01931_));
 sky130_fd_sc_hd__xor2_2 _08840_ (.A(_01928_),
    .B(_01930_),
    .X(_01932_));
 sky130_fd_sc_hd__o22a_1 _08841_ (.A1(net63),
    .A2(net134),
    .B1(net132),
    .B2(net61),
    .X(_01933_));
 sky130_fd_sc_hd__xnor2_1 _08842_ (.A(net181),
    .B(_01933_),
    .Y(_01934_));
 sky130_fd_sc_hd__inv_2 _08843_ (.A(_01934_),
    .Y(_01935_));
 sky130_fd_sc_hd__xnor2_1 _08844_ (.A(_01932_),
    .B(_01934_),
    .Y(_01936_));
 sky130_fd_sc_hd__o22a_1 _08845_ (.A1(net100),
    .A2(net86),
    .B1(net82),
    .B2(net98),
    .X(_01937_));
 sky130_fd_sc_hd__xnor2_1 _08846_ (.A(net137),
    .B(_01937_),
    .Y(_01938_));
 sky130_fd_sc_hd__o22a_1 _08847_ (.A1(net35),
    .A2(net77),
    .B1(net73),
    .B2(net33),
    .X(_01939_));
 sky130_fd_sc_hd__xnor2_1 _08848_ (.A(net125),
    .B(_01939_),
    .Y(_01940_));
 sky130_fd_sc_hd__and2b_1 _08849_ (.A_N(_01938_),
    .B(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__xor2_1 _08850_ (.A(_01938_),
    .B(_01940_),
    .X(_01942_));
 sky130_fd_sc_hd__o22a_1 _08851_ (.A1(net84),
    .A2(net78),
    .B1(net74),
    .B2(net80),
    .X(_01943_));
 sky130_fd_sc_hd__xnor2_1 _08852_ (.A(net121),
    .B(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__or2_1 _08853_ (.A(_01942_),
    .B(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__nand2_1 _08854_ (.A(_01942_),
    .B(_01944_),
    .Y(_01946_));
 sky130_fd_sc_hd__nand2_1 _08855_ (.A(_01945_),
    .B(_01946_),
    .Y(_01947_));
 sky130_fd_sc_hd__o22a_1 _08856_ (.A1(net150),
    .A2(net56),
    .B1(net17),
    .B2(net152),
    .X(_01948_));
 sky130_fd_sc_hd__xnor2_2 _08857_ (.A(net205),
    .B(_01948_),
    .Y(_01949_));
 sky130_fd_sc_hd__a31o_2 _08858_ (.A1(_04926_),
    .A2(_05013_),
    .A3(_00139_),
    .B1(net183),
    .X(_01950_));
 sky130_fd_sc_hd__xnor2_4 _08859_ (.A(_05100_),
    .B(_01950_),
    .Y(_01951_));
 sky130_fd_sc_hd__xnor2_1 _08860_ (.A(_05089_),
    .B(_01950_),
    .Y(_01952_));
 sky130_fd_sc_hd__a22o_1 _08861_ (.A1(_06519_),
    .A2(_00700_),
    .B1(_01951_),
    .B2(net292),
    .X(_01953_));
 sky130_fd_sc_hd__xnor2_2 _08862_ (.A(_06493_),
    .B(_01953_),
    .Y(_01954_));
 sky130_fd_sc_hd__o22a_1 _08863_ (.A1(net68),
    .A2(net156),
    .B1(net154),
    .B2(net65),
    .X(_01955_));
 sky130_fd_sc_hd__xnor2_2 _08864_ (.A(net207),
    .B(_01955_),
    .Y(_01956_));
 sky130_fd_sc_hd__or2_1 _08865_ (.A(_01954_),
    .B(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__xnor2_2 _08866_ (.A(_01954_),
    .B(_01956_),
    .Y(_01958_));
 sky130_fd_sc_hd__xor2_2 _08867_ (.A(_01949_),
    .B(_01958_),
    .X(_01959_));
 sky130_fd_sc_hd__xnor2_1 _08868_ (.A(_01947_),
    .B(_01959_),
    .Y(_01960_));
 sky130_fd_sc_hd__xnor2_1 _08869_ (.A(_01936_),
    .B(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__or4_1 _08870_ (.A(reg1_val[28]),
    .B(reg1_val[29]),
    .C(_00233_),
    .D(_00449_),
    .X(_01962_));
 sky130_fd_sc_hd__o41a_1 _08871_ (.A1(reg1_val[28]),
    .A2(reg1_val[29]),
    .A3(_00233_),
    .A4(_00449_),
    .B1(net262),
    .X(_01963_));
 sky130_fd_sc_hd__xnor2_2 _08872_ (.A(reg1_val[30]),
    .B(_01963_),
    .Y(_01964_));
 sky130_fd_sc_hd__or2_1 _08873_ (.A(net69),
    .B(_01964_),
    .X(_01965_));
 sky130_fd_sc_hd__nand2_1 _08874_ (.A(net69),
    .B(_01964_),
    .Y(_01966_));
 sky130_fd_sc_hd__and2_1 _08875_ (.A(_01965_),
    .B(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__nand2_1 _08876_ (.A(_01965_),
    .B(_01966_),
    .Y(_01968_));
 sky130_fd_sc_hd__nor2_2 _08877_ (.A(net216),
    .B(net11),
    .Y(_01969_));
 sky130_fd_sc_hd__o22a_1 _08878_ (.A1(_00264_),
    .A2(net24),
    .B1(net16),
    .B2(net144),
    .X(_01970_));
 sky130_fd_sc_hd__xnor2_2 _08879_ (.A(net71),
    .B(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__xor2_2 _08880_ (.A(_01969_),
    .B(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__or2_1 _08881_ (.A(_01961_),
    .B(_01972_),
    .X(_01973_));
 sky130_fd_sc_hd__xnor2_1 _08882_ (.A(_01961_),
    .B(_01972_),
    .Y(_01974_));
 sky130_fd_sc_hd__xor2_1 _08883_ (.A(_01926_),
    .B(_01974_),
    .X(_01975_));
 sky130_fd_sc_hd__a21oi_1 _08884_ (.A1(_00673_),
    .A2(_00675_),
    .B1(_00671_),
    .Y(_01976_));
 sky130_fd_sc_hd__o22a_1 _08885_ (.A1(net120),
    .A2(net27),
    .B1(net25),
    .B2(_00290_),
    .X(_01977_));
 sky130_fd_sc_hd__xnor2_1 _08886_ (.A(net88),
    .B(_01977_),
    .Y(_01978_));
 sky130_fd_sc_hd__a22o_1 _08887_ (.A1(net31),
    .A2(_00324_),
    .B1(_00330_),
    .B2(net29),
    .X(_01979_));
 sky130_fd_sc_hd__xnor2_1 _08888_ (.A(net49),
    .B(_01979_),
    .Y(_01980_));
 sky130_fd_sc_hd__and2_2 _08889_ (.A(_01978_),
    .B(_01980_),
    .X(_01981_));
 sky130_fd_sc_hd__nor2_1 _08890_ (.A(_01978_),
    .B(_01980_),
    .Y(_01982_));
 sky130_fd_sc_hd__or2_1 _08891_ (.A(_01981_),
    .B(_01982_),
    .X(_01983_));
 sky130_fd_sc_hd__a21oi_1 _08892_ (.A1(_00725_),
    .A2(_00730_),
    .B1(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__and3_1 _08893_ (.A(_00725_),
    .B(_00730_),
    .C(_01983_),
    .X(_01985_));
 sky130_fd_sc_hd__nor2_1 _08894_ (.A(_01984_),
    .B(_01985_),
    .Y(_01986_));
 sky130_fd_sc_hd__and2b_1 _08895_ (.A_N(_01976_),
    .B(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__xnor2_1 _08896_ (.A(_01976_),
    .B(_01986_),
    .Y(_01988_));
 sky130_fd_sc_hd__and2_1 _08897_ (.A(_01975_),
    .B(_01988_),
    .X(_01989_));
 sky130_fd_sc_hd__nor2_1 _08898_ (.A(_01975_),
    .B(_01988_),
    .Y(_01990_));
 sky130_fd_sc_hd__nor2_2 _08899_ (.A(_01989_),
    .B(_01990_),
    .Y(_01991_));
 sky130_fd_sc_hd__xor2_4 _08900_ (.A(_01921_),
    .B(_01991_),
    .X(_01992_));
 sky130_fd_sc_hd__a32o_1 _08901_ (.A1(_00735_),
    .A2(_00736_),
    .A3(_00750_),
    .B1(_00751_),
    .B2(_00684_),
    .X(_01993_));
 sky130_fd_sc_hd__o21bai_4 _08902_ (.A1(_00666_),
    .A2(_00682_),
    .B1_N(_00681_),
    .Y(_01994_));
 sky130_fd_sc_hd__a21o_2 _08903_ (.A1(_00694_),
    .A2(_00734_),
    .B1(_00733_),
    .X(_01995_));
 sky130_fd_sc_hd__nor2_2 _08904_ (.A(_00746_),
    .B(_00749_),
    .Y(_01996_));
 sky130_fd_sc_hd__o21ai_1 _08905_ (.A1(_00746_),
    .A2(_00749_),
    .B1(_01995_),
    .Y(_01997_));
 sky130_fd_sc_hd__xnor2_4 _08906_ (.A(_01995_),
    .B(_01996_),
    .Y(_01998_));
 sky130_fd_sc_hd__xnor2_4 _08907_ (.A(_01994_),
    .B(_01998_),
    .Y(_01999_));
 sky130_fd_sc_hd__a21oi_2 _08908_ (.A1(_00754_),
    .A2(_00758_),
    .B1(_00757_),
    .Y(_02000_));
 sky130_fd_sc_hd__xnor2_2 _08909_ (.A(_01999_),
    .B(_02000_),
    .Y(_02001_));
 sky130_fd_sc_hd__nand2b_1 _08910_ (.A_N(_02001_),
    .B(_01993_),
    .Y(_02002_));
 sky130_fd_sc_hd__xnor2_2 _08911_ (.A(_01993_),
    .B(_02001_),
    .Y(_02003_));
 sky130_fd_sc_hd__xnor2_2 _08912_ (.A(_01992_),
    .B(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__nand2b_1 _08913_ (.A_N(_02004_),
    .B(_01905_),
    .Y(_02005_));
 sky130_fd_sc_hd__xor2_4 _08914_ (.A(_01905_),
    .B(_02004_),
    .X(_02006_));
 sky130_fd_sc_hd__or2_1 _08915_ (.A(_01904_),
    .B(_02006_),
    .X(_02007_));
 sky130_fd_sc_hd__and2_1 _08916_ (.A(_01904_),
    .B(_02006_),
    .X(_02008_));
 sky130_fd_sc_hd__xnor2_4 _08917_ (.A(_01904_),
    .B(_02006_),
    .Y(_02009_));
 sky130_fd_sc_hd__o22a_1 _08918_ (.A1(_00664_),
    .A2(_00766_),
    .B1(_00769_),
    .B2(_00838_),
    .X(_02010_));
 sky130_fd_sc_hd__a21o_1 _08919_ (.A1(_00664_),
    .A2(_00766_),
    .B1(_02010_),
    .X(_02011_));
 sky130_fd_sc_hd__or2_1 _08920_ (.A(_00768_),
    .B(_01800_),
    .X(_02012_));
 sky130_fd_sc_hd__a211o_1 _08921_ (.A1(_01888_),
    .A2(_01889_),
    .B1(_00768_),
    .C1(_01800_),
    .X(_02013_));
 sky130_fd_sc_hd__o221a_2 _08922_ (.A1(_01896_),
    .A2(_02012_),
    .B1(_02013_),
    .B2(_01897_),
    .C1(_02011_),
    .X(_02014_));
 sky130_fd_sc_hd__xnor2_2 _08923_ (.A(_02009_),
    .B(_02014_),
    .Y(_02015_));
 sky130_fd_sc_hd__and3_1 _08924_ (.A(_01895_),
    .B(_01903_),
    .C(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__a21bo_2 _08925_ (.A1(_01992_),
    .A2(_02003_),
    .B1_N(_02005_),
    .X(_02017_));
 sky130_fd_sc_hd__o21ai_4 _08926_ (.A1(_01999_),
    .A2(_02000_),
    .B1(_02002_),
    .Y(_02018_));
 sky130_fd_sc_hd__a32o_1 _08927_ (.A1(_01945_),
    .A2(_01946_),
    .A3(_01959_),
    .B1(_01960_),
    .B2(_01936_),
    .X(_02019_));
 sky130_fd_sc_hd__o22a_1 _08928_ (.A1(net46),
    .A2(_00309_),
    .B1(net110),
    .B2(net48),
    .X(_02020_));
 sky130_fd_sc_hd__xnor2_1 _08929_ (.A(net97),
    .B(_02020_),
    .Y(_02021_));
 sky130_fd_sc_hd__a22o_1 _08930_ (.A1(_00213_),
    .A2(net44),
    .B1(net42),
    .B2(_00226_),
    .X(_02022_));
 sky130_fd_sc_hd__xor2_1 _08931_ (.A(net94),
    .B(_02022_),
    .X(_02023_));
 sky130_fd_sc_hd__and2_1 _08932_ (.A(_02021_),
    .B(_02023_),
    .X(_02024_));
 sky130_fd_sc_hd__nor2_1 _08933_ (.A(_02021_),
    .B(_02023_),
    .Y(_02025_));
 sky130_fd_sc_hd__nor2_1 _08934_ (.A(_02024_),
    .B(_02025_),
    .Y(_02026_));
 sky130_fd_sc_hd__a22o_1 _08935_ (.A1(net39),
    .A2(net113),
    .B1(_00374_),
    .B2(net37),
    .X(_02027_));
 sky130_fd_sc_hd__xor2_2 _08936_ (.A(net91),
    .B(_02027_),
    .X(_02028_));
 sky130_fd_sc_hd__xor2_2 _08937_ (.A(_02026_),
    .B(_02028_),
    .X(_02029_));
 sky130_fd_sc_hd__a21bo_1 _08938_ (.A1(_01922_),
    .A2(_01925_),
    .B1_N(_01924_),
    .X(_02030_));
 sky130_fd_sc_hd__xnor2_1 _08939_ (.A(_02029_),
    .B(_02030_),
    .Y(_02031_));
 sky130_fd_sc_hd__and2b_1 _08940_ (.A_N(_02031_),
    .B(_02019_),
    .X(_02032_));
 sky130_fd_sc_hd__and2b_1 _08941_ (.A_N(_02019_),
    .B(_02031_),
    .X(_02033_));
 sky130_fd_sc_hd__nor2_2 _08942_ (.A(_02032_),
    .B(_02033_),
    .Y(_02034_));
 sky130_fd_sc_hd__and2b_1 _08943_ (.A_N(_01941_),
    .B(_01945_),
    .X(_02035_));
 sky130_fd_sc_hd__a21oi_2 _08944_ (.A1(_01932_),
    .A2(_01935_),
    .B1(_01931_),
    .Y(_02036_));
 sky130_fd_sc_hd__nand2b_1 _08945_ (.A_N(_02036_),
    .B(_01981_),
    .Y(_02037_));
 sky130_fd_sc_hd__xnor2_2 _08946_ (.A(_01981_),
    .B(_02036_),
    .Y(_02038_));
 sky130_fd_sc_hd__nand2b_1 _08947_ (.A_N(_02035_),
    .B(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__xnor2_2 _08948_ (.A(_02035_),
    .B(_02038_),
    .Y(_02040_));
 sky130_fd_sc_hd__o22a_1 _08949_ (.A1(net61),
    .A2(net106),
    .B1(net104),
    .B2(net53),
    .X(_02041_));
 sky130_fd_sc_hd__xnor2_1 _08950_ (.A(net135),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__o22a_1 _08951_ (.A1(net65),
    .A2(_00160_),
    .B1(net146),
    .B2(net59),
    .X(_02043_));
 sky130_fd_sc_hd__xnor2_1 _08952_ (.A(net202),
    .B(_02043_),
    .Y(_02044_));
 sky130_fd_sc_hd__nor2_1 _08953_ (.A(_02042_),
    .B(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__xor2_1 _08954_ (.A(_02042_),
    .B(_02044_),
    .X(_02046_));
 sky130_fd_sc_hd__o22a_1 _08955_ (.A1(net57),
    .A2(net134),
    .B1(net132),
    .B2(net63),
    .X(_02047_));
 sky130_fd_sc_hd__xnor2_1 _08956_ (.A(net181),
    .B(_02047_),
    .Y(_02048_));
 sky130_fd_sc_hd__and2b_1 _08957_ (.A_N(_02048_),
    .B(_02046_),
    .X(_02049_));
 sky130_fd_sc_hd__and2b_1 _08958_ (.A_N(_02046_),
    .B(_02048_),
    .X(_02050_));
 sky130_fd_sc_hd__nor2_1 _08959_ (.A(_02049_),
    .B(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hd__o22a_1 _08960_ (.A1(net51),
    .A2(net86),
    .B1(net82),
    .B2(net100),
    .X(_02052_));
 sky130_fd_sc_hd__xnor2_1 _08961_ (.A(net137),
    .B(_02052_),
    .Y(_02053_));
 sky130_fd_sc_hd__o22a_1 _08962_ (.A1(net35),
    .A2(net81),
    .B1(net77),
    .B2(net33),
    .X(_02054_));
 sky130_fd_sc_hd__xnor2_1 _08963_ (.A(net125),
    .B(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__and2b_1 _08964_ (.A_N(_02053_),
    .B(_02055_),
    .X(_02056_));
 sky130_fd_sc_hd__xor2_1 _08965_ (.A(_02053_),
    .B(_02055_),
    .X(_02057_));
 sky130_fd_sc_hd__o22a_1 _08966_ (.A1(net98),
    .A2(net78),
    .B1(net74),
    .B2(net84),
    .X(_02058_));
 sky130_fd_sc_hd__xnor2_1 _08967_ (.A(net121),
    .B(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__or2_1 _08968_ (.A(_02057_),
    .B(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__nand2_1 _08969_ (.A(_02057_),
    .B(_02059_),
    .Y(_02061_));
 sky130_fd_sc_hd__nand2_1 _08970_ (.A(_02060_),
    .B(_02061_),
    .Y(_02062_));
 sky130_fd_sc_hd__o22a_2 _08971_ (.A1(net150),
    .A2(net17),
    .B1(net14),
    .B2(net152),
    .X(_02063_));
 sky130_fd_sc_hd__xnor2_4 _08972_ (.A(net205),
    .B(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__or4_2 _08973_ (.A(_04937_),
    .B(_05024_),
    .C(_05100_),
    .D(_00140_),
    .X(_02065_));
 sky130_fd_sc_hd__a21oi_4 _08974_ (.A1(net295),
    .A2(_02065_),
    .B1(_05371_),
    .Y(_02066_));
 sky130_fd_sc_hd__a21o_2 _08975_ (.A1(net295),
    .A2(_02065_),
    .B1(_05371_),
    .X(_02067_));
 sky130_fd_sc_hd__o22a_2 _08976_ (.A1(_06520_),
    .A2(net13),
    .B1(net8),
    .B2(net288),
    .X(_02068_));
 sky130_fd_sc_hd__xnor2_4 _08977_ (.A(net239),
    .B(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__o22a_2 _08978_ (.A1(net68),
    .A2(net154),
    .B1(net56),
    .B2(_06538_),
    .X(_02070_));
 sky130_fd_sc_hd__xnor2_4 _08979_ (.A(net207),
    .B(_02070_),
    .Y(_02071_));
 sky130_fd_sc_hd__or2_1 _08980_ (.A(_02069_),
    .B(_02071_),
    .X(_02072_));
 sky130_fd_sc_hd__xnor2_4 _08981_ (.A(_02069_),
    .B(_02071_),
    .Y(_02073_));
 sky130_fd_sc_hd__xor2_4 _08982_ (.A(_02064_),
    .B(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__xnor2_2 _08983_ (.A(_02062_),
    .B(_02074_),
    .Y(_02075_));
 sky130_fd_sc_hd__xnor2_2 _08984_ (.A(_02051_),
    .B(_02075_),
    .Y(_02076_));
 sky130_fd_sc_hd__nor2_1 _08985_ (.A(reg1_val[30]),
    .B(_01962_),
    .Y(_02077_));
 sky130_fd_sc_hd__o21a_4 _08986_ (.A1(net286),
    .A2(_02077_),
    .B1(reg1_val[31]),
    .X(_02078_));
 sky130_fd_sc_hd__o21ai_4 _08987_ (.A1(net286),
    .A2(_02077_),
    .B1(reg1_val[31]),
    .Y(_02079_));
 sky130_fd_sc_hd__a2111o_1 _08988_ (.A1(net294),
    .A2(_01962_),
    .B1(_00678_),
    .C1(reg1_val[30]),
    .D1(_04531_),
    .X(_02080_));
 sky130_fd_sc_hd__o21a_1 _08989_ (.A1(_01965_),
    .A2(_02078_),
    .B1(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__o21ai_1 _08990_ (.A1(_01965_),
    .A2(net22),
    .B1(_02080_),
    .Y(_02082_));
 sky130_fd_sc_hd__o22a_2 _08991_ (.A1(net144),
    .A2(net11),
    .B1(net6),
    .B2(net216),
    .X(_02083_));
 sky130_fd_sc_hd__xnor2_4 _08992_ (.A(net21),
    .B(_02083_),
    .Y(_02084_));
 sky130_fd_sc_hd__o21a_2 _08993_ (.A1(_01949_),
    .A2(_01958_),
    .B1(_01957_),
    .X(_02085_));
 sky130_fd_sc_hd__o22a_1 _08994_ (.A1(net142),
    .A2(net24),
    .B1(net16),
    .B2(_00264_),
    .X(_02086_));
 sky130_fd_sc_hd__xnor2_2 _08995_ (.A(_00678_),
    .B(_02086_),
    .Y(_02087_));
 sky130_fd_sc_hd__and2b_1 _08996_ (.A_N(_02085_),
    .B(_02087_),
    .X(_02088_));
 sky130_fd_sc_hd__xor2_4 _08997_ (.A(_02085_),
    .B(_02087_),
    .X(_02089_));
 sky130_fd_sc_hd__xnor2_4 _08998_ (.A(_02084_),
    .B(_02089_),
    .Y(_02090_));
 sky130_fd_sc_hd__nor2_1 _08999_ (.A(_02076_),
    .B(_02090_),
    .Y(_02091_));
 sky130_fd_sc_hd__xor2_2 _09000_ (.A(_02076_),
    .B(_02090_),
    .X(_02092_));
 sky130_fd_sc_hd__xor2_1 _09001_ (.A(_02040_),
    .B(_02092_),
    .X(_02093_));
 sky130_fd_sc_hd__a21o_1 _09002_ (.A1(_01914_),
    .A2(_01916_),
    .B1(_01912_),
    .X(_02094_));
 sky130_fd_sc_hd__o22a_1 _09003_ (.A1(net120),
    .A2(net25),
    .B1(net73),
    .B2(net27),
    .X(_02095_));
 sky130_fd_sc_hd__xnor2_1 _09004_ (.A(net88),
    .B(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__a22o_1 _09005_ (.A1(net116),
    .A2(net31),
    .B1(net29),
    .B2(_00324_),
    .X(_02097_));
 sky130_fd_sc_hd__xnor2_1 _09006_ (.A(net49),
    .B(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__and2_1 _09007_ (.A(_02096_),
    .B(_02098_),
    .X(_02099_));
 sky130_fd_sc_hd__nor2_1 _09008_ (.A(_02096_),
    .B(_02098_),
    .Y(_02100_));
 sky130_fd_sc_hd__nor2_1 _09009_ (.A(_02099_),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__nor2_1 _09010_ (.A(_01969_),
    .B(net22),
    .Y(_02102_));
 sky130_fd_sc_hd__a21oi_2 _09011_ (.A1(_01969_),
    .A2(_01971_),
    .B1(_02102_),
    .Y(_02103_));
 sky130_fd_sc_hd__xnor2_1 _09012_ (.A(_02101_),
    .B(_02103_),
    .Y(_02104_));
 sky130_fd_sc_hd__and2b_1 _09013_ (.A_N(_02104_),
    .B(_02094_),
    .X(_02105_));
 sky130_fd_sc_hd__xnor2_1 _09014_ (.A(_02094_),
    .B(_02104_),
    .Y(_02106_));
 sky130_fd_sc_hd__nand2_1 _09015_ (.A(_02093_),
    .B(_02106_),
    .Y(_02107_));
 sky130_fd_sc_hd__or2_1 _09016_ (.A(_02093_),
    .B(_02106_),
    .X(_02108_));
 sky130_fd_sc_hd__and2_2 _09017_ (.A(_02107_),
    .B(_02108_),
    .X(_02109_));
 sky130_fd_sc_hd__xor2_4 _09018_ (.A(_02034_),
    .B(_02109_),
    .X(_02110_));
 sky130_fd_sc_hd__a21o_2 _09019_ (.A1(_01921_),
    .A2(_01991_),
    .B1(_01989_),
    .X(_02111_));
 sky130_fd_sc_hd__a21o_2 _09020_ (.A1(_01907_),
    .A2(_01917_),
    .B1(_01919_),
    .X(_02112_));
 sky130_fd_sc_hd__o21a_2 _09021_ (.A1(_01926_),
    .A2(_01974_),
    .B1(_01973_),
    .X(_02113_));
 sky130_fd_sc_hd__nor2_2 _09022_ (.A(_01984_),
    .B(_01987_),
    .Y(_02114_));
 sky130_fd_sc_hd__nor2_1 _09023_ (.A(_02113_),
    .B(_02114_),
    .Y(_02115_));
 sky130_fd_sc_hd__xor2_4 _09024_ (.A(_02113_),
    .B(_02114_),
    .X(_02116_));
 sky130_fd_sc_hd__xnor2_4 _09025_ (.A(_02112_),
    .B(_02116_),
    .Y(_02117_));
 sky130_fd_sc_hd__a21boi_4 _09026_ (.A1(_01994_),
    .A2(_01998_),
    .B1_N(_01997_),
    .Y(_02118_));
 sky130_fd_sc_hd__xnor2_4 _09027_ (.A(_02117_),
    .B(_02118_),
    .Y(_02119_));
 sky130_fd_sc_hd__nand2b_1 _09028_ (.A_N(_02119_),
    .B(_02111_),
    .Y(_02120_));
 sky130_fd_sc_hd__xnor2_4 _09029_ (.A(_02111_),
    .B(_02119_),
    .Y(_02121_));
 sky130_fd_sc_hd__and2_1 _09030_ (.A(_02110_),
    .B(_02121_),
    .X(_02122_));
 sky130_fd_sc_hd__xor2_4 _09031_ (.A(_02110_),
    .B(_02121_),
    .X(_02123_));
 sky130_fd_sc_hd__xor2_4 _09032_ (.A(_02018_),
    .B(_02123_),
    .X(_02124_));
 sky130_fd_sc_hd__nor2_1 _09033_ (.A(_02017_),
    .B(_02124_),
    .Y(_02125_));
 sky130_fd_sc_hd__xnor2_4 _09034_ (.A(_02017_),
    .B(_02124_),
    .Y(_02126_));
 sky130_fd_sc_hd__a21o_1 _09035_ (.A1(_00767_),
    .A2(_02007_),
    .B1(_02008_),
    .X(_02127_));
 sky130_fd_sc_hd__nor2_1 _09036_ (.A(_00768_),
    .B(_02009_),
    .Y(_02128_));
 sky130_fd_sc_hd__or2_1 _09037_ (.A(_00768_),
    .B(_02009_),
    .X(_02129_));
 sky130_fd_sc_hd__a21boi_2 _09038_ (.A1(_01801_),
    .A2(_02128_),
    .B1_N(_02127_),
    .Y(_02130_));
 sky130_fd_sc_hd__xnor2_2 _09039_ (.A(_02126_),
    .B(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__nand4_2 _09040_ (.A(_01895_),
    .B(_01903_),
    .C(_02015_),
    .D(_02131_),
    .Y(_02132_));
 sky130_fd_sc_hd__a2111o_1 _09041_ (.A1(_01896_),
    .A2(_01898_),
    .B1(_02009_),
    .C1(_02012_),
    .D1(_02126_),
    .X(_02133_));
 sky130_fd_sc_hd__a21boi_1 _09042_ (.A1(_02017_),
    .A2(_02124_),
    .B1_N(_02007_),
    .Y(_02134_));
 sky130_fd_sc_hd__o32a_1 _09043_ (.A1(_02009_),
    .A2(_02011_),
    .A3(_02126_),
    .B1(_02134_),
    .B2(_02125_),
    .X(_02135_));
 sky130_fd_sc_hd__nand2_1 _09044_ (.A(_02133_),
    .B(_02135_),
    .Y(_02136_));
 sky130_fd_sc_hd__a21oi_4 _09045_ (.A1(_02018_),
    .A2(_02123_),
    .B1(_02122_),
    .Y(_02137_));
 sky130_fd_sc_hd__o21ai_4 _09046_ (.A1(_02117_),
    .A2(_02118_),
    .B1(_02120_),
    .Y(_02138_));
 sky130_fd_sc_hd__a32o_2 _09047_ (.A1(_02060_),
    .A2(_02061_),
    .A3(_02074_),
    .B1(_02075_),
    .B2(_02051_),
    .X(_02139_));
 sky130_fd_sc_hd__o22a_1 _09048_ (.A1(net128),
    .A2(net24),
    .B1(net16),
    .B2(net142),
    .X(_02140_));
 sky130_fd_sc_hd__xnor2_2 _09049_ (.A(net71),
    .B(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__inv_2 _09050_ (.A(_02141_),
    .Y(_02142_));
 sky130_fd_sc_hd__a22o_1 _09051_ (.A1(net39),
    .A2(_00308_),
    .B1(net113),
    .B2(net37),
    .X(_02143_));
 sky130_fd_sc_hd__xor2_1 _09052_ (.A(net91),
    .B(_02143_),
    .X(_02144_));
 sky130_fd_sc_hd__xor2_1 _09053_ (.A(_02141_),
    .B(_02144_),
    .X(_02145_));
 sky130_fd_sc_hd__a22o_1 _09054_ (.A1(_00213_),
    .A2(net42),
    .B1(_00374_),
    .B2(net44),
    .X(_02146_));
 sky130_fd_sc_hd__xor2_1 _09055_ (.A(net94),
    .B(_02146_),
    .X(_02147_));
 sky130_fd_sc_hd__and2b_1 _09056_ (.A_N(_02145_),
    .B(_02147_),
    .X(_02148_));
 sky130_fd_sc_hd__and2b_1 _09057_ (.A_N(_02147_),
    .B(_02145_),
    .X(_02149_));
 sky130_fd_sc_hd__or2_1 _09058_ (.A(_02148_),
    .B(_02149_),
    .X(_02150_));
 sky130_fd_sc_hd__a21o_1 _09059_ (.A1(_02037_),
    .A2(_02039_),
    .B1(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__nand3_1 _09060_ (.A(_02037_),
    .B(_02039_),
    .C(_02150_),
    .Y(_02152_));
 sky130_fd_sc_hd__nand2_2 _09061_ (.A(_02151_),
    .B(_02152_),
    .Y(_02153_));
 sky130_fd_sc_hd__nand2b_1 _09062_ (.A_N(_02153_),
    .B(_02139_),
    .Y(_02154_));
 sky130_fd_sc_hd__xnor2_4 _09063_ (.A(_02139_),
    .B(_02153_),
    .Y(_02155_));
 sky130_fd_sc_hd__and2b_1 _09064_ (.A_N(_02056_),
    .B(_02060_),
    .X(_02156_));
 sky130_fd_sc_hd__o21ai_1 _09065_ (.A1(_02045_),
    .A2(_02049_),
    .B1(_02099_),
    .Y(_02157_));
 sky130_fd_sc_hd__or3_1 _09066_ (.A(_02045_),
    .B(_02049_),
    .C(_02099_),
    .X(_02158_));
 sky130_fd_sc_hd__and2_1 _09067_ (.A(_02157_),
    .B(_02158_),
    .X(_02159_));
 sky130_fd_sc_hd__nand2b_1 _09068_ (.A_N(_02156_),
    .B(_02159_),
    .Y(_02160_));
 sky130_fd_sc_hd__xnor2_2 _09069_ (.A(_02156_),
    .B(_02159_),
    .Y(_02161_));
 sky130_fd_sc_hd__o22a_1 _09070_ (.A1(net68),
    .A2(_00160_),
    .B1(net146),
    .B2(net65),
    .X(_02162_));
 sky130_fd_sc_hd__xnor2_2 _09071_ (.A(net202),
    .B(_02162_),
    .Y(_02163_));
 sky130_fd_sc_hd__o22a_1 _09072_ (.A1(net63),
    .A2(net106),
    .B1(net104),
    .B2(net61),
    .X(_02164_));
 sky130_fd_sc_hd__xnor2_2 _09073_ (.A(net135),
    .B(_02164_),
    .Y(_02165_));
 sky130_fd_sc_hd__nor2_1 _09074_ (.A(_02163_),
    .B(_02165_),
    .Y(_02166_));
 sky130_fd_sc_hd__xor2_2 _09075_ (.A(_02163_),
    .B(_02165_),
    .X(_02167_));
 sky130_fd_sc_hd__o22a_1 _09076_ (.A1(net59),
    .A2(net134),
    .B1(net132),
    .B2(net57),
    .X(_02168_));
 sky130_fd_sc_hd__xnor2_2 _09077_ (.A(net181),
    .B(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__inv_2 _09078_ (.A(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__xnor2_2 _09079_ (.A(_02167_),
    .B(_02169_),
    .Y(_02171_));
 sky130_fd_sc_hd__o22a_1 _09080_ (.A1(net53),
    .A2(net86),
    .B1(net82),
    .B2(net51),
    .X(_02172_));
 sky130_fd_sc_hd__xnor2_1 _09081_ (.A(net137),
    .B(_02172_),
    .Y(_02173_));
 sky130_fd_sc_hd__o22a_1 _09082_ (.A1(net35),
    .A2(net84),
    .B1(net81),
    .B2(net33),
    .X(_02174_));
 sky130_fd_sc_hd__xnor2_1 _09083_ (.A(net125),
    .B(_02174_),
    .Y(_02175_));
 sky130_fd_sc_hd__and2b_1 _09084_ (.A_N(_02173_),
    .B(_02175_),
    .X(_02176_));
 sky130_fd_sc_hd__xor2_1 _09085_ (.A(_02173_),
    .B(_02175_),
    .X(_02177_));
 sky130_fd_sc_hd__o22a_1 _09086_ (.A1(net100),
    .A2(net78),
    .B1(net74),
    .B2(net98),
    .X(_02178_));
 sky130_fd_sc_hd__xnor2_1 _09087_ (.A(net121),
    .B(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hd__or2_1 _09088_ (.A(_02177_),
    .B(_02179_),
    .X(_02180_));
 sky130_fd_sc_hd__nand2_1 _09089_ (.A(_02177_),
    .B(_02179_),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2_1 _09090_ (.A(_02180_),
    .B(_02181_),
    .Y(_02182_));
 sky130_fd_sc_hd__o22a_1 _09091_ (.A1(net150),
    .A2(net14),
    .B1(net13),
    .B2(net152),
    .X(_02183_));
 sky130_fd_sc_hd__xor2_1 _09092_ (.A(net205),
    .B(_02183_),
    .X(_02184_));
 sky130_fd_sc_hd__o32a_1 _09093_ (.A1(net156),
    .A2(_00405_),
    .A3(_00407_),
    .B1(net154),
    .B2(net56),
    .X(_02185_));
 sky130_fd_sc_hd__xnor2_1 _09094_ (.A(_06532_),
    .B(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__a21oi_1 _09095_ (.A1(net288),
    .A2(net9),
    .B1(net239),
    .Y(_02187_));
 sky130_fd_sc_hd__nand2_1 _09096_ (.A(_02186_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__xor2_1 _09097_ (.A(_02186_),
    .B(_02187_),
    .X(_02189_));
 sky130_fd_sc_hd__nand2_1 _09098_ (.A(_02184_),
    .B(_02189_),
    .Y(_02190_));
 sky130_fd_sc_hd__or2_1 _09099_ (.A(_02184_),
    .B(_02189_),
    .X(_02191_));
 sky130_fd_sc_hd__and2_2 _09100_ (.A(_02190_),
    .B(_02191_),
    .X(_02192_));
 sky130_fd_sc_hd__xnor2_2 _09101_ (.A(_02182_),
    .B(_02192_),
    .Y(_02193_));
 sky130_fd_sc_hd__xnor2_2 _09102_ (.A(_02171_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__nor2_1 _09103_ (.A(_06364_),
    .B(net21),
    .Y(_02195_));
 sky130_fd_sc_hd__o21ai_2 _09104_ (.A1(_02064_),
    .A2(_02073_),
    .B1(_02072_),
    .Y(_02196_));
 sky130_fd_sc_hd__o22a_1 _09105_ (.A1(_00264_),
    .A2(net11),
    .B1(net6),
    .B2(net144),
    .X(_02197_));
 sky130_fd_sc_hd__xnor2_2 _09106_ (.A(net22),
    .B(_02197_),
    .Y(_02198_));
 sky130_fd_sc_hd__nand2_1 _09107_ (.A(_02196_),
    .B(_02198_),
    .Y(_02199_));
 sky130_fd_sc_hd__xor2_2 _09108_ (.A(_02196_),
    .B(_02198_),
    .X(_02200_));
 sky130_fd_sc_hd__xnor2_2 _09109_ (.A(_02195_),
    .B(_02200_),
    .Y(_02201_));
 sky130_fd_sc_hd__nor2_1 _09110_ (.A(_02194_),
    .B(_02201_),
    .Y(_02202_));
 sky130_fd_sc_hd__xor2_2 _09111_ (.A(_02194_),
    .B(_02201_),
    .X(_02203_));
 sky130_fd_sc_hd__xnor2_1 _09112_ (.A(_02161_),
    .B(_02203_),
    .Y(_02204_));
 sky130_fd_sc_hd__a21o_1 _09113_ (.A1(_02026_),
    .A2(_02028_),
    .B1(_02024_),
    .X(_02205_));
 sky130_fd_sc_hd__o22a_1 _09114_ (.A1(net27),
    .A2(net77),
    .B1(net73),
    .B2(net25),
    .X(_02206_));
 sky130_fd_sc_hd__xnor2_2 _09115_ (.A(net88),
    .B(_02206_),
    .Y(_02207_));
 sky130_fd_sc_hd__o22a_1 _09116_ (.A1(net48),
    .A2(net112),
    .B1(net110),
    .B2(net46),
    .X(_02208_));
 sky130_fd_sc_hd__xnor2_2 _09117_ (.A(net97),
    .B(_02208_),
    .Y(_02209_));
 sky130_fd_sc_hd__and2_1 _09118_ (.A(_02207_),
    .B(_02209_),
    .X(_02210_));
 sky130_fd_sc_hd__xor2_2 _09119_ (.A(_02207_),
    .B(_02209_),
    .X(_02211_));
 sky130_fd_sc_hd__a22o_1 _09120_ (.A1(net118),
    .A2(net31),
    .B1(net29),
    .B2(net116),
    .X(_02212_));
 sky130_fd_sc_hd__xnor2_2 _09121_ (.A(net50),
    .B(_02212_),
    .Y(_02213_));
 sky130_fd_sc_hd__xor2_2 _09122_ (.A(_02211_),
    .B(_02213_),
    .X(_02214_));
 sky130_fd_sc_hd__o21ba_1 _09123_ (.A1(_02084_),
    .A2(_02089_),
    .B1_N(_02088_),
    .X(_02215_));
 sky130_fd_sc_hd__and2b_1 _09124_ (.A_N(_02215_),
    .B(_02214_),
    .X(_02216_));
 sky130_fd_sc_hd__xnor2_2 _09125_ (.A(_02214_),
    .B(_02215_),
    .Y(_02217_));
 sky130_fd_sc_hd__xnor2_1 _09126_ (.A(_02205_),
    .B(_02217_),
    .Y(_02218_));
 sky130_fd_sc_hd__nor2_1 _09127_ (.A(_02204_),
    .B(_02218_),
    .Y(_02219_));
 sky130_fd_sc_hd__nand2_1 _09128_ (.A(_02204_),
    .B(_02218_),
    .Y(_02220_));
 sky130_fd_sc_hd__and2b_1 _09129_ (.A_N(_02219_),
    .B(_02220_),
    .X(_02221_));
 sky130_fd_sc_hd__xor2_4 _09130_ (.A(_02155_),
    .B(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__a21bo_2 _09131_ (.A1(_02034_),
    .A2(_02109_),
    .B1_N(_02107_),
    .X(_02223_));
 sky130_fd_sc_hd__a21o_2 _09132_ (.A1(_02029_),
    .A2(_02030_),
    .B1(_02032_),
    .X(_02224_));
 sky130_fd_sc_hd__a21oi_4 _09133_ (.A1(_02040_),
    .A2(_02092_),
    .B1(_02091_),
    .Y(_02225_));
 sky130_fd_sc_hd__a21oi_4 _09134_ (.A1(_02101_),
    .A2(_02103_),
    .B1(_02105_),
    .Y(_02226_));
 sky130_fd_sc_hd__nor2_1 _09135_ (.A(_02225_),
    .B(_02226_),
    .Y(_02227_));
 sky130_fd_sc_hd__xor2_4 _09136_ (.A(_02225_),
    .B(_02226_),
    .X(_02228_));
 sky130_fd_sc_hd__xnor2_4 _09137_ (.A(_02224_),
    .B(_02228_),
    .Y(_02229_));
 sky130_fd_sc_hd__a21oi_4 _09138_ (.A1(_02112_),
    .A2(_02116_),
    .B1(_02115_),
    .Y(_02230_));
 sky130_fd_sc_hd__xnor2_2 _09139_ (.A(_02229_),
    .B(_02230_),
    .Y(_02231_));
 sky130_fd_sc_hd__nand2b_1 _09140_ (.A_N(_02231_),
    .B(_02223_),
    .Y(_02232_));
 sky130_fd_sc_hd__xnor2_4 _09141_ (.A(_02223_),
    .B(_02231_),
    .Y(_02233_));
 sky130_fd_sc_hd__and2_1 _09142_ (.A(_02222_),
    .B(_02233_),
    .X(_02234_));
 sky130_fd_sc_hd__xor2_4 _09143_ (.A(_02222_),
    .B(_02233_),
    .X(_02235_));
 sky130_fd_sc_hd__xnor2_4 _09144_ (.A(_02138_),
    .B(_02235_),
    .Y(_02236_));
 sky130_fd_sc_hd__and2_1 _09145_ (.A(_02137_),
    .B(_02236_),
    .X(_02237_));
 sky130_fd_sc_hd__xnor2_4 _09146_ (.A(_02137_),
    .B(_02236_),
    .Y(_02238_));
 sky130_fd_sc_hd__xnor2_2 _09147_ (.A(_02136_),
    .B(_02238_),
    .Y(_02239_));
 sky130_fd_sc_hd__a21oi_1 _09148_ (.A1(net163),
    .A2(_02132_),
    .B1(_02239_),
    .Y(_02240_));
 sky130_fd_sc_hd__nor2_4 _09149_ (.A(_06455_),
    .B(_06461_),
    .Y(_02241_));
 sky130_fd_sc_hd__or2_4 _09150_ (.A(_06455_),
    .B(_06461_),
    .X(_02242_));
 sky130_fd_sc_hd__a31o_1 _09151_ (.A1(net163),
    .A2(_02132_),
    .A3(_02239_),
    .B1(_02242_),
    .X(_02243_));
 sky130_fd_sc_hd__nor2_2 _09152_ (.A(net285),
    .B(_06480_),
    .Y(_02244_));
 sky130_fd_sc_hd__nand2_1 _09153_ (.A(net294),
    .B(_06479_),
    .Y(_02245_));
 sky130_fd_sc_hd__mux2_1 _09154_ (.A0(net289),
    .A1(reg1_val[30]),
    .S(net178),
    .X(_02246_));
 sky130_fd_sc_hd__mux2_1 _09155_ (.A0(net293),
    .A1(reg1_val[31]),
    .S(net178),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _09156_ (.A0(_02246_),
    .A1(_02247_),
    .S(net216),
    .X(_02248_));
 sky130_fd_sc_hd__mux2_1 _09157_ (.A0(reg1_val[2]),
    .A1(reg1_val[29]),
    .S(net178),
    .X(_02249_));
 sky130_fd_sc_hd__mux2_1 _09158_ (.A0(reg1_val[3]),
    .A1(reg1_val[28]),
    .S(net178),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _09159_ (.A0(_02249_),
    .A1(_02250_),
    .S(net212),
    .X(_02251_));
 sky130_fd_sc_hd__mux2_1 _09160_ (.A0(_02248_),
    .A1(_02251_),
    .S(net218),
    .X(_02252_));
 sky130_fd_sc_hd__mux2_1 _09161_ (.A0(reg1_val[4]),
    .A1(reg1_val[27]),
    .S(net178),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _09162_ (.A0(reg1_val[5]),
    .A1(reg1_val[26]),
    .S(net178),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _09163_ (.A0(_02253_),
    .A1(_02254_),
    .S(net212),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _09164_ (.A0(reg1_val[6]),
    .A1(reg1_val[25]),
    .S(net178),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _09165_ (.A0(reg1_val[7]),
    .A1(reg1_val[24]),
    .S(net178),
    .X(_02257_));
 sky130_fd_sc_hd__mux2_1 _09166_ (.A0(_02256_),
    .A1(_02257_),
    .S(net212),
    .X(_02258_));
 sky130_fd_sc_hd__mux2_1 _09167_ (.A0(_02255_),
    .A1(_02258_),
    .S(net217),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _09168_ (.A0(_02252_),
    .A1(_02259_),
    .S(net220),
    .X(_02260_));
 sky130_fd_sc_hd__mux2_1 _09169_ (.A0(reg1_val[8]),
    .A1(reg1_val[23]),
    .S(net178),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _09170_ (.A0(reg1_val[9]),
    .A1(reg1_val[22]),
    .S(net178),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _09171_ (.A0(_02261_),
    .A1(_02262_),
    .S(net212),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _09172_ (.A0(reg1_val[10]),
    .A1(reg1_val[21]),
    .S(net178),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _09173_ (.A0(reg1_val[11]),
    .A1(reg1_val[20]),
    .S(net178),
    .X(_02265_));
 sky130_fd_sc_hd__mux2_1 _09174_ (.A0(_02264_),
    .A1(_02265_),
    .S(net211),
    .X(_02266_));
 sky130_fd_sc_hd__mux2_1 _09175_ (.A0(_02263_),
    .A1(_02266_),
    .S(net217),
    .X(_02267_));
 sky130_fd_sc_hd__mux2_1 _09176_ (.A0(reg1_val[12]),
    .A1(reg1_val[19]),
    .S(net178),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _09177_ (.A0(reg1_val[13]),
    .A1(reg1_val[18]),
    .S(net178),
    .X(_02269_));
 sky130_fd_sc_hd__mux2_1 _09178_ (.A0(_02268_),
    .A1(_02269_),
    .S(net211),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_1 _09179_ (.A0(net291),
    .A1(reg1_val[17]),
    .S(net178),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _09180_ (.A0(net290),
    .A1(reg1_val[16]),
    .S(net178),
    .X(_02272_));
 sky130_fd_sc_hd__mux2_1 _09181_ (.A0(_02271_),
    .A1(_02272_),
    .S(net211),
    .X(_02273_));
 sky130_fd_sc_hd__mux2_1 _09182_ (.A0(_02270_),
    .A1(_02273_),
    .S(net217),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _09183_ (.A0(_02267_),
    .A1(_02274_),
    .S(net219),
    .X(_02275_));
 sky130_fd_sc_hd__mux2_1 _09184_ (.A0(_02260_),
    .A1(_02275_),
    .S(net222),
    .X(_02276_));
 sky130_fd_sc_hd__mux2_1 _09185_ (.A0(reg1_val[7]),
    .A1(reg1_val[24]),
    .S(net176),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _09186_ (.A0(reg1_val[6]),
    .A1(reg1_val[25]),
    .S(net176),
    .X(_02278_));
 sky130_fd_sc_hd__mux2_1 _09187_ (.A0(_02277_),
    .A1(_02278_),
    .S(net211),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_1 _09188_ (.A0(reg1_val[5]),
    .A1(reg1_val[26]),
    .S(net176),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _09189_ (.A0(reg1_val[4]),
    .A1(reg1_val[27]),
    .S(net176),
    .X(_02281_));
 sky130_fd_sc_hd__mux2_1 _09190_ (.A0(_02280_),
    .A1(_02281_),
    .S(net212),
    .X(_02282_));
 sky130_fd_sc_hd__mux2_1 _09191_ (.A0(_02279_),
    .A1(_02282_),
    .S(net218),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _09192_ (.A0(reg1_val[3]),
    .A1(reg1_val[28]),
    .S(net176),
    .X(_02284_));
 sky130_fd_sc_hd__mux2_1 _09193_ (.A0(reg1_val[2]),
    .A1(reg1_val[29]),
    .S(net176),
    .X(_02285_));
 sky130_fd_sc_hd__mux2_1 _09194_ (.A0(_02284_),
    .A1(_02285_),
    .S(net213),
    .X(_02286_));
 sky130_fd_sc_hd__mux2_1 _09195_ (.A0(net289),
    .A1(reg1_val[30]),
    .S(net176),
    .X(_02287_));
 sky130_fd_sc_hd__mux2_1 _09196_ (.A0(net293),
    .A1(reg1_val[31]),
    .S(net176),
    .X(_02288_));
 sky130_fd_sc_hd__mux2_1 _09197_ (.A0(_02287_),
    .A1(_02288_),
    .S(net213),
    .X(_02289_));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(_02286_),
    .A1(_02289_),
    .S(net218),
    .X(_02290_));
 sky130_fd_sc_hd__mux2_1 _09199_ (.A0(_02283_),
    .A1(_02290_),
    .S(net219),
    .X(_02291_));
 sky130_fd_sc_hd__mux2_1 _09200_ (.A0(net290),
    .A1(reg1_val[16]),
    .S(net176),
    .X(_02292_));
 sky130_fd_sc_hd__mux2_1 _09201_ (.A0(net291),
    .A1(reg1_val[17]),
    .S(net176),
    .X(_02293_));
 sky130_fd_sc_hd__mux2_1 _09202_ (.A0(_02292_),
    .A1(_02293_),
    .S(net211),
    .X(_02294_));
 sky130_fd_sc_hd__mux2_1 _09203_ (.A0(reg1_val[13]),
    .A1(reg1_val[18]),
    .S(net176),
    .X(_02295_));
 sky130_fd_sc_hd__mux2_1 _09204_ (.A0(reg1_val[12]),
    .A1(reg1_val[19]),
    .S(net176),
    .X(_02296_));
 sky130_fd_sc_hd__mux2_1 _09205_ (.A0(_02295_),
    .A1(_02296_),
    .S(net211),
    .X(_02297_));
 sky130_fd_sc_hd__mux2_1 _09206_ (.A0(_02294_),
    .A1(_02297_),
    .S(net217),
    .X(_02298_));
 sky130_fd_sc_hd__mux2_1 _09207_ (.A0(reg1_val[11]),
    .A1(reg1_val[20]),
    .S(net176),
    .X(_02299_));
 sky130_fd_sc_hd__mux2_1 _09208_ (.A0(reg1_val[10]),
    .A1(reg1_val[21]),
    .S(net176),
    .X(_02300_));
 sky130_fd_sc_hd__mux2_1 _09209_ (.A0(_02299_),
    .A1(_02300_),
    .S(net211),
    .X(_02301_));
 sky130_fd_sc_hd__mux2_1 _09210_ (.A0(reg1_val[9]),
    .A1(reg1_val[22]),
    .S(net176),
    .X(_02302_));
 sky130_fd_sc_hd__mux2_1 _09211_ (.A0(reg1_val[8]),
    .A1(reg1_val[23]),
    .S(net176),
    .X(_02303_));
 sky130_fd_sc_hd__mux2_1 _09212_ (.A0(_02302_),
    .A1(_02303_),
    .S(net211),
    .X(_02304_));
 sky130_fd_sc_hd__mux2_1 _09213_ (.A0(_02301_),
    .A1(_02304_),
    .S(net217),
    .X(_02305_));
 sky130_fd_sc_hd__mux2_1 _09214_ (.A0(_02298_),
    .A1(_02305_),
    .S(net219),
    .X(_02306_));
 sky130_fd_sc_hd__mux2_1 _09215_ (.A0(_02291_),
    .A1(_02306_),
    .S(net224),
    .X(_02307_));
 sky130_fd_sc_hd__mux2_2 _09216_ (.A0(_02276_),
    .A1(_02307_),
    .S(net226),
    .X(_02308_));
 sky130_fd_sc_hd__nand2_1 _09217_ (.A(net293),
    .B(curr_PC[0]),
    .Y(_02309_));
 sky130_fd_sc_hd__or2_1 _09218_ (.A(net293),
    .B(curr_PC[0]),
    .X(_02310_));
 sky130_fd_sc_hd__a21o_1 _09219_ (.A1(_02309_),
    .A2(_02310_),
    .B1(net229),
    .X(_02311_));
 sky130_fd_sc_hd__o211a_1 _09220_ (.A1(net249),
    .A2(_02308_),
    .B1(_02311_),
    .C1(net210),
    .X(_02312_));
 sky130_fd_sc_hd__nor2_8 _09221_ (.A(net295),
    .B(_06480_),
    .Y(_02313_));
 sky130_fd_sc_hd__nand2_8 _09222_ (.A(net284),
    .B(_06479_),
    .Y(_02314_));
 sky130_fd_sc_hd__nor2_4 _09223_ (.A(_06478_),
    .B(_06486_),
    .Y(_02315_));
 sky130_fd_sc_hd__or2_1 _09224_ (.A(_06478_),
    .B(_06486_),
    .X(_02316_));
 sky130_fd_sc_hd__nor2_8 _09225_ (.A(_06440_),
    .B(_06477_),
    .Y(_02317_));
 sky130_fd_sc_hd__or2_1 _09226_ (.A(_06440_),
    .B(_06477_),
    .X(_02318_));
 sky130_fd_sc_hd__nor2_4 _09227_ (.A(_06453_),
    .B(_06486_),
    .Y(_02319_));
 sky130_fd_sc_hd__or2_4 _09228_ (.A(_06453_),
    .B(_06486_),
    .X(_02320_));
 sky130_fd_sc_hd__a21o_1 _09229_ (.A1(net236),
    .A2(net197),
    .B1(_06441_),
    .X(_02321_));
 sky130_fd_sc_hd__a21oi_1 _09230_ (.A1(net199),
    .A2(_02321_),
    .B1(_06442_),
    .Y(_02322_));
 sky130_fd_sc_hd__nor2_8 _09231_ (.A(_06440_),
    .B(_06461_),
    .Y(_02323_));
 sky130_fd_sc_hd__or2_4 _09232_ (.A(_06440_),
    .B(_06461_),
    .X(_02324_));
 sky130_fd_sc_hd__and3b_4 _09233_ (.A_N(_06455_),
    .B(_04487_),
    .C(instruction[5]),
    .X(_02325_));
 sky130_fd_sc_hd__or3_4 _09234_ (.A(instruction[6]),
    .B(_04498_),
    .C(_06455_),
    .X(_02326_));
 sky130_fd_sc_hd__o21a_1 _09235_ (.A1(_02323_),
    .A2(_02325_),
    .B1(_06441_),
    .X(_02327_));
 sky130_fd_sc_hd__nor2_1 _09236_ (.A(_06461_),
    .B(_06478_),
    .Y(_02328_));
 sky130_fd_sc_hd__or2_1 _09237_ (.A(_06461_),
    .B(_06478_),
    .X(_02329_));
 sky130_fd_sc_hd__nor2_4 _09238_ (.A(_06453_),
    .B(_06461_),
    .Y(_02330_));
 sky130_fd_sc_hd__or2_1 _09239_ (.A(_06453_),
    .B(_06461_),
    .X(_02331_));
 sky130_fd_sc_hd__a221o_1 _09240_ (.A1(\div_res[0] ),
    .A2(_02328_),
    .B1(_02330_),
    .B2(\div_shifter[32] ),
    .C1(_02327_),
    .X(_02332_));
 sky130_fd_sc_hd__or2_1 _09241_ (.A(_02322_),
    .B(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__nor2_2 _09242_ (.A(_04531_),
    .B(_06476_),
    .Y(_02334_));
 sky130_fd_sc_hd__or2_4 _09243_ (.A(net225),
    .B(_02334_),
    .X(_02335_));
 sky130_fd_sc_hd__mux2_1 _09244_ (.A0(_02288_),
    .A1(_02334_),
    .S(net213),
    .X(_02336_));
 sky130_fd_sc_hd__o21ai_1 _09245_ (.A1(_06359_),
    .A2(_02334_),
    .B1(_02336_),
    .Y(_02337_));
 sky130_fd_sc_hd__inv_2 _09246_ (.A(_02337_),
    .Y(_02338_));
 sky130_fd_sc_hd__or2_1 _09247_ (.A(_06352_),
    .B(_02334_),
    .X(_02339_));
 sky130_fd_sc_hd__and2_1 _09248_ (.A(_02338_),
    .B(_02339_),
    .X(_02340_));
 sky130_fd_sc_hd__nor2_1 _09249_ (.A(net224),
    .B(_02334_),
    .Y(_02341_));
 sky130_fd_sc_hd__or2_2 _09250_ (.A(net224),
    .B(_02334_),
    .X(_02342_));
 sky130_fd_sc_hd__nand3_2 _09251_ (.A(_02335_),
    .B(_02340_),
    .C(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__inv_2 _09252_ (.A(_02343_),
    .Y(_02344_));
 sky130_fd_sc_hd__a221o_1 _09253_ (.A1(_02308_),
    .A2(_02313_),
    .B1(_02344_),
    .B2(net179),
    .C1(_02333_),
    .X(_02345_));
 sky130_fd_sc_hd__a311o_1 _09254_ (.A1(_04498_),
    .A2(_06429_),
    .A3(_06454_),
    .B1(_02312_),
    .C1(_02345_),
    .X(_02346_));
 sky130_fd_sc_hd__a41o_1 _09255_ (.A1(_04487_),
    .A2(instruction[5]),
    .A3(_06437_),
    .A4(_06439_),
    .B1(_02346_),
    .X(_02347_));
 sky130_fd_sc_hd__o21ba_1 _09256_ (.A1(_02240_),
    .A2(_02243_),
    .B1_N(_02347_),
    .X(_02348_));
 sky130_fd_sc_hd__mux2_2 _09257_ (.A0(net216),
    .A1(_02348_),
    .S(net209),
    .X(_02349_));
 sky130_fd_sc_hd__or2_1 _09258_ (.A(curr_PC[0]),
    .B(net242),
    .X(_02350_));
 sky130_fd_sc_hd__o21ai_4 _09259_ (.A1(net248),
    .A2(_02349_),
    .B1(_02350_),
    .Y(dest_val[0]));
 sky130_fd_sc_hd__xor2_1 _09260_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .X(_02351_));
 sky130_fd_sc_hd__or2_2 _09261_ (.A(_02132_),
    .B(_02239_),
    .X(_02352_));
 sky130_fd_sc_hd__a21oi_4 _09262_ (.A1(_02138_),
    .A2(_02235_),
    .B1(_02234_),
    .Y(_02353_));
 sky130_fd_sc_hd__o21ai_4 _09263_ (.A1(_02229_),
    .A2(_02230_),
    .B1(_02232_),
    .Y(_02354_));
 sky130_fd_sc_hd__a32o_1 _09264_ (.A1(_02180_),
    .A2(_02181_),
    .A3(_02192_),
    .B1(_02193_),
    .B2(_02171_),
    .X(_02355_));
 sky130_fd_sc_hd__o22a_1 _09265_ (.A1(net130),
    .A2(net24),
    .B1(net16),
    .B2(net128),
    .X(_02356_));
 sky130_fd_sc_hd__xnor2_1 _09266_ (.A(net71),
    .B(_02356_),
    .Y(_02357_));
 sky130_fd_sc_hd__a22o_1 _09267_ (.A1(net37),
    .A2(_00308_),
    .B1(_00330_),
    .B2(net39),
    .X(_02358_));
 sky130_fd_sc_hd__xor2_1 _09268_ (.A(net91),
    .B(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__and2b_1 _09269_ (.A_N(_02357_),
    .B(_02359_),
    .X(_02360_));
 sky130_fd_sc_hd__and2b_1 _09270_ (.A_N(_02359_),
    .B(_02357_),
    .X(_02361_));
 sky130_fd_sc_hd__or2_1 _09271_ (.A(_02360_),
    .B(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__a22o_1 _09272_ (.A1(net44),
    .A2(net113),
    .B1(_00374_),
    .B2(net42),
    .X(_02363_));
 sky130_fd_sc_hd__xor2_1 _09273_ (.A(net94),
    .B(_02363_),
    .X(_02364_));
 sky130_fd_sc_hd__and2b_1 _09274_ (.A_N(_02362_),
    .B(_02364_),
    .X(_02365_));
 sky130_fd_sc_hd__and2b_1 _09275_ (.A_N(_02364_),
    .B(_02362_),
    .X(_02366_));
 sky130_fd_sc_hd__or2_1 _09276_ (.A(_02365_),
    .B(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__a21oi_1 _09277_ (.A1(_02157_),
    .A2(_02160_),
    .B1(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hd__and3_1 _09278_ (.A(_02157_),
    .B(_02160_),
    .C(_02367_),
    .X(_02369_));
 sky130_fd_sc_hd__nor2_1 _09279_ (.A(_02368_),
    .B(_02369_),
    .Y(_02370_));
 sky130_fd_sc_hd__xnor2_1 _09280_ (.A(_02355_),
    .B(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__and2b_1 _09281_ (.A_N(_02176_),
    .B(_02180_),
    .X(_02372_));
 sky130_fd_sc_hd__a21o_1 _09282_ (.A1(_02211_),
    .A2(_02213_),
    .B1(_02210_),
    .X(_02373_));
 sky130_fd_sc_hd__a21o_1 _09283_ (.A1(_02167_),
    .A2(_02170_),
    .B1(_02166_),
    .X(_02374_));
 sky130_fd_sc_hd__xor2_1 _09284_ (.A(_02373_),
    .B(_02374_),
    .X(_02375_));
 sky130_fd_sc_hd__and2b_1 _09285_ (.A_N(_02372_),
    .B(_02375_),
    .X(_02376_));
 sky130_fd_sc_hd__xnor2_1 _09286_ (.A(_02372_),
    .B(_02375_),
    .Y(_02377_));
 sky130_fd_sc_hd__o22a_1 _09287_ (.A1(net56),
    .A2(net148),
    .B1(net146),
    .B2(net68),
    .X(_02378_));
 sky130_fd_sc_hd__xnor2_1 _09288_ (.A(net202),
    .B(_02378_),
    .Y(_02379_));
 sky130_fd_sc_hd__o22a_1 _09289_ (.A1(net57),
    .A2(net106),
    .B1(net104),
    .B2(net63),
    .X(_02380_));
 sky130_fd_sc_hd__xnor2_1 _09290_ (.A(net135),
    .B(_02380_),
    .Y(_02381_));
 sky130_fd_sc_hd__nor2_1 _09291_ (.A(_02379_),
    .B(_02381_),
    .Y(_02382_));
 sky130_fd_sc_hd__xor2_1 _09292_ (.A(_02379_),
    .B(_02381_),
    .X(_02383_));
 sky130_fd_sc_hd__o22a_1 _09293_ (.A1(net65),
    .A2(_00184_),
    .B1(net132),
    .B2(net59),
    .X(_02384_));
 sky130_fd_sc_hd__xnor2_1 _09294_ (.A(net181),
    .B(_02384_),
    .Y(_02385_));
 sky130_fd_sc_hd__and2b_1 _09295_ (.A_N(_02385_),
    .B(_02383_),
    .X(_02386_));
 sky130_fd_sc_hd__and2b_1 _09296_ (.A_N(_02383_),
    .B(_02385_),
    .X(_02387_));
 sky130_fd_sc_hd__nor2_1 _09297_ (.A(_02386_),
    .B(_02387_),
    .Y(_02388_));
 sky130_fd_sc_hd__o22a_1 _09298_ (.A1(net150),
    .A2(net13),
    .B1(net8),
    .B2(net152),
    .X(_02389_));
 sky130_fd_sc_hd__xor2_1 _09299_ (.A(net205),
    .B(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__a21o_1 _09300_ (.A1(_00697_),
    .A2(_00698_),
    .B1(net156),
    .X(_02391_));
 sky130_fd_sc_hd__or3_1 _09301_ (.A(net154),
    .B(_00405_),
    .C(_00407_),
    .X(_02392_));
 sky130_fd_sc_hd__nand3_1 _09302_ (.A(_06532_),
    .B(_02391_),
    .C(_02392_),
    .Y(_02393_));
 sky130_fd_sc_hd__a21o_1 _09303_ (.A1(_02391_),
    .A2(_02392_),
    .B1(_06532_),
    .X(_02394_));
 sky130_fd_sc_hd__a21oi_1 _09304_ (.A1(_02393_),
    .A2(_02394_),
    .B1(net239),
    .Y(_02395_));
 sky130_fd_sc_hd__a21o_1 _09305_ (.A1(_02393_),
    .A2(_02394_),
    .B1(net239),
    .X(_02396_));
 sky130_fd_sc_hd__nand3_1 _09306_ (.A(net239),
    .B(_02393_),
    .C(_02394_),
    .Y(_02397_));
 sky130_fd_sc_hd__and3_1 _09307_ (.A(_02390_),
    .B(_02396_),
    .C(_02397_),
    .X(_02398_));
 sky130_fd_sc_hd__a21oi_1 _09308_ (.A1(_02396_),
    .A2(_02397_),
    .B1(_02390_),
    .Y(_02399_));
 sky130_fd_sc_hd__nor2_2 _09309_ (.A(_02398_),
    .B(_02399_),
    .Y(_02400_));
 sky130_fd_sc_hd__o22a_1 _09310_ (.A1(net61),
    .A2(net86),
    .B1(net82),
    .B2(net53),
    .X(_02401_));
 sky130_fd_sc_hd__xnor2_1 _09311_ (.A(net137),
    .B(_02401_),
    .Y(_02402_));
 sky130_fd_sc_hd__o22a_1 _09312_ (.A1(net98),
    .A2(net35),
    .B1(net33),
    .B2(net84),
    .X(_02403_));
 sky130_fd_sc_hd__xnor2_1 _09313_ (.A(net124),
    .B(_02403_),
    .Y(_02404_));
 sky130_fd_sc_hd__or2_1 _09314_ (.A(_02402_),
    .B(_02404_),
    .X(_02405_));
 sky130_fd_sc_hd__nand2_1 _09315_ (.A(_02402_),
    .B(_02404_),
    .Y(_02406_));
 sky130_fd_sc_hd__nand2_1 _09316_ (.A(_02405_),
    .B(_02406_),
    .Y(_02407_));
 sky130_fd_sc_hd__o22a_1 _09317_ (.A1(net51),
    .A2(net78),
    .B1(net74),
    .B2(net100),
    .X(_02408_));
 sky130_fd_sc_hd__xnor2_2 _09318_ (.A(net121),
    .B(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__xor2_2 _09319_ (.A(_02407_),
    .B(_02409_),
    .X(_02410_));
 sky130_fd_sc_hd__nand2_1 _09320_ (.A(_02400_),
    .B(_02410_),
    .Y(_02411_));
 sky130_fd_sc_hd__xor2_2 _09321_ (.A(_02400_),
    .B(_02410_),
    .X(_02412_));
 sky130_fd_sc_hd__and2_1 _09322_ (.A(_02388_),
    .B(_02412_),
    .X(_02413_));
 sky130_fd_sc_hd__inv_2 _09323_ (.A(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__xnor2_2 _09324_ (.A(_02388_),
    .B(_02412_),
    .Y(_02415_));
 sky130_fd_sc_hd__nor2_1 _09325_ (.A(net144),
    .B(net21),
    .Y(_02416_));
 sky130_fd_sc_hd__o22a_1 _09326_ (.A1(net142),
    .A2(net11),
    .B1(net6),
    .B2(net140),
    .X(_02417_));
 sky130_fd_sc_hd__xnor2_1 _09327_ (.A(net21),
    .B(_02417_),
    .Y(_02418_));
 sky130_fd_sc_hd__a21oi_1 _09328_ (.A1(_02188_),
    .A2(_02190_),
    .B1(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__a21o_1 _09329_ (.A1(_02188_),
    .A2(_02190_),
    .B1(_02418_),
    .X(_02420_));
 sky130_fd_sc_hd__and3_1 _09330_ (.A(_02188_),
    .B(_02190_),
    .C(_02418_),
    .X(_02421_));
 sky130_fd_sc_hd__nor2_1 _09331_ (.A(_02419_),
    .B(_02421_),
    .Y(_02422_));
 sky130_fd_sc_hd__xnor2_2 _09332_ (.A(_02416_),
    .B(_02422_),
    .Y(_02423_));
 sky130_fd_sc_hd__or2_1 _09333_ (.A(_02415_),
    .B(_02423_),
    .X(_02424_));
 sky130_fd_sc_hd__nand2_1 _09334_ (.A(_02415_),
    .B(_02423_),
    .Y(_02425_));
 sky130_fd_sc_hd__xnor2_1 _09335_ (.A(_02415_),
    .B(_02423_),
    .Y(_02426_));
 sky130_fd_sc_hd__xnor2_1 _09336_ (.A(_02377_),
    .B(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__a21o_1 _09337_ (.A1(_02142_),
    .A2(_02144_),
    .B1(_02148_),
    .X(_02428_));
 sky130_fd_sc_hd__o22a_1 _09338_ (.A1(net48),
    .A2(_00290_),
    .B1(net112),
    .B2(net46),
    .X(_02429_));
 sky130_fd_sc_hd__xnor2_1 _09339_ (.A(net97),
    .B(_02429_),
    .Y(_02430_));
 sky130_fd_sc_hd__o22a_1 _09340_ (.A1(net27),
    .A2(net81),
    .B1(net77),
    .B2(net25),
    .X(_02431_));
 sky130_fd_sc_hd__xnor2_1 _09341_ (.A(net88),
    .B(_02431_),
    .Y(_02432_));
 sky130_fd_sc_hd__and2_1 _09342_ (.A(_02430_),
    .B(_02432_),
    .X(_02433_));
 sky130_fd_sc_hd__nor2_1 _09343_ (.A(_02430_),
    .B(_02432_),
    .Y(_02434_));
 sky130_fd_sc_hd__nor2_1 _09344_ (.A(_02433_),
    .B(_02434_),
    .Y(_02435_));
 sky130_fd_sc_hd__a22o_1 _09345_ (.A1(net118),
    .A2(net29),
    .B1(_00366_),
    .B2(net31),
    .X(_02436_));
 sky130_fd_sc_hd__xnor2_1 _09346_ (.A(net50),
    .B(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__xnor2_1 _09347_ (.A(_02435_),
    .B(_02437_),
    .Y(_02438_));
 sky130_fd_sc_hd__a21boi_2 _09348_ (.A1(_02195_),
    .A2(_02200_),
    .B1_N(_02199_),
    .Y(_02439_));
 sky130_fd_sc_hd__nor2_1 _09349_ (.A(_02438_),
    .B(_02439_),
    .Y(_02440_));
 sky130_fd_sc_hd__xor2_1 _09350_ (.A(_02438_),
    .B(_02439_),
    .X(_02441_));
 sky130_fd_sc_hd__xor2_1 _09351_ (.A(_02428_),
    .B(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__xnor2_1 _09352_ (.A(_02427_),
    .B(_02442_),
    .Y(_02443_));
 sky130_fd_sc_hd__nor2_1 _09353_ (.A(_02371_),
    .B(_02443_),
    .Y(_02444_));
 sky130_fd_sc_hd__and2_1 _09354_ (.A(_02371_),
    .B(_02443_),
    .X(_02445_));
 sky130_fd_sc_hd__nor2_2 _09355_ (.A(_02444_),
    .B(_02445_),
    .Y(_02446_));
 sky130_fd_sc_hd__a21o_2 _09356_ (.A1(_02155_),
    .A2(_02220_),
    .B1(_02219_),
    .X(_02447_));
 sky130_fd_sc_hd__nand2_2 _09357_ (.A(_02151_),
    .B(_02154_),
    .Y(_02448_));
 sky130_fd_sc_hd__a21oi_4 _09358_ (.A1(_02161_),
    .A2(_02203_),
    .B1(_02202_),
    .Y(_02449_));
 sky130_fd_sc_hd__a21oi_2 _09359_ (.A1(_02205_),
    .A2(_02217_),
    .B1(_02216_),
    .Y(_02450_));
 sky130_fd_sc_hd__nor2_1 _09360_ (.A(_02449_),
    .B(_02450_),
    .Y(_02451_));
 sky130_fd_sc_hd__xor2_4 _09361_ (.A(_02449_),
    .B(_02450_),
    .X(_02452_));
 sky130_fd_sc_hd__xnor2_4 _09362_ (.A(_02448_),
    .B(_02452_),
    .Y(_02453_));
 sky130_fd_sc_hd__a21oi_4 _09363_ (.A1(_02224_),
    .A2(_02228_),
    .B1(_02227_),
    .Y(_02454_));
 sky130_fd_sc_hd__xnor2_4 _09364_ (.A(_02453_),
    .B(_02454_),
    .Y(_02455_));
 sky130_fd_sc_hd__nand2b_1 _09365_ (.A_N(_02455_),
    .B(_02447_),
    .Y(_02456_));
 sky130_fd_sc_hd__xnor2_4 _09366_ (.A(_02447_),
    .B(_02455_),
    .Y(_02457_));
 sky130_fd_sc_hd__and2_1 _09367_ (.A(_02446_),
    .B(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__xor2_4 _09368_ (.A(_02446_),
    .B(_02457_),
    .X(_02459_));
 sky130_fd_sc_hd__xnor2_4 _09369_ (.A(_02354_),
    .B(_02459_),
    .Y(_02460_));
 sky130_fd_sc_hd__or2_1 _09370_ (.A(_02353_),
    .B(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__xnor2_4 _09371_ (.A(_02353_),
    .B(_02460_),
    .Y(_02462_));
 sky130_fd_sc_hd__or4b_2 _09372_ (.A(_02126_),
    .B(_02129_),
    .C(_02238_),
    .D_N(_01801_),
    .X(_02463_));
 sky130_fd_sc_hd__o2bb2a_1 _09373_ (.A1_N(_02017_),
    .A2_N(_02124_),
    .B1(_02137_),
    .B2(_02236_),
    .X(_02464_));
 sky130_fd_sc_hd__o32a_2 _09374_ (.A1(_02126_),
    .A2(_02127_),
    .A3(_02238_),
    .B1(_02464_),
    .B2(_02237_),
    .X(_02465_));
 sky130_fd_sc_hd__nand2_4 _09375_ (.A(_02463_),
    .B(_02465_),
    .Y(_02466_));
 sky130_fd_sc_hd__xnor2_4 _09376_ (.A(_02462_),
    .B(_02466_),
    .Y(_02467_));
 sky130_fd_sc_hd__a21oi_1 _09377_ (.A1(net163),
    .A2(_02352_),
    .B1(_02467_),
    .Y(_02468_));
 sky130_fd_sc_hd__a31o_1 _09378_ (.A1(net163),
    .A2(_02352_),
    .A3(_02467_),
    .B1(_02242_),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _09379_ (.A0(_02246_),
    .A1(_02249_),
    .S(net212),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _09380_ (.A0(_02250_),
    .A1(_02253_),
    .S(net212),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _09381_ (.A0(_02470_),
    .A1(_02471_),
    .S(net218),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _09382_ (.A0(_02254_),
    .A1(_02256_),
    .S(net212),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _09383_ (.A0(_02257_),
    .A1(_02261_),
    .S(net212),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _09384_ (.A0(_02473_),
    .A1(_02474_),
    .S(net218),
    .X(_02475_));
 sky130_fd_sc_hd__mux2_1 _09385_ (.A0(_02472_),
    .A1(_02475_),
    .S(net220),
    .X(_02476_));
 sky130_fd_sc_hd__mux2_1 _09386_ (.A0(_02262_),
    .A1(_02264_),
    .S(net211),
    .X(_02477_));
 sky130_fd_sc_hd__mux2_1 _09387_ (.A0(_02265_),
    .A1(_02268_),
    .S(net211),
    .X(_02478_));
 sky130_fd_sc_hd__mux2_1 _09388_ (.A0(_02477_),
    .A1(_02478_),
    .S(net217),
    .X(_02479_));
 sky130_fd_sc_hd__mux2_1 _09389_ (.A0(_02269_),
    .A1(_02271_),
    .S(net211),
    .X(_02480_));
 sky130_fd_sc_hd__mux2_1 _09390_ (.A0(_02272_),
    .A1(_02292_),
    .S(net211),
    .X(_02481_));
 sky130_fd_sc_hd__mux2_1 _09391_ (.A0(_02480_),
    .A1(_02481_),
    .S(net217),
    .X(_02482_));
 sky130_fd_sc_hd__mux2_1 _09392_ (.A0(_02479_),
    .A1(_02482_),
    .S(net220),
    .X(_02483_));
 sky130_fd_sc_hd__mux2_1 _09393_ (.A0(_02476_),
    .A1(_02483_),
    .S(net223),
    .X(_02484_));
 sky130_fd_sc_hd__mux2_1 _09394_ (.A0(_02278_),
    .A1(_02280_),
    .S(net211),
    .X(_02485_));
 sky130_fd_sc_hd__mux2_1 _09395_ (.A0(_02281_),
    .A1(_02284_),
    .S(net213),
    .X(_02486_));
 sky130_fd_sc_hd__mux2_1 _09396_ (.A0(_02485_),
    .A1(_02486_),
    .S(net218),
    .X(_02487_));
 sky130_fd_sc_hd__mux2_1 _09397_ (.A0(_02285_),
    .A1(_02287_),
    .S(net213),
    .X(_02488_));
 sky130_fd_sc_hd__mux2_1 _09398_ (.A0(_02336_),
    .A1(_02488_),
    .S(_06359_),
    .X(_02489_));
 sky130_fd_sc_hd__mux2_1 _09399_ (.A0(_02487_),
    .A1(_02489_),
    .S(net219),
    .X(_02490_));
 sky130_fd_sc_hd__mux2_1 _09400_ (.A0(_02293_),
    .A1(_02295_),
    .S(net211),
    .X(_02491_));
 sky130_fd_sc_hd__mux2_1 _09401_ (.A0(_02296_),
    .A1(_02299_),
    .S(net211),
    .X(_02492_));
 sky130_fd_sc_hd__mux2_1 _09402_ (.A0(_02491_),
    .A1(_02492_),
    .S(net217),
    .X(_02493_));
 sky130_fd_sc_hd__mux2_1 _09403_ (.A0(_02300_),
    .A1(_02302_),
    .S(net211),
    .X(_02494_));
 sky130_fd_sc_hd__mux2_1 _09404_ (.A0(_02277_),
    .A1(_02303_),
    .S(net215),
    .X(_02495_));
 sky130_fd_sc_hd__mux2_1 _09405_ (.A0(_02494_),
    .A1(_02495_),
    .S(net218),
    .X(_02496_));
 sky130_fd_sc_hd__mux2_1 _09406_ (.A0(_02493_),
    .A1(_02496_),
    .S(net220),
    .X(_02497_));
 sky130_fd_sc_hd__mux2_1 _09407_ (.A0(_02490_),
    .A1(_02497_),
    .S(net224),
    .X(_02498_));
 sky130_fd_sc_hd__mux2_1 _09408_ (.A0(_02484_),
    .A1(_02498_),
    .S(net226),
    .X(_02499_));
 sky130_fd_sc_hd__inv_2 _09409_ (.A(_02499_),
    .Y(_02500_));
 sky130_fd_sc_hd__or2_1 _09410_ (.A(net289),
    .B(curr_PC[1]),
    .X(_02501_));
 sky130_fd_sc_hd__nand2_1 _09411_ (.A(net289),
    .B(curr_PC[1]),
    .Y(_02502_));
 sky130_fd_sc_hd__nand2_1 _09412_ (.A(_02501_),
    .B(_02502_),
    .Y(_02503_));
 sky130_fd_sc_hd__xnor2_1 _09413_ (.A(_02309_),
    .B(_02503_),
    .Y(_02504_));
 sky130_fd_sc_hd__a21o_1 _09414_ (.A1(net249),
    .A2(_02504_),
    .B1(_06476_),
    .X(_02505_));
 sky130_fd_sc_hd__a21oi_1 _09415_ (.A1(_02314_),
    .A2(_02505_),
    .B1(_02500_),
    .Y(_02506_));
 sky130_fd_sc_hd__a21oi_1 _09416_ (.A1(\div_res[0] ),
    .A2(net162),
    .B1(\div_res[1] ),
    .Y(_02507_));
 sky130_fd_sc_hd__a311o_1 _09417_ (.A1(\div_res[1] ),
    .A2(\div_res[0] ),
    .A3(net162),
    .B1(net195),
    .C1(_02507_),
    .X(_02508_));
 sky130_fd_sc_hd__xnor2_1 _09418_ (.A(_06362_),
    .B(_06366_),
    .Y(_02509_));
 sky130_fd_sc_hd__nand2_1 _09419_ (.A(net285),
    .B(net213),
    .Y(_02510_));
 sky130_fd_sc_hd__a21oi_1 _09420_ (.A1(_02509_),
    .A2(_02510_),
    .B1(net236),
    .Y(_02511_));
 sky130_fd_sc_hd__o21ai_1 _09421_ (.A1(_02509_),
    .A2(_02510_),
    .B1(_02511_),
    .Y(_02512_));
 sky130_fd_sc_hd__or3b_1 _09422_ (.A(_06359_),
    .B(net196),
    .C_N(net289),
    .X(_02513_));
 sky130_fd_sc_hd__and2_1 _09423_ (.A(divi1_sign),
    .B(net295),
    .X(_02514_));
 sky130_fd_sc_hd__a21oi_1 _09424_ (.A1(\div_shifter[32] ),
    .A2(net235),
    .B1(\div_shifter[33] ),
    .Y(_02515_));
 sky130_fd_sc_hd__and3_1 _09425_ (.A(\div_shifter[33] ),
    .B(\div_shifter[32] ),
    .C(net235),
    .X(_02516_));
 sky130_fd_sc_hd__o32a_1 _09426_ (.A1(net193),
    .A2(_02515_),
    .A3(_02516_),
    .B1(net209),
    .B2(_06359_),
    .X(_02517_));
 sky130_fd_sc_hd__o2bb2a_1 _09427_ (.A1_N(_06361_),
    .A2_N(_02315_),
    .B1(_02505_),
    .B2(net229),
    .X(_02518_));
 sky130_fd_sc_hd__o2111a_1 _09428_ (.A1(_06362_),
    .A2(net197),
    .B1(_02513_),
    .C1(_02517_),
    .D1(_02518_),
    .X(_02519_));
 sky130_fd_sc_hd__and4b_1 _09429_ (.A_N(_02506_),
    .B(_02508_),
    .C(_02512_),
    .D(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__o21ai_1 _09430_ (.A1(net159),
    .A2(_06494_),
    .B1(_06441_),
    .Y(_02521_));
 sky130_fd_sc_hd__a21o_1 _09431_ (.A1(net159),
    .A2(net238),
    .B1(_02521_),
    .X(_02522_));
 sky130_fd_sc_hd__xnor2_1 _09432_ (.A(_01754_),
    .B(_02522_),
    .Y(_02523_));
 sky130_fd_sc_hd__nand2_1 _09433_ (.A(_02323_),
    .B(_02523_),
    .Y(_02524_));
 sky130_fd_sc_hd__mux2_1 _09434_ (.A0(_02289_),
    .A1(_02334_),
    .S(net218),
    .X(_02525_));
 sky130_fd_sc_hd__o21ai_2 _09435_ (.A1(net221),
    .A2(_02525_),
    .B1(_02339_),
    .Y(_02526_));
 sky130_fd_sc_hd__inv_2 _09436_ (.A(_02526_),
    .Y(_02527_));
 sky130_fd_sc_hd__a21oi_2 _09437_ (.A1(net224),
    .A2(_02526_),
    .B1(_02341_),
    .Y(_02528_));
 sky130_fd_sc_hd__o21ai_2 _09438_ (.A1(net227),
    .A2(_02528_),
    .B1(_02335_),
    .Y(_02529_));
 sky130_fd_sc_hd__o211a_1 _09439_ (.A1(net177),
    .A2(_02529_),
    .B1(_02524_),
    .C1(_02520_),
    .X(_02530_));
 sky130_fd_sc_hd__o21ai_2 _09440_ (.A1(_02468_),
    .A2(_02469_),
    .B1(_02530_),
    .Y(_02531_));
 sky130_fd_sc_hd__mux2_8 _09441_ (.A0(_02351_),
    .A1(_02531_),
    .S(net242),
    .X(dest_val[1]));
 sky130_fd_sc_hd__and3_1 _09442_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .C(curr_PC[2]),
    .X(_02532_));
 sky130_fd_sc_hd__a21oi_1 _09443_ (.A1(curr_PC[0]),
    .A2(curr_PC[1]),
    .B1(curr_PC[2]),
    .Y(_02533_));
 sky130_fd_sc_hd__or3_1 _09444_ (.A(net242),
    .B(_02532_),
    .C(_02533_),
    .X(_02534_));
 sky130_fd_sc_hd__o21ai_1 _09445_ (.A1(_02352_),
    .A2(_02467_),
    .B1(net163),
    .Y(_02535_));
 sky130_fd_sc_hd__a21oi_4 _09446_ (.A1(_02354_),
    .A2(_02459_),
    .B1(_02458_),
    .Y(_02536_));
 sky130_fd_sc_hd__o21ai_4 _09447_ (.A1(_02453_),
    .A2(_02454_),
    .B1(_02456_),
    .Y(_02537_));
 sky130_fd_sc_hd__o22a_1 _09448_ (.A1(_00375_),
    .A2(net24),
    .B1(net16),
    .B2(net130),
    .X(_02538_));
 sky130_fd_sc_hd__xnor2_1 _09449_ (.A(net71),
    .B(_02538_),
    .Y(_02539_));
 sky130_fd_sc_hd__a22o_1 _09450_ (.A1(net39),
    .A2(_00324_),
    .B1(_00330_),
    .B2(net37),
    .X(_02540_));
 sky130_fd_sc_hd__xor2_1 _09451_ (.A(net91),
    .B(_02540_),
    .X(_02541_));
 sky130_fd_sc_hd__and2b_1 _09452_ (.A_N(_02539_),
    .B(_02541_),
    .X(_02542_));
 sky130_fd_sc_hd__and2b_1 _09453_ (.A_N(_02541_),
    .B(_02539_),
    .X(_02543_));
 sky130_fd_sc_hd__or2_1 _09454_ (.A(_02542_),
    .B(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__a22o_1 _09455_ (.A1(net44),
    .A2(_00308_),
    .B1(net113),
    .B2(net42),
    .X(_02545_));
 sky130_fd_sc_hd__xor2_1 _09456_ (.A(net94),
    .B(_02545_),
    .X(_02546_));
 sky130_fd_sc_hd__and2b_1 _09457_ (.A_N(_02544_),
    .B(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__and2b_1 _09458_ (.A_N(_02546_),
    .B(_02544_),
    .X(_02548_));
 sky130_fd_sc_hd__or2_2 _09459_ (.A(_02547_),
    .B(_02548_),
    .X(_02549_));
 sky130_fd_sc_hd__a21oi_2 _09460_ (.A1(_02373_),
    .A2(_02374_),
    .B1(_02376_),
    .Y(_02550_));
 sky130_fd_sc_hd__xnor2_1 _09461_ (.A(_02549_),
    .B(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__a21o_1 _09462_ (.A1(_02411_),
    .A2(_02414_),
    .B1(_02551_),
    .X(_02552_));
 sky130_fd_sc_hd__nand3_1 _09463_ (.A(_02411_),
    .B(_02414_),
    .C(_02551_),
    .Y(_02553_));
 sky130_fd_sc_hd__and2_2 _09464_ (.A(_02552_),
    .B(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__o21a_1 _09465_ (.A1(_02407_),
    .A2(_02409_),
    .B1(_02405_),
    .X(_02555_));
 sky130_fd_sc_hd__a21o_1 _09466_ (.A1(_02435_),
    .A2(_02437_),
    .B1(_02433_),
    .X(_02556_));
 sky130_fd_sc_hd__nor2_1 _09467_ (.A(_02382_),
    .B(_02386_),
    .Y(_02557_));
 sky130_fd_sc_hd__o21ai_1 _09468_ (.A1(_02382_),
    .A2(_02386_),
    .B1(_02556_),
    .Y(_02558_));
 sky130_fd_sc_hd__xnor2_1 _09469_ (.A(_02556_),
    .B(_02557_),
    .Y(_02559_));
 sky130_fd_sc_hd__nand2b_1 _09470_ (.A_N(_02555_),
    .B(_02559_),
    .Y(_02560_));
 sky130_fd_sc_hd__xnor2_1 _09471_ (.A(_02555_),
    .B(_02559_),
    .Y(_02561_));
 sky130_fd_sc_hd__nor2_1 _09472_ (.A(net140),
    .B(net21),
    .Y(_02562_));
 sky130_fd_sc_hd__o22a_1 _09473_ (.A1(net128),
    .A2(net11),
    .B1(net6),
    .B2(net142),
    .X(_02563_));
 sky130_fd_sc_hd__xnor2_1 _09474_ (.A(net22),
    .B(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__o21a_1 _09475_ (.A1(_02395_),
    .A2(_02398_),
    .B1(_02564_),
    .X(_02565_));
 sky130_fd_sc_hd__or3_1 _09476_ (.A(_02395_),
    .B(_02398_),
    .C(_02564_),
    .X(_02566_));
 sky130_fd_sc_hd__and2b_1 _09477_ (.A_N(_02565_),
    .B(_02566_),
    .X(_02567_));
 sky130_fd_sc_hd__xnor2_2 _09478_ (.A(_02562_),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__o22a_1 _09479_ (.A1(net59),
    .A2(net106),
    .B1(net105),
    .B2(net57),
    .X(_02569_));
 sky130_fd_sc_hd__xnor2_1 _09480_ (.A(net135),
    .B(_02569_),
    .Y(_02570_));
 sky130_fd_sc_hd__o22a_1 _09481_ (.A1(net56),
    .A2(net146),
    .B1(net17),
    .B2(net148),
    .X(_02571_));
 sky130_fd_sc_hd__xnor2_1 _09482_ (.A(net202),
    .B(_02571_),
    .Y(_02572_));
 sky130_fd_sc_hd__nor2_1 _09483_ (.A(_02570_),
    .B(_02572_),
    .Y(_02573_));
 sky130_fd_sc_hd__and2_1 _09484_ (.A(_02570_),
    .B(_02572_),
    .X(_02574_));
 sky130_fd_sc_hd__nor2_1 _09485_ (.A(_02573_),
    .B(_02574_),
    .Y(_02575_));
 sky130_fd_sc_hd__o22a_1 _09486_ (.A1(net68),
    .A2(net134),
    .B1(net132),
    .B2(net65),
    .X(_02576_));
 sky130_fd_sc_hd__xnor2_1 _09487_ (.A(net181),
    .B(_02576_),
    .Y(_02577_));
 sky130_fd_sc_hd__xnor2_1 _09488_ (.A(_02575_),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__o22a_1 _09489_ (.A1(net63),
    .A2(net86),
    .B1(net82),
    .B2(net61),
    .X(_02579_));
 sky130_fd_sc_hd__xnor2_1 _09490_ (.A(net137),
    .B(_02579_),
    .Y(_02580_));
 sky130_fd_sc_hd__o22a_1 _09491_ (.A1(net100),
    .A2(net35),
    .B1(net33),
    .B2(net98),
    .X(_02581_));
 sky130_fd_sc_hd__xnor2_1 _09492_ (.A(net124),
    .B(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__or2_1 _09493_ (.A(_02580_),
    .B(_02582_),
    .X(_02583_));
 sky130_fd_sc_hd__nand2_1 _09494_ (.A(_02580_),
    .B(_02582_),
    .Y(_02584_));
 sky130_fd_sc_hd__nand2_1 _09495_ (.A(_02583_),
    .B(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__o22a_1 _09496_ (.A1(net53),
    .A2(net78),
    .B1(net74),
    .B2(net51),
    .X(_02586_));
 sky130_fd_sc_hd__xnor2_1 _09497_ (.A(net121),
    .B(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__xnor2_1 _09498_ (.A(_02585_),
    .B(_02587_),
    .Y(_02588_));
 sky130_fd_sc_hd__o22a_1 _09499_ (.A1(net154),
    .A2(net14),
    .B1(net13),
    .B2(net156),
    .X(_02589_));
 sky130_fd_sc_hd__xnor2_2 _09500_ (.A(net207),
    .B(_02589_),
    .Y(_02590_));
 sky130_fd_sc_hd__nor2_1 _09501_ (.A(net239),
    .B(_02590_),
    .Y(_02591_));
 sky130_fd_sc_hd__xnor2_2 _09502_ (.A(_06493_),
    .B(_02590_),
    .Y(_02592_));
 sky130_fd_sc_hd__a21oi_1 _09503_ (.A1(_06565_),
    .A2(net9),
    .B1(net205),
    .Y(_02593_));
 sky130_fd_sc_hd__a31o_2 _09504_ (.A1(net205),
    .A2(_06555_),
    .A3(net9),
    .B1(_02593_),
    .X(_02594_));
 sky130_fd_sc_hd__xnor2_2 _09505_ (.A(_02592_),
    .B(_02594_),
    .Y(_02595_));
 sky130_fd_sc_hd__nor2_1 _09506_ (.A(_02588_),
    .B(_02595_),
    .Y(_02596_));
 sky130_fd_sc_hd__xor2_1 _09507_ (.A(_02588_),
    .B(_02595_),
    .X(_02597_));
 sky130_fd_sc_hd__xnor2_1 _09508_ (.A(_02578_),
    .B(_02597_),
    .Y(_02598_));
 sky130_fd_sc_hd__nor2_1 _09509_ (.A(_02568_),
    .B(_02598_),
    .Y(_02599_));
 sky130_fd_sc_hd__xor2_1 _09510_ (.A(_02568_),
    .B(_02598_),
    .X(_02600_));
 sky130_fd_sc_hd__xor2_1 _09511_ (.A(_02561_),
    .B(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__nor2_1 _09512_ (.A(_02360_),
    .B(_02365_),
    .Y(_02602_));
 sky130_fd_sc_hd__o22a_1 _09513_ (.A1(net28),
    .A2(net85),
    .B1(net81),
    .B2(net25),
    .X(_02603_));
 sky130_fd_sc_hd__xnor2_1 _09514_ (.A(_00301_),
    .B(_02603_),
    .Y(_02604_));
 sky130_fd_sc_hd__o22a_1 _09515_ (.A1(net48),
    .A2(net119),
    .B1(net117),
    .B2(net46),
    .X(_02605_));
 sky130_fd_sc_hd__xnor2_1 _09516_ (.A(net97),
    .B(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__and2_1 _09517_ (.A(_02604_),
    .B(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__nor2_1 _09518_ (.A(_02604_),
    .B(_02606_),
    .Y(_02608_));
 sky130_fd_sc_hd__nor2_1 _09519_ (.A(_02607_),
    .B(_02608_),
    .Y(_02609_));
 sky130_fd_sc_hd__a22o_1 _09520_ (.A1(net32),
    .A2(_00361_),
    .B1(_00366_),
    .B2(net29),
    .X(_02610_));
 sky130_fd_sc_hd__xnor2_1 _09521_ (.A(net50),
    .B(_02610_),
    .Y(_02611_));
 sky130_fd_sc_hd__xnor2_1 _09522_ (.A(_02609_),
    .B(_02611_),
    .Y(_02612_));
 sky130_fd_sc_hd__o31a_1 _09523_ (.A1(net144),
    .A2(net21),
    .A3(_02421_),
    .B1(_02420_),
    .X(_02613_));
 sky130_fd_sc_hd__nor2_1 _09524_ (.A(_02612_),
    .B(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__xor2_1 _09525_ (.A(_02612_),
    .B(_02613_),
    .X(_02615_));
 sky130_fd_sc_hd__and2b_1 _09526_ (.A_N(_02602_),
    .B(_02615_),
    .X(_02616_));
 sky130_fd_sc_hd__xnor2_1 _09527_ (.A(_02602_),
    .B(_02615_),
    .Y(_02617_));
 sky130_fd_sc_hd__and2_1 _09528_ (.A(_02601_),
    .B(_02617_),
    .X(_02618_));
 sky130_fd_sc_hd__nor2_1 _09529_ (.A(_02601_),
    .B(_02617_),
    .Y(_02619_));
 sky130_fd_sc_hd__nor2_2 _09530_ (.A(_02618_),
    .B(_02619_),
    .Y(_02620_));
 sky130_fd_sc_hd__xor2_4 _09531_ (.A(_02554_),
    .B(_02620_),
    .X(_02621_));
 sky130_fd_sc_hd__a21o_2 _09532_ (.A1(_02427_),
    .A2(_02442_),
    .B1(_02444_),
    .X(_02622_));
 sky130_fd_sc_hd__a21o_1 _09533_ (.A1(_02448_),
    .A2(_02452_),
    .B1(_02451_),
    .X(_02623_));
 sky130_fd_sc_hd__a21o_1 _09534_ (.A1(_02355_),
    .A2(_02370_),
    .B1(_02368_),
    .X(_02624_));
 sky130_fd_sc_hd__a21bo_1 _09535_ (.A1(_02377_),
    .A2(_02425_),
    .B1_N(_02424_),
    .X(_02625_));
 sky130_fd_sc_hd__a21o_1 _09536_ (.A1(_02428_),
    .A2(_02441_),
    .B1(_02440_),
    .X(_02626_));
 sky130_fd_sc_hd__and2_1 _09537_ (.A(_02625_),
    .B(_02626_),
    .X(_02627_));
 sky130_fd_sc_hd__xor2_2 _09538_ (.A(_02625_),
    .B(_02626_),
    .X(_02628_));
 sky130_fd_sc_hd__xor2_2 _09539_ (.A(_02624_),
    .B(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__xnor2_2 _09540_ (.A(_02623_),
    .B(_02629_),
    .Y(_02630_));
 sky130_fd_sc_hd__nand2b_1 _09541_ (.A_N(_02630_),
    .B(_02622_),
    .Y(_02631_));
 sky130_fd_sc_hd__xnor2_4 _09542_ (.A(_02622_),
    .B(_02630_),
    .Y(_02632_));
 sky130_fd_sc_hd__and2_1 _09543_ (.A(_02621_),
    .B(_02632_),
    .X(_02633_));
 sky130_fd_sc_hd__xor2_4 _09544_ (.A(_02621_),
    .B(_02632_),
    .X(_02634_));
 sky130_fd_sc_hd__xnor2_4 _09545_ (.A(_02537_),
    .B(_02634_),
    .Y(_02635_));
 sky130_fd_sc_hd__or2_2 _09546_ (.A(_02536_),
    .B(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__and2_1 _09547_ (.A(_02536_),
    .B(_02635_),
    .X(_02637_));
 sky130_fd_sc_hd__xnor2_4 _09548_ (.A(_02536_),
    .B(_02635_),
    .Y(_02638_));
 sky130_fd_sc_hd__or4_1 _09549_ (.A(_02009_),
    .B(_02126_),
    .C(_02238_),
    .D(_02462_),
    .X(_02639_));
 sky130_fd_sc_hd__o22ai_1 _09550_ (.A1(_02137_),
    .A2(_02236_),
    .B1(_02353_),
    .B2(_02460_),
    .Y(_02640_));
 sky130_fd_sc_hd__a21bo_1 _09551_ (.A1(_02353_),
    .A2(_02460_),
    .B1_N(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__or4_1 _09552_ (.A(_02125_),
    .B(_02134_),
    .C(_02238_),
    .D(_02462_),
    .X(_02642_));
 sky130_fd_sc_hd__o211a_4 _09553_ (.A1(_02014_),
    .A2(_02639_),
    .B1(_02641_),
    .C1(_02642_),
    .X(_02643_));
 sky130_fd_sc_hd__xor2_4 _09554_ (.A(_02638_),
    .B(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__xnor2_1 _09555_ (.A(_02535_),
    .B(_02644_),
    .Y(_02645_));
 sky130_fd_sc_hd__nand2_1 _09556_ (.A(net163),
    .B(_01755_),
    .Y(_02646_));
 sky130_fd_sc_hd__mux2_1 _09557_ (.A0(_01753_),
    .A1(_01806_),
    .S(_02646_),
    .X(_02647_));
 sky130_fd_sc_hd__o21ai_1 _09558_ (.A1(net219),
    .A2(_02489_),
    .B1(_02339_),
    .Y(_02648_));
 sky130_fd_sc_hd__a21oi_2 _09559_ (.A1(net224),
    .A2(_02648_),
    .B1(_02341_),
    .Y(_02649_));
 sky130_fd_sc_hd__inv_2 _09560_ (.A(_02649_),
    .Y(_02650_));
 sky130_fd_sc_hd__o21ai_2 _09561_ (.A1(net227),
    .A2(_02649_),
    .B1(_02335_),
    .Y(_02651_));
 sky130_fd_sc_hd__inv_2 _09562_ (.A(_02651_),
    .Y(_02652_));
 sky130_fd_sc_hd__mux2_1 _09563_ (.A0(_02251_),
    .A1(_02255_),
    .S(net218),
    .X(_02653_));
 sky130_fd_sc_hd__mux2_1 _09564_ (.A0(_02258_),
    .A1(_02263_),
    .S(net217),
    .X(_02654_));
 sky130_fd_sc_hd__mux2_1 _09565_ (.A0(_02653_),
    .A1(_02654_),
    .S(net220),
    .X(_02655_));
 sky130_fd_sc_hd__mux2_1 _09566_ (.A0(_02266_),
    .A1(_02270_),
    .S(net217),
    .X(_02656_));
 sky130_fd_sc_hd__mux2_1 _09567_ (.A0(_02273_),
    .A1(_02294_),
    .S(net217),
    .X(_02657_));
 sky130_fd_sc_hd__mux2_1 _09568_ (.A0(_02656_),
    .A1(_02657_),
    .S(net219),
    .X(_02658_));
 sky130_fd_sc_hd__mux2_1 _09569_ (.A0(_02655_),
    .A1(_02658_),
    .S(net222),
    .X(_02659_));
 sky130_fd_sc_hd__mux2_1 _09570_ (.A0(_02282_),
    .A1(_02286_),
    .S(net218),
    .X(_02660_));
 sky130_fd_sc_hd__mux2_1 _09571_ (.A0(_02525_),
    .A1(_02660_),
    .S(_06352_),
    .X(_02661_));
 sky130_fd_sc_hd__mux2_1 _09572_ (.A0(_02297_),
    .A1(_02301_),
    .S(net217),
    .X(_02662_));
 sky130_fd_sc_hd__mux2_1 _09573_ (.A0(_02279_),
    .A1(_02304_),
    .S(_06359_),
    .X(_02663_));
 sky130_fd_sc_hd__mux2_1 _09574_ (.A0(_02662_),
    .A1(_02663_),
    .S(net219),
    .X(_02664_));
 sky130_fd_sc_hd__mux2_1 _09575_ (.A0(_02661_),
    .A1(_02664_),
    .S(net224),
    .X(_02665_));
 sky130_fd_sc_hd__mux2_2 _09576_ (.A0(_02659_),
    .A1(_02665_),
    .S(net226),
    .X(_02666_));
 sky130_fd_sc_hd__o21a_1 _09577_ (.A1(_02309_),
    .A2(_02503_),
    .B1(_02502_),
    .X(_02667_));
 sky130_fd_sc_hd__nor2_1 _09578_ (.A(reg1_val[2]),
    .B(curr_PC[2]),
    .Y(_02668_));
 sky130_fd_sc_hd__nand2_1 _09579_ (.A(reg1_val[2]),
    .B(curr_PC[2]),
    .Y(_02669_));
 sky130_fd_sc_hd__nand2b_1 _09580_ (.A_N(_02668_),
    .B(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__xnor2_1 _09581_ (.A(_02667_),
    .B(_02670_),
    .Y(_02671_));
 sky130_fd_sc_hd__or2_1 _09582_ (.A(\div_res[1] ),
    .B(\div_res[0] ),
    .X(_02672_));
 sky130_fd_sc_hd__a21oi_1 _09583_ (.A1(net167),
    .A2(_02672_),
    .B1(\div_res[2] ),
    .Y(_02673_));
 sky130_fd_sc_hd__a31o_1 _09584_ (.A1(\div_res[2] ),
    .A2(net167),
    .A3(_02672_),
    .B1(net195),
    .X(_02674_));
 sky130_fd_sc_hd__a22o_1 _09585_ (.A1(reg1_val[1]),
    .A2(_06360_),
    .B1(net214),
    .B2(net292),
    .X(_02675_));
 sky130_fd_sc_hd__nand2_1 _09586_ (.A(_06361_),
    .B(_02675_),
    .Y(_02676_));
 sky130_fd_sc_hd__mux2_1 _09587_ (.A0(_06368_),
    .A1(_02676_),
    .S(net285),
    .X(_02677_));
 sky130_fd_sc_hd__a21oi_1 _09588_ (.A1(_06357_),
    .A2(_02677_),
    .B1(net236),
    .Y(_02678_));
 sky130_fd_sc_hd__o21ai_1 _09589_ (.A1(_06357_),
    .A2(_02677_),
    .B1(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__or2_1 _09590_ (.A(\div_shifter[33] ),
    .B(\div_shifter[32] ),
    .X(_02680_));
 sky130_fd_sc_hd__a21oi_1 _09591_ (.A1(net235),
    .A2(_02680_),
    .B1(\div_shifter[34] ),
    .Y(_02681_));
 sky130_fd_sc_hd__a31o_1 _09592_ (.A1(\div_shifter[34] ),
    .A2(net235),
    .A3(_02680_),
    .B1(net193),
    .X(_02682_));
 sky130_fd_sc_hd__or2_1 _09593_ (.A(_02681_),
    .B(_02682_),
    .X(_02683_));
 sky130_fd_sc_hd__or2_1 _09594_ (.A(net294),
    .B(_02666_),
    .X(_02684_));
 sky130_fd_sc_hd__o211a_1 _09595_ (.A1(net284),
    .A2(_02652_),
    .B1(_02684_),
    .C1(_06479_),
    .X(_02685_));
 sky130_fd_sc_hd__nor2_1 _09596_ (.A(net249),
    .B(_02666_),
    .Y(_02686_));
 sky130_fd_sc_hd__a211o_1 _09597_ (.A1(net249),
    .A2(_02671_),
    .B1(_02686_),
    .C1(_06476_),
    .X(_02687_));
 sky130_fd_sc_hd__o221a_1 _09598_ (.A1(_06355_),
    .A2(net199),
    .B1(net196),
    .B2(_06354_),
    .C1(_02683_),
    .X(_02688_));
 sky130_fd_sc_hd__o211a_1 _09599_ (.A1(_06357_),
    .A2(net197),
    .B1(_02679_),
    .C1(_02688_),
    .X(_02689_));
 sky130_fd_sc_hd__o211a_1 _09600_ (.A1(_02673_),
    .A2(_02674_),
    .B1(_02687_),
    .C1(_02689_),
    .X(_02690_));
 sky130_fd_sc_hd__a22o_1 _09601_ (.A1(net221),
    .A2(net241),
    .B1(net200),
    .B2(_02645_),
    .X(_02691_));
 sky130_fd_sc_hd__or3b_1 _09602_ (.A(_02691_),
    .B(_02685_),
    .C_N(_02690_),
    .X(_02692_));
 sky130_fd_sc_hd__a21oi_2 _09603_ (.A1(_02323_),
    .A2(_02647_),
    .B1(_02692_),
    .Y(_02693_));
 sky130_fd_sc_hd__o21ai_4 _09604_ (.A1(net248),
    .A2(_02693_),
    .B1(_02534_),
    .Y(dest_val[2]));
 sky130_fd_sc_hd__o31ai_1 _09605_ (.A1(_02352_),
    .A2(_02467_),
    .A3(_02644_),
    .B1(net163),
    .Y(_02694_));
 sky130_fd_sc_hd__a21oi_4 _09606_ (.A1(_02537_),
    .A2(_02634_),
    .B1(_02633_),
    .Y(_02695_));
 sky130_fd_sc_hd__a21bo_2 _09607_ (.A1(_02623_),
    .A2(_02629_),
    .B1_N(_02631_),
    .X(_02696_));
 sky130_fd_sc_hd__a21o_2 _09608_ (.A1(_02578_),
    .A2(_02597_),
    .B1(_02596_),
    .X(_02697_));
 sky130_fd_sc_hd__o22a_1 _09609_ (.A1(net114),
    .A2(net24),
    .B1(net16),
    .B2(_00375_),
    .X(_02698_));
 sky130_fd_sc_hd__xnor2_2 _09610_ (.A(net71),
    .B(_02698_),
    .Y(_02699_));
 sky130_fd_sc_hd__inv_2 _09611_ (.A(_02699_),
    .Y(_02700_));
 sky130_fd_sc_hd__a22o_1 _09612_ (.A1(net39),
    .A2(net116),
    .B1(_00324_),
    .B2(net37),
    .X(_02701_));
 sky130_fd_sc_hd__xor2_1 _09613_ (.A(net91),
    .B(_02701_),
    .X(_02702_));
 sky130_fd_sc_hd__xor2_1 _09614_ (.A(_02699_),
    .B(_02702_),
    .X(_02703_));
 sky130_fd_sc_hd__a22o_1 _09615_ (.A1(net42),
    .A2(_00308_),
    .B1(_00330_),
    .B2(net44),
    .X(_02704_));
 sky130_fd_sc_hd__xor2_1 _09616_ (.A(net94),
    .B(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__and2b_1 _09617_ (.A_N(_02703_),
    .B(_02705_),
    .X(_02706_));
 sky130_fd_sc_hd__and2b_1 _09618_ (.A_N(_02705_),
    .B(_02703_),
    .X(_02707_));
 sky130_fd_sc_hd__or2_1 _09619_ (.A(_02706_),
    .B(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__a21oi_1 _09620_ (.A1(_02558_),
    .A2(_02560_),
    .B1(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__and3_1 _09621_ (.A(_02558_),
    .B(_02560_),
    .C(_02708_),
    .X(_02710_));
 sky130_fd_sc_hd__nor2_2 _09622_ (.A(_02709_),
    .B(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__xor2_4 _09623_ (.A(_02697_),
    .B(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__or2_1 _09624_ (.A(_02542_),
    .B(_02547_),
    .X(_02713_));
 sky130_fd_sc_hd__o22a_1 _09625_ (.A1(net99),
    .A2(net28),
    .B1(net26),
    .B2(net85),
    .X(_02714_));
 sky130_fd_sc_hd__xnor2_2 _09626_ (.A(net89),
    .B(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__o22a_1 _09627_ (.A1(net46),
    .A2(net120),
    .B1(net73),
    .B2(net48),
    .X(_02716_));
 sky130_fd_sc_hd__xnor2_2 _09628_ (.A(net97),
    .B(_02716_),
    .Y(_02717_));
 sky130_fd_sc_hd__and2_1 _09629_ (.A(_02715_),
    .B(_02717_),
    .X(_02718_));
 sky130_fd_sc_hd__xor2_2 _09630_ (.A(_02715_),
    .B(_02717_),
    .X(_02719_));
 sky130_fd_sc_hd__a22o_1 _09631_ (.A1(net31),
    .A2(_00354_),
    .B1(_00361_),
    .B2(net29),
    .X(_02720_));
 sky130_fd_sc_hd__xnor2_2 _09632_ (.A(net49),
    .B(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__xnor2_1 _09633_ (.A(_02719_),
    .B(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__a21o_1 _09634_ (.A1(_02562_),
    .A2(_02566_),
    .B1(_02565_),
    .X(_02723_));
 sky130_fd_sc_hd__nand2b_1 _09635_ (.A_N(_02722_),
    .B(_02723_),
    .Y(_02724_));
 sky130_fd_sc_hd__xnor2_1 _09636_ (.A(_02722_),
    .B(_02723_),
    .Y(_02725_));
 sky130_fd_sc_hd__nand2_1 _09637_ (.A(_02713_),
    .B(_02725_),
    .Y(_02726_));
 sky130_fd_sc_hd__or2_1 _09638_ (.A(_02713_),
    .B(_02725_),
    .X(_02727_));
 sky130_fd_sc_hd__nand2_1 _09639_ (.A(_02726_),
    .B(_02727_),
    .Y(_02728_));
 sky130_fd_sc_hd__o21a_1 _09640_ (.A1(_02585_),
    .A2(_02587_),
    .B1(_02583_),
    .X(_02729_));
 sky130_fd_sc_hd__o21bai_2 _09641_ (.A1(_02574_),
    .A2(_02577_),
    .B1_N(_02573_),
    .Y(_02730_));
 sky130_fd_sc_hd__a21o_1 _09642_ (.A1(_02609_),
    .A2(_02611_),
    .B1(_02607_),
    .X(_02731_));
 sky130_fd_sc_hd__nand2_1 _09643_ (.A(_02730_),
    .B(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__xor2_1 _09644_ (.A(_02730_),
    .B(_02731_),
    .X(_02733_));
 sky130_fd_sc_hd__nand2b_1 _09645_ (.A_N(_02729_),
    .B(_02733_),
    .Y(_02734_));
 sky130_fd_sc_hd__xnor2_1 _09646_ (.A(_02729_),
    .B(_02733_),
    .Y(_02735_));
 sky130_fd_sc_hd__o22a_1 _09647_ (.A1(net65),
    .A2(net106),
    .B1(net104),
    .B2(net59),
    .X(_02736_));
 sky130_fd_sc_hd__xnor2_1 _09648_ (.A(_00342_),
    .B(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__a21o_1 _09649_ (.A1(_00697_),
    .A2(_00698_),
    .B1(net148),
    .X(_02738_));
 sky130_fd_sc_hd__or3_1 _09650_ (.A(net146),
    .B(_00405_),
    .C(_00407_),
    .X(_02739_));
 sky130_fd_sc_hd__a21o_1 _09651_ (.A1(_02738_),
    .A2(_02739_),
    .B1(net202),
    .X(_02740_));
 sky130_fd_sc_hd__nand3_1 _09652_ (.A(net202),
    .B(_02738_),
    .C(_02739_),
    .Y(_02741_));
 sky130_fd_sc_hd__and3_1 _09653_ (.A(_02737_),
    .B(_02740_),
    .C(_02741_),
    .X(_02742_));
 sky130_fd_sc_hd__a21oi_1 _09654_ (.A1(_02740_),
    .A2(_02741_),
    .B1(_02737_),
    .Y(_02743_));
 sky130_fd_sc_hd__nor2_1 _09655_ (.A(_02742_),
    .B(_02743_),
    .Y(_02744_));
 sky130_fd_sc_hd__o22a_1 _09656_ (.A1(net56),
    .A2(net134),
    .B1(net132),
    .B2(net68),
    .X(_02745_));
 sky130_fd_sc_hd__xnor2_2 _09657_ (.A(net182),
    .B(_02745_),
    .Y(_02746_));
 sky130_fd_sc_hd__xnor2_2 _09658_ (.A(_02744_),
    .B(_02746_),
    .Y(_02747_));
 sky130_fd_sc_hd__o22a_1 _09659_ (.A1(net57),
    .A2(net86),
    .B1(net82),
    .B2(net63),
    .X(_02748_));
 sky130_fd_sc_hd__xnor2_1 _09660_ (.A(_00338_),
    .B(_02748_),
    .Y(_02749_));
 sky130_fd_sc_hd__o22a_1 _09661_ (.A1(net51),
    .A2(net35),
    .B1(net33),
    .B2(net100),
    .X(_02750_));
 sky130_fd_sc_hd__xnor2_1 _09662_ (.A(net124),
    .B(_02750_),
    .Y(_02751_));
 sky130_fd_sc_hd__or2_1 _09663_ (.A(_02749_),
    .B(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__nand2_1 _09664_ (.A(_02749_),
    .B(_02751_),
    .Y(_02753_));
 sky130_fd_sc_hd__nand2_1 _09665_ (.A(_02752_),
    .B(_02753_),
    .Y(_02754_));
 sky130_fd_sc_hd__o22a_1 _09666_ (.A1(net61),
    .A2(_00360_),
    .B1(net75),
    .B2(net53),
    .X(_02755_));
 sky130_fd_sc_hd__xnor2_2 _09667_ (.A(net121),
    .B(_02755_),
    .Y(_02756_));
 sky130_fd_sc_hd__xnor2_2 _09668_ (.A(_02754_),
    .B(_02756_),
    .Y(_02757_));
 sky130_fd_sc_hd__o22a_1 _09669_ (.A1(net154),
    .A2(net13),
    .B1(net8),
    .B2(net156),
    .X(_02758_));
 sky130_fd_sc_hd__xnor2_2 _09670_ (.A(net208),
    .B(_02758_),
    .Y(_02759_));
 sky130_fd_sc_hd__nor2_1 _09671_ (.A(_06493_),
    .B(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__xnor2_2 _09672_ (.A(net239),
    .B(_02759_),
    .Y(_02761_));
 sky130_fd_sc_hd__xnor2_2 _09673_ (.A(net205),
    .B(_02761_),
    .Y(_02762_));
 sky130_fd_sc_hd__nor2_1 _09674_ (.A(_02757_),
    .B(_02762_),
    .Y(_02763_));
 sky130_fd_sc_hd__xor2_2 _09675_ (.A(_02757_),
    .B(_02762_),
    .X(_02764_));
 sky130_fd_sc_hd__xnor2_2 _09676_ (.A(_02747_),
    .B(_02764_),
    .Y(_02765_));
 sky130_fd_sc_hd__nor2_1 _09677_ (.A(net142),
    .B(net21),
    .Y(_02766_));
 sky130_fd_sc_hd__a21oi_2 _09678_ (.A1(_02592_),
    .A2(_02594_),
    .B1(_02591_),
    .Y(_02767_));
 sky130_fd_sc_hd__o22a_1 _09679_ (.A1(net130),
    .A2(net11),
    .B1(net6),
    .B2(net128),
    .X(_02768_));
 sky130_fd_sc_hd__xnor2_2 _09680_ (.A(net22),
    .B(_02768_),
    .Y(_02769_));
 sky130_fd_sc_hd__nand2b_1 _09681_ (.A_N(_02767_),
    .B(_02769_),
    .Y(_02770_));
 sky130_fd_sc_hd__xnor2_2 _09682_ (.A(_02767_),
    .B(_02769_),
    .Y(_02771_));
 sky130_fd_sc_hd__xnor2_2 _09683_ (.A(_02766_),
    .B(_02771_),
    .Y(_02772_));
 sky130_fd_sc_hd__nor2_1 _09684_ (.A(_02765_),
    .B(_02772_),
    .Y(_02773_));
 sky130_fd_sc_hd__xor2_2 _09685_ (.A(_02765_),
    .B(_02772_),
    .X(_02774_));
 sky130_fd_sc_hd__xnor2_1 _09686_ (.A(_02735_),
    .B(_02774_),
    .Y(_02775_));
 sky130_fd_sc_hd__nor2_1 _09687_ (.A(_02728_),
    .B(_02775_),
    .Y(_02776_));
 sky130_fd_sc_hd__nand2_1 _09688_ (.A(_02728_),
    .B(_02775_),
    .Y(_02777_));
 sky130_fd_sc_hd__and2b_1 _09689_ (.A_N(_02776_),
    .B(_02777_),
    .X(_02778_));
 sky130_fd_sc_hd__xor2_4 _09690_ (.A(_02712_),
    .B(_02778_),
    .X(_02779_));
 sky130_fd_sc_hd__a21o_1 _09691_ (.A1(_02554_),
    .A2(_02620_),
    .B1(_02618_),
    .X(_02780_));
 sky130_fd_sc_hd__o21ai_4 _09692_ (.A1(_02549_),
    .A2(_02550_),
    .B1(_02552_),
    .Y(_02781_));
 sky130_fd_sc_hd__a21o_2 _09693_ (.A1(_02561_),
    .A2(_02600_),
    .B1(_02599_),
    .X(_02782_));
 sky130_fd_sc_hd__nor2_2 _09694_ (.A(_02614_),
    .B(_02616_),
    .Y(_02783_));
 sky130_fd_sc_hd__o21ai_1 _09695_ (.A1(_02614_),
    .A2(_02616_),
    .B1(_02782_),
    .Y(_02784_));
 sky130_fd_sc_hd__xnor2_4 _09696_ (.A(_02782_),
    .B(_02783_),
    .Y(_02785_));
 sky130_fd_sc_hd__xnor2_4 _09697_ (.A(_02781_),
    .B(_02785_),
    .Y(_02786_));
 sky130_fd_sc_hd__a21oi_2 _09698_ (.A1(_02624_),
    .A2(_02628_),
    .B1(_02627_),
    .Y(_02787_));
 sky130_fd_sc_hd__xnor2_2 _09699_ (.A(_02786_),
    .B(_02787_),
    .Y(_02788_));
 sky130_fd_sc_hd__nand2b_1 _09700_ (.A_N(_02788_),
    .B(_02780_),
    .Y(_02789_));
 sky130_fd_sc_hd__xnor2_2 _09701_ (.A(_02780_),
    .B(_02788_),
    .Y(_02790_));
 sky130_fd_sc_hd__and2_1 _09702_ (.A(_02779_),
    .B(_02790_),
    .X(_02791_));
 sky130_fd_sc_hd__xor2_4 _09703_ (.A(_02779_),
    .B(_02790_),
    .X(_02792_));
 sky130_fd_sc_hd__xnor2_4 _09704_ (.A(_02696_),
    .B(_02792_),
    .Y(_02793_));
 sky130_fd_sc_hd__or2_1 _09705_ (.A(_02695_),
    .B(_02793_),
    .X(_02794_));
 sky130_fd_sc_hd__and2_1 _09706_ (.A(_02695_),
    .B(_02793_),
    .X(_02795_));
 sky130_fd_sc_hd__xnor2_4 _09707_ (.A(_02695_),
    .B(_02793_),
    .Y(_02796_));
 sky130_fd_sc_hd__or4_1 _09708_ (.A(_02126_),
    .B(_02238_),
    .C(_02462_),
    .D(_02638_),
    .X(_02797_));
 sky130_fd_sc_hd__a21oi_1 _09709_ (.A1(_02461_),
    .A2(_02636_),
    .B1(_02637_),
    .Y(_02798_));
 sky130_fd_sc_hd__a21o_1 _09710_ (.A1(_02461_),
    .A2(_02636_),
    .B1(_02637_),
    .X(_02799_));
 sky130_fd_sc_hd__or4_1 _09711_ (.A(_02237_),
    .B(_02462_),
    .C(_02464_),
    .D(_02638_),
    .X(_02800_));
 sky130_fd_sc_hd__o211a_2 _09712_ (.A1(_02130_),
    .A2(_02797_),
    .B1(_02799_),
    .C1(_02800_),
    .X(_02801_));
 sky130_fd_sc_hd__xnor2_2 _09713_ (.A(_02796_),
    .B(_02801_),
    .Y(_02802_));
 sky130_fd_sc_hd__or2_1 _09714_ (.A(_02694_),
    .B(_02802_),
    .X(_02803_));
 sky130_fd_sc_hd__nand2_1 _09715_ (.A(_02694_),
    .B(_02802_),
    .Y(_02804_));
 sky130_fd_sc_hd__o21ai_1 _09716_ (.A1(net159),
    .A2(_01807_),
    .B1(_01809_),
    .Y(_02805_));
 sky130_fd_sc_hd__or3_1 _09717_ (.A(net159),
    .B(_01807_),
    .C(_01809_),
    .X(_02806_));
 sky130_fd_sc_hd__mux2_1 _09718_ (.A0(_02471_),
    .A1(_02473_),
    .S(net218),
    .X(_02807_));
 sky130_fd_sc_hd__mux2_1 _09719_ (.A0(_02474_),
    .A1(_02477_),
    .S(net217),
    .X(_02808_));
 sky130_fd_sc_hd__mux2_1 _09720_ (.A0(_02807_),
    .A1(_02808_),
    .S(net220),
    .X(_02809_));
 sky130_fd_sc_hd__mux2_1 _09721_ (.A0(_02478_),
    .A1(_02480_),
    .S(net217),
    .X(_02810_));
 sky130_fd_sc_hd__mux2_1 _09722_ (.A0(_02481_),
    .A1(_02491_),
    .S(net217),
    .X(_02811_));
 sky130_fd_sc_hd__mux2_1 _09723_ (.A0(_02810_),
    .A1(_02811_),
    .S(net219),
    .X(_02812_));
 sky130_fd_sc_hd__mux2_1 _09724_ (.A0(_02809_),
    .A1(_02812_),
    .S(net222),
    .X(_02813_));
 sky130_fd_sc_hd__mux2_1 _09725_ (.A0(_02486_),
    .A1(_02488_),
    .S(net218),
    .X(_02814_));
 sky130_fd_sc_hd__mux2_1 _09726_ (.A0(_02338_),
    .A1(_02814_),
    .S(_06352_),
    .X(_02815_));
 sky130_fd_sc_hd__mux2_1 _09727_ (.A0(_02492_),
    .A1(_02494_),
    .S(net217),
    .X(_02816_));
 sky130_fd_sc_hd__mux2_1 _09728_ (.A0(_02485_),
    .A1(_02495_),
    .S(_06359_),
    .X(_02817_));
 sky130_fd_sc_hd__mux2_1 _09729_ (.A0(_02816_),
    .A1(_02817_),
    .S(net219),
    .X(_02818_));
 sky130_fd_sc_hd__mux2_1 _09730_ (.A0(_02815_),
    .A1(_02818_),
    .S(net224),
    .X(_02819_));
 sky130_fd_sc_hd__mux2_2 _09731_ (.A0(_02813_),
    .A1(_02819_),
    .S(net226),
    .X(_02820_));
 sky130_fd_sc_hd__or2_1 _09732_ (.A(net250),
    .B(_02820_),
    .X(_02821_));
 sky130_fd_sc_hd__o21a_1 _09733_ (.A1(_02667_),
    .A2(_02668_),
    .B1(_02669_),
    .X(_02822_));
 sky130_fd_sc_hd__nor2_1 _09734_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .Y(_02823_));
 sky130_fd_sc_hd__nand2_1 _09735_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .Y(_02824_));
 sky130_fd_sc_hd__and2b_1 _09736_ (.A_N(_02823_),
    .B(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__o21ai_1 _09737_ (.A1(_02822_),
    .A2(_02825_),
    .B1(net249),
    .Y(_02826_));
 sky130_fd_sc_hd__a21o_1 _09738_ (.A1(_02822_),
    .A2(_02825_),
    .B1(_02826_),
    .X(_02827_));
 sky130_fd_sc_hd__o21a_1 _09739_ (.A1(net219),
    .A2(_02290_),
    .B1(_02339_),
    .X(_02828_));
 sky130_fd_sc_hd__o21a_1 _09740_ (.A1(net222),
    .A2(_02828_),
    .B1(_02342_),
    .X(_02829_));
 sky130_fd_sc_hd__o21a_2 _09741_ (.A1(net227),
    .A2(_02829_),
    .B1(_02335_),
    .X(_02830_));
 sky130_fd_sc_hd__a21boi_1 _09742_ (.A1(_06361_),
    .A2(_02675_),
    .B1_N(_06354_),
    .Y(_02831_));
 sky130_fd_sc_hd__or3_1 _09743_ (.A(net294),
    .B(_06355_),
    .C(_02831_),
    .X(_02832_));
 sky130_fd_sc_hd__o21ai_1 _09744_ (.A1(net285),
    .A2(_06370_),
    .B1(_02832_),
    .Y(_02833_));
 sky130_fd_sc_hd__nand2b_1 _09745_ (.A_N(_02833_),
    .B(_06350_),
    .Y(_02834_));
 sky130_fd_sc_hd__nand2b_1 _09746_ (.A_N(_06350_),
    .B(_02833_),
    .Y(_02835_));
 sky130_fd_sc_hd__or3_1 _09747_ (.A(\div_res[2] ),
    .B(\div_res[1] ),
    .C(\div_res[0] ),
    .X(_02836_));
 sky130_fd_sc_hd__a21oi_1 _09748_ (.A1(net167),
    .A2(_02836_),
    .B1(\div_res[3] ),
    .Y(_02837_));
 sky130_fd_sc_hd__a31o_1 _09749_ (.A1(\div_res[3] ),
    .A2(net167),
    .A3(_02836_),
    .B1(net195),
    .X(_02838_));
 sky130_fd_sc_hd__o31a_1 _09750_ (.A1(\div_shifter[34] ),
    .A2(\div_shifter[33] ),
    .A3(\div_shifter[32] ),
    .B1(net235),
    .X(_02839_));
 sky130_fd_sc_hd__o21ai_1 _09751_ (.A1(\div_shifter[35] ),
    .A2(_02839_),
    .B1(_02330_),
    .Y(_02840_));
 sky130_fd_sc_hd__a21o_1 _09752_ (.A1(\div_shifter[35] ),
    .A2(_02839_),
    .B1(_02840_),
    .X(_02841_));
 sky130_fd_sc_hd__o221a_1 _09753_ (.A1(net224),
    .A2(net209),
    .B1(net196),
    .B2(_06349_),
    .C1(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__o221a_1 _09754_ (.A1(_06348_),
    .A2(net199),
    .B1(net197),
    .B2(_06350_),
    .C1(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__o21ai_1 _09755_ (.A1(_02837_),
    .A2(_02838_),
    .B1(_02843_),
    .Y(_02844_));
 sky130_fd_sc_hd__a31o_1 _09756_ (.A1(_02317_),
    .A2(_02834_),
    .A3(_02835_),
    .B1(_02844_),
    .X(_02845_));
 sky130_fd_sc_hd__a221o_1 _09757_ (.A1(_02313_),
    .A2(_02820_),
    .B1(_02830_),
    .B2(net179),
    .C1(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__a31o_1 _09758_ (.A1(net210),
    .A2(_02821_),
    .A3(_02827_),
    .B1(_02846_),
    .X(_02847_));
 sky130_fd_sc_hd__a31o_1 _09759_ (.A1(_02323_),
    .A2(_02805_),
    .A3(_02806_),
    .B1(_02847_),
    .X(_02848_));
 sky130_fd_sc_hd__a31o_1 _09760_ (.A1(net200),
    .A2(_02803_),
    .A3(_02804_),
    .B1(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__or2_1 _09761_ (.A(curr_PC[3]),
    .B(_02532_),
    .X(_02850_));
 sky130_fd_sc_hd__and2_1 _09762_ (.A(curr_PC[3]),
    .B(_02532_),
    .X(_02851_));
 sky130_fd_sc_hd__nor2_1 _09763_ (.A(net242),
    .B(_02851_),
    .Y(_02852_));
 sky130_fd_sc_hd__a22o_4 _09764_ (.A1(net242),
    .A2(_02849_),
    .B1(_02850_),
    .B2(_02852_),
    .X(dest_val[3]));
 sky130_fd_sc_hd__nor4b_1 _09765_ (.A(_02352_),
    .B(_02467_),
    .C(_02644_),
    .D_N(_02802_),
    .Y(_02853_));
 sky130_fd_sc_hd__or2_1 _09766_ (.A(net159),
    .B(_02853_),
    .X(_02854_));
 sky130_fd_sc_hd__a21oi_4 _09767_ (.A1(_02696_),
    .A2(_02792_),
    .B1(_02791_),
    .Y(_02855_));
 sky130_fd_sc_hd__o21ai_4 _09768_ (.A1(_02786_),
    .A2(_02787_),
    .B1(_02789_),
    .Y(_02856_));
 sky130_fd_sc_hd__a21o_2 _09769_ (.A1(_02747_),
    .A2(_02764_),
    .B1(_02763_),
    .X(_02857_));
 sky130_fd_sc_hd__o22a_1 _09770_ (.A1(_00309_),
    .A2(net24),
    .B1(net16),
    .B2(net114),
    .X(_02858_));
 sky130_fd_sc_hd__xnor2_1 _09771_ (.A(net71),
    .B(_02858_),
    .Y(_02859_));
 sky130_fd_sc_hd__a22o_1 _09772_ (.A1(net39),
    .A2(net118),
    .B1(net116),
    .B2(net37),
    .X(_02860_));
 sky130_fd_sc_hd__xor2_1 _09773_ (.A(net91),
    .B(_02860_),
    .X(_02861_));
 sky130_fd_sc_hd__and2b_1 _09774_ (.A_N(_02859_),
    .B(_02861_),
    .X(_02862_));
 sky130_fd_sc_hd__and2b_1 _09775_ (.A_N(_02861_),
    .B(_02859_),
    .X(_02863_));
 sky130_fd_sc_hd__or2_1 _09776_ (.A(_02862_),
    .B(_02863_),
    .X(_02864_));
 sky130_fd_sc_hd__inv_2 _09777_ (.A(_02864_),
    .Y(_02865_));
 sky130_fd_sc_hd__a22o_1 _09778_ (.A1(net44),
    .A2(_00324_),
    .B1(_00330_),
    .B2(net42),
    .X(_02866_));
 sky130_fd_sc_hd__xor2_1 _09779_ (.A(net94),
    .B(_02866_),
    .X(_02867_));
 sky130_fd_sc_hd__xor2_1 _09780_ (.A(_02864_),
    .B(_02867_),
    .X(_02868_));
 sky130_fd_sc_hd__a21oi_1 _09781_ (.A1(_02732_),
    .A2(_02734_),
    .B1(_02868_),
    .Y(_02869_));
 sky130_fd_sc_hd__and3_1 _09782_ (.A(_02732_),
    .B(_02734_),
    .C(_02868_),
    .X(_02870_));
 sky130_fd_sc_hd__nor2_2 _09783_ (.A(_02869_),
    .B(_02870_),
    .Y(_02871_));
 sky130_fd_sc_hd__xor2_4 _09784_ (.A(_02857_),
    .B(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__o21a_1 _09785_ (.A1(_02754_),
    .A2(_02756_),
    .B1(_02752_),
    .X(_02873_));
 sky130_fd_sc_hd__a21oi_2 _09786_ (.A1(_02719_),
    .A2(_02721_),
    .B1(_02718_),
    .Y(_02874_));
 sky130_fd_sc_hd__o21ba_1 _09787_ (.A1(_02743_),
    .A2(_02746_),
    .B1_N(_02742_),
    .X(_02875_));
 sky130_fd_sc_hd__xor2_2 _09788_ (.A(_02874_),
    .B(_02875_),
    .X(_02876_));
 sky130_fd_sc_hd__and2b_1 _09789_ (.A_N(_02873_),
    .B(_02876_),
    .X(_02877_));
 sky130_fd_sc_hd__xnor2_2 _09790_ (.A(_02873_),
    .B(_02876_),
    .Y(_02878_));
 sky130_fd_sc_hd__o22a_1 _09791_ (.A1(net68),
    .A2(net106),
    .B1(net104),
    .B2(net65),
    .X(_02879_));
 sky130_fd_sc_hd__xnor2_1 _09792_ (.A(net135),
    .B(_02879_),
    .Y(_02880_));
 sky130_fd_sc_hd__o22a_1 _09793_ (.A1(net59),
    .A2(net86),
    .B1(net82),
    .B2(net57),
    .X(_02881_));
 sky130_fd_sc_hd__xnor2_1 _09794_ (.A(_00338_),
    .B(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__o32a_1 _09795_ (.A1(net134),
    .A2(_00405_),
    .A3(_00407_),
    .B1(net132),
    .B2(net56),
    .X(_02883_));
 sky130_fd_sc_hd__xnor2_1 _09796_ (.A(net182),
    .B(_02883_),
    .Y(_02884_));
 sky130_fd_sc_hd__xnor2_1 _09797_ (.A(_02882_),
    .B(_02884_),
    .Y(_02885_));
 sky130_fd_sc_hd__or2_1 _09798_ (.A(_02880_),
    .B(_02885_),
    .X(_02886_));
 sky130_fd_sc_hd__nand2_1 _09799_ (.A(_02880_),
    .B(_02885_),
    .Y(_02887_));
 sky130_fd_sc_hd__and2_1 _09800_ (.A(_02886_),
    .B(_02887_),
    .X(_02888_));
 sky130_fd_sc_hd__o22a_1 _09801_ (.A1(net101),
    .A2(net28),
    .B1(net26),
    .B2(net99),
    .X(_02889_));
 sky130_fd_sc_hd__xnor2_1 _09802_ (.A(net89),
    .B(_02889_),
    .Y(_02890_));
 sky130_fd_sc_hd__inv_2 _09803_ (.A(_02890_),
    .Y(_02891_));
 sky130_fd_sc_hd__o22a_1 _09804_ (.A1(net63),
    .A2(net78),
    .B1(net74),
    .B2(net62),
    .X(_02892_));
 sky130_fd_sc_hd__xnor2_1 _09805_ (.A(net122),
    .B(_02892_),
    .Y(_02893_));
 sky130_fd_sc_hd__nor2_1 _09806_ (.A(_02891_),
    .B(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__xnor2_1 _09807_ (.A(_02890_),
    .B(_02893_),
    .Y(_02895_));
 sky130_fd_sc_hd__o22a_1 _09808_ (.A1(net53),
    .A2(net35),
    .B1(net34),
    .B2(net51),
    .X(_02896_));
 sky130_fd_sc_hd__xnor2_1 _09809_ (.A(net126),
    .B(_02896_),
    .Y(_02897_));
 sky130_fd_sc_hd__and2_1 _09810_ (.A(_02895_),
    .B(_02897_),
    .X(_02898_));
 sky130_fd_sc_hd__xor2_1 _09811_ (.A(_02895_),
    .B(_02897_),
    .X(_02899_));
 sky130_fd_sc_hd__o22a_1 _09812_ (.A1(net146),
    .A2(net14),
    .B1(net13),
    .B2(net148),
    .X(_02900_));
 sky130_fd_sc_hd__xnor2_1 _09813_ (.A(net202),
    .B(_02900_),
    .Y(_02901_));
 sky130_fd_sc_hd__o21ai_2 _09814_ (.A1(_06537_),
    .A2(net8),
    .B1(_06532_),
    .Y(_02902_));
 sky130_fd_sc_hd__o31ai_4 _09815_ (.A1(_06532_),
    .A2(_06536_),
    .A3(net8),
    .B1(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__and2b_1 _09816_ (.A_N(_02903_),
    .B(_02901_),
    .X(_02904_));
 sky130_fd_sc_hd__xor2_1 _09817_ (.A(_02901_),
    .B(_02903_),
    .X(_02905_));
 sky130_fd_sc_hd__and2_1 _09818_ (.A(_02899_),
    .B(_02905_),
    .X(_02906_));
 sky130_fd_sc_hd__nor2_1 _09819_ (.A(_02899_),
    .B(_02905_),
    .Y(_02907_));
 sky130_fd_sc_hd__nor2_1 _09820_ (.A(_02906_),
    .B(_02907_),
    .Y(_02908_));
 sky130_fd_sc_hd__xnor2_2 _09821_ (.A(_02888_),
    .B(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__nor2_1 _09822_ (.A(net128),
    .B(net21),
    .Y(_02910_));
 sky130_fd_sc_hd__a21oi_2 _09823_ (.A1(net205),
    .A2(_02761_),
    .B1(_02760_),
    .Y(_02911_));
 sky130_fd_sc_hd__o22a_1 _09824_ (.A1(_00375_),
    .A2(net11),
    .B1(net6),
    .B2(net130),
    .X(_02912_));
 sky130_fd_sc_hd__xnor2_2 _09825_ (.A(net21),
    .B(_02912_),
    .Y(_02913_));
 sky130_fd_sc_hd__nor2_1 _09826_ (.A(_02911_),
    .B(_02913_),
    .Y(_02914_));
 sky130_fd_sc_hd__xor2_2 _09827_ (.A(_02911_),
    .B(_02913_),
    .X(_02915_));
 sky130_fd_sc_hd__xnor2_2 _09828_ (.A(_02910_),
    .B(_02915_),
    .Y(_02916_));
 sky130_fd_sc_hd__nor2_1 _09829_ (.A(_02909_),
    .B(_02916_),
    .Y(_02917_));
 sky130_fd_sc_hd__xor2_2 _09830_ (.A(_02909_),
    .B(_02916_),
    .X(_02918_));
 sky130_fd_sc_hd__xnor2_1 _09831_ (.A(_02878_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__a21o_1 _09832_ (.A1(_02700_),
    .A2(_02702_),
    .B1(_02706_),
    .X(_02920_));
 sky130_fd_sc_hd__o22a_1 _09833_ (.A1(net48),
    .A2(net77),
    .B1(net72),
    .B2(net46),
    .X(_02921_));
 sky130_fd_sc_hd__xnor2_2 _09834_ (.A(net97),
    .B(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__a22o_1 _09835_ (.A1(net31),
    .A2(_00348_),
    .B1(_00354_),
    .B2(net29),
    .X(_02923_));
 sky130_fd_sc_hd__xnor2_2 _09836_ (.A(net49),
    .B(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__nand2_1 _09837_ (.A(_02922_),
    .B(_02924_),
    .Y(_02925_));
 sky130_fd_sc_hd__or2_1 _09838_ (.A(_02922_),
    .B(_02924_),
    .X(_02926_));
 sky130_fd_sc_hd__nand2_1 _09839_ (.A(_02925_),
    .B(_02926_),
    .Y(_02927_));
 sky130_fd_sc_hd__a21bo_1 _09840_ (.A1(_02766_),
    .A2(_02771_),
    .B1_N(_02770_),
    .X(_02928_));
 sky130_fd_sc_hd__and3_1 _09841_ (.A(_02925_),
    .B(_02926_),
    .C(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__xnor2_2 _09842_ (.A(_02927_),
    .B(_02928_),
    .Y(_02930_));
 sky130_fd_sc_hd__xnor2_1 _09843_ (.A(_02920_),
    .B(_02930_),
    .Y(_02931_));
 sky130_fd_sc_hd__nor2_1 _09844_ (.A(_02919_),
    .B(_02931_),
    .Y(_02932_));
 sky130_fd_sc_hd__nand2_1 _09845_ (.A(_02919_),
    .B(_02931_),
    .Y(_02933_));
 sky130_fd_sc_hd__and2b_1 _09846_ (.A_N(_02932_),
    .B(_02933_),
    .X(_02934_));
 sky130_fd_sc_hd__xor2_4 _09847_ (.A(_02872_),
    .B(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__a21o_1 _09848_ (.A1(_02712_),
    .A2(_02777_),
    .B1(_02776_),
    .X(_02936_));
 sky130_fd_sc_hd__a21o_1 _09849_ (.A1(_02697_),
    .A2(_02711_),
    .B1(_02709_),
    .X(_02937_));
 sky130_fd_sc_hd__nand2_1 _09850_ (.A(_02724_),
    .B(_02726_),
    .Y(_02938_));
 sky130_fd_sc_hd__a21oi_2 _09851_ (.A1(_02735_),
    .A2(_02774_),
    .B1(_02773_),
    .Y(_02939_));
 sky130_fd_sc_hd__a21oi_1 _09852_ (.A1(_02724_),
    .A2(_02726_),
    .B1(_02939_),
    .Y(_02940_));
 sky130_fd_sc_hd__xnor2_2 _09853_ (.A(_02938_),
    .B(_02939_),
    .Y(_02941_));
 sky130_fd_sc_hd__xnor2_2 _09854_ (.A(_02937_),
    .B(_02941_),
    .Y(_02942_));
 sky130_fd_sc_hd__a21boi_2 _09855_ (.A1(_02781_),
    .A2(_02785_),
    .B1_N(_02784_),
    .Y(_02943_));
 sky130_fd_sc_hd__xnor2_1 _09856_ (.A(_02942_),
    .B(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__nand2b_1 _09857_ (.A_N(_02944_),
    .B(_02936_),
    .Y(_02945_));
 sky130_fd_sc_hd__xnor2_2 _09858_ (.A(_02936_),
    .B(_02944_),
    .Y(_02946_));
 sky130_fd_sc_hd__and2_1 _09859_ (.A(_02935_),
    .B(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__xor2_4 _09860_ (.A(_02935_),
    .B(_02946_),
    .X(_02948_));
 sky130_fd_sc_hd__xnor2_4 _09861_ (.A(_02856_),
    .B(_02948_),
    .Y(_02949_));
 sky130_fd_sc_hd__xnor2_4 _09862_ (.A(_02855_),
    .B(_02949_),
    .Y(_02950_));
 sky130_fd_sc_hd__or4_1 _09863_ (.A(_02238_),
    .B(_02462_),
    .C(_02638_),
    .D(_02796_),
    .X(_02951_));
 sky130_fd_sc_hd__a21o_1 _09864_ (.A1(_02133_),
    .A2(_02135_),
    .B1(_02951_),
    .X(_02952_));
 sky130_fd_sc_hd__a21o_1 _09865_ (.A1(_02636_),
    .A2(_02794_),
    .B1(_02795_),
    .X(_02953_));
 sky130_fd_sc_hd__o31a_2 _09866_ (.A1(_02638_),
    .A2(_02641_),
    .A3(_02796_),
    .B1(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__a21oi_1 _09867_ (.A1(_02952_),
    .A2(_02954_),
    .B1(_02950_),
    .Y(_02955_));
 sky130_fd_sc_hd__and3_1 _09868_ (.A(_02950_),
    .B(_02952_),
    .C(_02954_),
    .X(_02956_));
 sky130_fd_sc_hd__or2_2 _09869_ (.A(_02955_),
    .B(_02956_),
    .X(_02957_));
 sky130_fd_sc_hd__o21ai_1 _09870_ (.A1(_02854_),
    .A2(_02957_),
    .B1(net200),
    .Y(_02958_));
 sky130_fd_sc_hd__a21oi_1 _09871_ (.A1(_02854_),
    .A2(_02957_),
    .B1(_02958_),
    .Y(_02959_));
 sky130_fd_sc_hd__a21oi_1 _09872_ (.A1(net163),
    .A2(_01810_),
    .B1(_01811_),
    .Y(_02960_));
 sky130_fd_sc_hd__a311oi_1 _09873_ (.A1(net163),
    .A2(_01810_),
    .A3(_01811_),
    .B1(_02324_),
    .C1(_02960_),
    .Y(_02961_));
 sky130_fd_sc_hd__o31ai_2 _09874_ (.A1(_06348_),
    .A2(_06355_),
    .A3(_02831_),
    .B1(_06349_),
    .Y(_02962_));
 sky130_fd_sc_hd__nand2_1 _09875_ (.A(net286),
    .B(_02962_),
    .Y(_02963_));
 sky130_fd_sc_hd__o21a_1 _09876_ (.A1(net286),
    .A2(_06372_),
    .B1(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__a21oi_1 _09877_ (.A1(_06344_),
    .A2(_02964_),
    .B1(net236),
    .Y(_02965_));
 sky130_fd_sc_hd__o21a_1 _09878_ (.A1(_06344_),
    .A2(_02964_),
    .B1(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__o21ai_2 _09879_ (.A1(net223),
    .A2(_02815_),
    .B1(_02342_),
    .Y(_02967_));
 sky130_fd_sc_hd__a21boi_4 _09880_ (.A1(net225),
    .A2(_02967_),
    .B1_N(_02335_),
    .Y(_02968_));
 sky130_fd_sc_hd__mux2_1 _09881_ (.A0(_02259_),
    .A1(_02267_),
    .S(net219),
    .X(_02969_));
 sky130_fd_sc_hd__mux2_1 _09882_ (.A0(_02274_),
    .A1(_02298_),
    .S(net219),
    .X(_02970_));
 sky130_fd_sc_hd__mux2_1 _09883_ (.A0(_02969_),
    .A1(_02970_),
    .S(net222),
    .X(_02971_));
 sky130_fd_sc_hd__mux2_1 _09884_ (.A0(_02283_),
    .A1(_02305_),
    .S(_06352_),
    .X(_02972_));
 sky130_fd_sc_hd__mux2_1 _09885_ (.A0(_02828_),
    .A1(_02972_),
    .S(net224),
    .X(_02973_));
 sky130_fd_sc_hd__mux2_2 _09886_ (.A0(_02971_),
    .A1(_02973_),
    .S(net226),
    .X(_02974_));
 sky130_fd_sc_hd__a21o_1 _09887_ (.A1(net229),
    .A2(net210),
    .B1(_02313_),
    .X(_02975_));
 sky130_fd_sc_hd__or4_2 _09888_ (.A(\div_res[3] ),
    .B(\div_res[2] ),
    .C(\div_res[1] ),
    .D(\div_res[0] ),
    .X(_02976_));
 sky130_fd_sc_hd__a21oi_1 _09889_ (.A1(net167),
    .A2(_02976_),
    .B1(\div_res[4] ),
    .Y(_02977_));
 sky130_fd_sc_hd__a31o_1 _09890_ (.A1(\div_res[4] ),
    .A2(net163),
    .A3(_02976_),
    .B1(net195),
    .X(_02978_));
 sky130_fd_sc_hd__or4_2 _09891_ (.A(\div_shifter[35] ),
    .B(\div_shifter[34] ),
    .C(\div_shifter[33] ),
    .D(\div_shifter[32] ),
    .X(_02979_));
 sky130_fd_sc_hd__a21oi_1 _09892_ (.A1(net235),
    .A2(_02979_),
    .B1(\div_shifter[36] ),
    .Y(_02980_));
 sky130_fd_sc_hd__a31o_1 _09893_ (.A1(\div_shifter[36] ),
    .A2(net235),
    .A3(_02979_),
    .B1(net193),
    .X(_02981_));
 sky130_fd_sc_hd__a2bb2o_1 _09894_ (.A1_N(_02980_),
    .A2_N(_02981_),
    .B1(net228),
    .B2(net241),
    .X(_02982_));
 sky130_fd_sc_hd__o21a_1 _09895_ (.A1(_02822_),
    .A2(_02823_),
    .B1(_02824_),
    .X(_02983_));
 sky130_fd_sc_hd__nor2_1 _09896_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .Y(_02984_));
 sky130_fd_sc_hd__nand2_1 _09897_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .Y(_02985_));
 sky130_fd_sc_hd__nand2b_1 _09898_ (.A_N(_02984_),
    .B(_02985_),
    .Y(_02986_));
 sky130_fd_sc_hd__xor2_2 _09899_ (.A(_02983_),
    .B(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__a32o_1 _09900_ (.A1(net250),
    .A2(net210),
    .A3(_02987_),
    .B1(_02315_),
    .B2(_06342_),
    .X(_02988_));
 sky130_fd_sc_hd__a311o_1 _09901_ (.A1(reg1_val[4]),
    .A2(net228),
    .A3(_02325_),
    .B1(_02982_),
    .C1(_02988_),
    .X(_02989_));
 sky130_fd_sc_hd__o21ba_1 _09902_ (.A1(_06344_),
    .A2(net197),
    .B1_N(_02989_),
    .X(_02990_));
 sky130_fd_sc_hd__o21ai_1 _09903_ (.A1(_02977_),
    .A2(_02978_),
    .B1(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hd__a221o_1 _09904_ (.A1(net179),
    .A2(_02968_),
    .B1(_02974_),
    .B2(_02975_),
    .C1(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__o41a_1 _09905_ (.A1(_02959_),
    .A2(_02961_),
    .A3(_02966_),
    .A4(_02992_),
    .B1(net247),
    .X(_02993_));
 sky130_fd_sc_hd__nand2_1 _09906_ (.A(curr_PC[4]),
    .B(_02851_),
    .Y(_02994_));
 sky130_fd_sc_hd__or2_1 _09907_ (.A(curr_PC[4]),
    .B(_02851_),
    .X(_02995_));
 sky130_fd_sc_hd__a31o_4 _09908_ (.A1(net248),
    .A2(_02994_),
    .A3(_02995_),
    .B1(_02993_),
    .X(dest_val[4]));
 sky130_fd_sc_hd__nand2_1 _09909_ (.A(_02853_),
    .B(_02957_),
    .Y(_02996_));
 sky130_fd_sc_hd__nand2_1 _09910_ (.A(net163),
    .B(_02996_),
    .Y(_02997_));
 sky130_fd_sc_hd__a21oi_4 _09911_ (.A1(_02856_),
    .A2(_02948_),
    .B1(_02947_),
    .Y(_02998_));
 sky130_fd_sc_hd__o21ai_4 _09912_ (.A1(_02942_),
    .A2(_02943_),
    .B1(_02945_),
    .Y(_02999_));
 sky130_fd_sc_hd__a21o_1 _09913_ (.A1(_02888_),
    .A2(_02908_),
    .B1(_02906_),
    .X(_03000_));
 sky130_fd_sc_hd__a22o_1 _09914_ (.A1(net44),
    .A2(net116),
    .B1(_00324_),
    .B2(net42),
    .X(_03001_));
 sky130_fd_sc_hd__xor2_1 _09915_ (.A(net92),
    .B(_03001_),
    .X(_03002_));
 sky130_fd_sc_hd__o22a_1 _09916_ (.A1(net47),
    .A2(net81),
    .B1(net77),
    .B2(net45),
    .X(_03003_));
 sky130_fd_sc_hd__xnor2_1 _09917_ (.A(net96),
    .B(_03003_),
    .Y(_03004_));
 sky130_fd_sc_hd__and2_1 _09918_ (.A(_03002_),
    .B(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__nor2_1 _09919_ (.A(_03002_),
    .B(_03004_),
    .Y(_03006_));
 sky130_fd_sc_hd__nor2_1 _09920_ (.A(_03005_),
    .B(_03006_),
    .Y(_03007_));
 sky130_fd_sc_hd__a22o_1 _09921_ (.A1(net37),
    .A2(net118),
    .B1(_00366_),
    .B2(net39),
    .X(_03008_));
 sky130_fd_sc_hd__xor2_1 _09922_ (.A(net91),
    .B(_03008_),
    .X(_03009_));
 sky130_fd_sc_hd__xor2_1 _09923_ (.A(_03007_),
    .B(_03009_),
    .X(_03010_));
 sky130_fd_sc_hd__o21bai_2 _09924_ (.A1(_02874_),
    .A2(_02875_),
    .B1_N(_02877_),
    .Y(_03011_));
 sky130_fd_sc_hd__xnor2_1 _09925_ (.A(_03010_),
    .B(_03011_),
    .Y(_03012_));
 sky130_fd_sc_hd__and2b_1 _09926_ (.A_N(_03012_),
    .B(_03000_),
    .X(_03013_));
 sky130_fd_sc_hd__and2b_1 _09927_ (.A_N(_03000_),
    .B(_03012_),
    .X(_03014_));
 sky130_fd_sc_hd__nor2_2 _09928_ (.A(_03013_),
    .B(_03014_),
    .Y(_03015_));
 sky130_fd_sc_hd__o21ai_1 _09929_ (.A1(_02882_),
    .A2(_02884_),
    .B1(_02886_),
    .Y(_03016_));
 sky130_fd_sc_hd__o21ba_1 _09930_ (.A1(_02894_),
    .A2(_02898_),
    .B1_N(_02904_),
    .X(_03017_));
 sky130_fd_sc_hd__or3b_1 _09931_ (.A(_02894_),
    .B(_02898_),
    .C_N(_02904_),
    .X(_03018_));
 sky130_fd_sc_hd__nand2b_1 _09932_ (.A_N(_03017_),
    .B(_03018_),
    .Y(_03019_));
 sky130_fd_sc_hd__xor2_1 _09933_ (.A(_03016_),
    .B(_03019_),
    .X(_03020_));
 sky130_fd_sc_hd__nor2_1 _09934_ (.A(net130),
    .B(net21),
    .Y(_03021_));
 sky130_fd_sc_hd__a32o_1 _09935_ (.A1(_00308_),
    .A2(_00686_),
    .A3(_00687_),
    .B1(_00330_),
    .B2(_00452_),
    .X(_03022_));
 sky130_fd_sc_hd__xnor2_1 _09936_ (.A(net71),
    .B(_03022_),
    .Y(_03023_));
 sky130_fd_sc_hd__nand2_1 _09937_ (.A(_03021_),
    .B(_03023_),
    .Y(_03024_));
 sky130_fd_sc_hd__or2_1 _09938_ (.A(_03021_),
    .B(_03023_),
    .X(_03025_));
 sky130_fd_sc_hd__nand2_1 _09939_ (.A(_03024_),
    .B(_03025_),
    .Y(_03026_));
 sky130_fd_sc_hd__o22a_1 _09940_ (.A1(_00313_),
    .A2(net11),
    .B1(net6),
    .B2(net108),
    .X(_03027_));
 sky130_fd_sc_hd__xnor2_2 _09941_ (.A(net21),
    .B(_03027_),
    .Y(_03028_));
 sky130_fd_sc_hd__xor2_2 _09942_ (.A(_03026_),
    .B(_03028_),
    .X(_03029_));
 sky130_fd_sc_hd__o22a_1 _09943_ (.A1(net146),
    .A2(net13),
    .B1(net8),
    .B2(net148),
    .X(_03030_));
 sky130_fd_sc_hd__xnor2_2 _09944_ (.A(net202),
    .B(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__o22a_1 _09945_ (.A1(net132),
    .A2(net17),
    .B1(net14),
    .B2(net134),
    .X(_03032_));
 sky130_fd_sc_hd__xnor2_2 _09946_ (.A(net181),
    .B(_03032_),
    .Y(_03033_));
 sky130_fd_sc_hd__xnor2_2 _09947_ (.A(net207),
    .B(_03033_),
    .Y(_03034_));
 sky130_fd_sc_hd__nand2b_1 _09948_ (.A_N(_03031_),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__xnor2_2 _09949_ (.A(_03031_),
    .B(_03034_),
    .Y(_03036_));
 sky130_fd_sc_hd__o22a_2 _09950_ (.A1(net65),
    .A2(net86),
    .B1(net82),
    .B2(net59),
    .X(_03037_));
 sky130_fd_sc_hd__xnor2_4 _09951_ (.A(net137),
    .B(_03037_),
    .Y(_03038_));
 sky130_fd_sc_hd__o22a_2 _09952_ (.A1(net56),
    .A2(net107),
    .B1(net104),
    .B2(net67),
    .X(_03039_));
 sky130_fd_sc_hd__xnor2_4 _09953_ (.A(_00341_),
    .B(_03039_),
    .Y(_03040_));
 sky130_fd_sc_hd__o22a_2 _09954_ (.A1(net58),
    .A2(net78),
    .B1(net74),
    .B2(net64),
    .X(_03041_));
 sky130_fd_sc_hd__xnor2_4 _09955_ (.A(net122),
    .B(_03041_),
    .Y(_03042_));
 sky130_fd_sc_hd__nor2_1 _09956_ (.A(_03040_),
    .B(_03042_),
    .Y(_03043_));
 sky130_fd_sc_hd__xnor2_4 _09957_ (.A(_03040_),
    .B(_03042_),
    .Y(_03044_));
 sky130_fd_sc_hd__nor2_1 _09958_ (.A(_03038_),
    .B(_03044_),
    .Y(_03045_));
 sky130_fd_sc_hd__xor2_4 _09959_ (.A(_03038_),
    .B(_03044_),
    .X(_03046_));
 sky130_fd_sc_hd__xnor2_2 _09960_ (.A(_02925_),
    .B(_03046_),
    .Y(_03047_));
 sky130_fd_sc_hd__xor2_1 _09961_ (.A(_03036_),
    .B(_03047_),
    .X(_03048_));
 sky130_fd_sc_hd__and2_1 _09962_ (.A(_03029_),
    .B(_03048_),
    .X(_03049_));
 sky130_fd_sc_hd__xnor2_1 _09963_ (.A(_03029_),
    .B(_03048_),
    .Y(_03050_));
 sky130_fd_sc_hd__nor2_1 _09964_ (.A(_03020_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__and2_1 _09965_ (.A(_03020_),
    .B(_03050_),
    .X(_03052_));
 sky130_fd_sc_hd__or2_1 _09966_ (.A(_03051_),
    .B(_03052_),
    .X(_03053_));
 sky130_fd_sc_hd__a21o_1 _09967_ (.A1(_02865_),
    .A2(_02867_),
    .B1(_02862_),
    .X(_03054_));
 sky130_fd_sc_hd__o22a_1 _09968_ (.A1(net61),
    .A2(net36),
    .B1(net33),
    .B2(net53),
    .X(_03055_));
 sky130_fd_sc_hd__xnor2_2 _09969_ (.A(net125),
    .B(_03055_),
    .Y(_03056_));
 sky130_fd_sc_hd__a22o_1 _09970_ (.A1(_00189_),
    .A2(net32),
    .B1(net30),
    .B2(_00348_),
    .X(_03057_));
 sky130_fd_sc_hd__xnor2_2 _09971_ (.A(net50),
    .B(_03057_),
    .Y(_03058_));
 sky130_fd_sc_hd__and2_1 _09972_ (.A(_03056_),
    .B(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__xor2_2 _09973_ (.A(_03056_),
    .B(_03058_),
    .X(_03060_));
 sky130_fd_sc_hd__o22a_1 _09974_ (.A1(net52),
    .A2(net28),
    .B1(net26),
    .B2(net101),
    .X(_03061_));
 sky130_fd_sc_hd__xnor2_2 _09975_ (.A(net89),
    .B(_03061_),
    .Y(_03062_));
 sky130_fd_sc_hd__xnor2_2 _09976_ (.A(_03060_),
    .B(_03062_),
    .Y(_03063_));
 sky130_fd_sc_hd__a21oi_2 _09977_ (.A1(_02910_),
    .A2(_02915_),
    .B1(_02914_),
    .Y(_03064_));
 sky130_fd_sc_hd__nor2_1 _09978_ (.A(_03063_),
    .B(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__xor2_2 _09979_ (.A(_03063_),
    .B(_03064_),
    .X(_03066_));
 sky130_fd_sc_hd__xnor2_1 _09980_ (.A(_03054_),
    .B(_03066_),
    .Y(_03067_));
 sky130_fd_sc_hd__nor2_1 _09981_ (.A(_03053_),
    .B(_03067_),
    .Y(_03068_));
 sky130_fd_sc_hd__nand2_1 _09982_ (.A(_03053_),
    .B(_03067_),
    .Y(_03069_));
 sky130_fd_sc_hd__and2b_1 _09983_ (.A_N(_03068_),
    .B(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__xor2_4 _09984_ (.A(_03015_),
    .B(_03070_),
    .X(_03071_));
 sky130_fd_sc_hd__a21o_1 _09985_ (.A1(_02872_),
    .A2(_02933_),
    .B1(_02932_),
    .X(_03072_));
 sky130_fd_sc_hd__a21o_1 _09986_ (.A1(_02937_),
    .A2(_02941_),
    .B1(_02940_),
    .X(_03073_));
 sky130_fd_sc_hd__a21o_2 _09987_ (.A1(_02857_),
    .A2(_02871_),
    .B1(_02869_),
    .X(_03074_));
 sky130_fd_sc_hd__a21oi_4 _09988_ (.A1(_02878_),
    .A2(_02918_),
    .B1(_02917_),
    .Y(_03075_));
 sky130_fd_sc_hd__a21oi_4 _09989_ (.A1(_02920_),
    .A2(_02930_),
    .B1(_02929_),
    .Y(_03076_));
 sky130_fd_sc_hd__nor2_1 _09990_ (.A(_03075_),
    .B(_03076_),
    .Y(_03077_));
 sky130_fd_sc_hd__xor2_4 _09991_ (.A(_03075_),
    .B(_03076_),
    .X(_03078_));
 sky130_fd_sc_hd__xor2_2 _09992_ (.A(_03074_),
    .B(_03078_),
    .X(_03079_));
 sky130_fd_sc_hd__xnor2_2 _09993_ (.A(_03073_),
    .B(_03079_),
    .Y(_03080_));
 sky130_fd_sc_hd__nand2b_1 _09994_ (.A_N(_03080_),
    .B(_03072_),
    .Y(_03081_));
 sky130_fd_sc_hd__xnor2_2 _09995_ (.A(_03072_),
    .B(_03080_),
    .Y(_03082_));
 sky130_fd_sc_hd__and2_1 _09996_ (.A(_03071_),
    .B(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__xor2_4 _09997_ (.A(_03071_),
    .B(_03082_),
    .X(_03084_));
 sky130_fd_sc_hd__xnor2_4 _09998_ (.A(_02999_),
    .B(_03084_),
    .Y(_03085_));
 sky130_fd_sc_hd__xnor2_4 _09999_ (.A(_02998_),
    .B(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__o22a_1 _10000_ (.A1(_02695_),
    .A2(_02793_),
    .B1(_02855_),
    .B2(_02949_),
    .X(_03087_));
 sky130_fd_sc_hd__a21oi_1 _10001_ (.A1(_02855_),
    .A2(_02949_),
    .B1(_03087_),
    .Y(_03088_));
 sky130_fd_sc_hd__nor2_1 _10002_ (.A(_02796_),
    .B(_02950_),
    .Y(_03089_));
 sky130_fd_sc_hd__a21o_1 _10003_ (.A1(_02798_),
    .A2(_03089_),
    .B1(_03088_),
    .X(_03090_));
 sky130_fd_sc_hd__nor4_2 _10004_ (.A(_02462_),
    .B(_02638_),
    .C(_02796_),
    .D(_02950_),
    .Y(_03091_));
 sky130_fd_sc_hd__a21oi_4 _10005_ (.A1(_02466_),
    .A2(_03091_),
    .B1(_03090_),
    .Y(_03092_));
 sky130_fd_sc_hd__xnor2_4 _10006_ (.A(_03086_),
    .B(_03092_),
    .Y(_03093_));
 sky130_fd_sc_hd__o21ai_1 _10007_ (.A1(_02997_),
    .A2(_03093_),
    .B1(net200),
    .Y(_03094_));
 sky130_fd_sc_hd__a21oi_1 _10008_ (.A1(_02997_),
    .A2(_03093_),
    .B1(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__o21ai_1 _10009_ (.A1(net157),
    .A2(_01812_),
    .B1(_01813_),
    .Y(_03096_));
 sky130_fd_sc_hd__or3_1 _10010_ (.A(net157),
    .B(_01812_),
    .C(_01813_),
    .X(_03097_));
 sky130_fd_sc_hd__a21boi_1 _10011_ (.A1(_06342_),
    .A2(_02962_),
    .B1_N(_06343_),
    .Y(_03098_));
 sky130_fd_sc_hd__nor2_1 _10012_ (.A(net294),
    .B(_03098_),
    .Y(_03099_));
 sky130_fd_sc_hd__a21oi_1 _10013_ (.A1(net294),
    .A2(_06374_),
    .B1(_03099_),
    .Y(_03100_));
 sky130_fd_sc_hd__xnor2_1 _10014_ (.A(_06337_),
    .B(_03100_),
    .Y(_03101_));
 sky130_fd_sc_hd__o21ai_1 _10015_ (.A1(net223),
    .A2(_02661_),
    .B1(_02342_),
    .Y(_03102_));
 sky130_fd_sc_hd__a21boi_2 _10016_ (.A1(net225),
    .A2(_03102_),
    .B1_N(_02335_),
    .Y(_03103_));
 sky130_fd_sc_hd__mux2_1 _10017_ (.A0(_02475_),
    .A1(_02479_),
    .S(net220),
    .X(_03104_));
 sky130_fd_sc_hd__or2_1 _10018_ (.A(net220),
    .B(_02482_),
    .X(_03105_));
 sky130_fd_sc_hd__o21ai_1 _10019_ (.A1(_06352_),
    .A2(_02493_),
    .B1(_03105_),
    .Y(_03106_));
 sky130_fd_sc_hd__nand2_1 _10020_ (.A(net222),
    .B(_03106_),
    .Y(_03107_));
 sky130_fd_sc_hd__o211a_1 _10021_ (.A1(net222),
    .A2(_03104_),
    .B1(_03107_),
    .C1(net225),
    .X(_03108_));
 sky130_fd_sc_hd__or2_1 _10022_ (.A(net219),
    .B(_02496_),
    .X(_03109_));
 sky130_fd_sc_hd__o21ai_1 _10023_ (.A1(_06352_),
    .A2(_02487_),
    .B1(_03109_),
    .Y(_03110_));
 sky130_fd_sc_hd__or2_1 _10024_ (.A(net224),
    .B(_02648_),
    .X(_03111_));
 sky130_fd_sc_hd__o21ai_1 _10025_ (.A1(net223),
    .A2(_03110_),
    .B1(_03111_),
    .Y(_03112_));
 sky130_fd_sc_hd__a21o_1 _10026_ (.A1(net227),
    .A2(_03112_),
    .B1(_03108_),
    .X(_03113_));
 sky130_fd_sc_hd__o21ai_1 _10027_ (.A1(\div_res[4] ),
    .A2(_02976_),
    .B1(net162),
    .Y(_03114_));
 sky130_fd_sc_hd__xnor2_1 _10028_ (.A(\div_res[5] ),
    .B(_03114_),
    .Y(_03115_));
 sky130_fd_sc_hd__o21a_1 _10029_ (.A1(\div_shifter[36] ),
    .A2(_02979_),
    .B1(net235),
    .X(_03116_));
 sky130_fd_sc_hd__and2_1 _10030_ (.A(\div_shifter[37] ),
    .B(_03116_),
    .X(_03117_));
 sky130_fd_sc_hd__nor2_1 _10031_ (.A(\div_shifter[37] ),
    .B(_03116_),
    .Y(_03118_));
 sky130_fd_sc_hd__o32a_1 _10032_ (.A1(net193),
    .A2(_03117_),
    .A3(_03118_),
    .B1(net209),
    .B2(_06332_),
    .X(_03119_));
 sky130_fd_sc_hd__o221a_1 _10033_ (.A1(_06334_),
    .A2(net199),
    .B1(net196),
    .B2(_06336_),
    .C1(_03119_),
    .X(_03120_));
 sky130_fd_sc_hd__o21ai_1 _10034_ (.A1(_06338_),
    .A2(net197),
    .B1(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__o21a_1 _10035_ (.A1(_02983_),
    .A2(_02984_),
    .B1(_02985_),
    .X(_03122_));
 sky130_fd_sc_hd__nor2_1 _10036_ (.A(reg1_val[5]),
    .B(curr_PC[5]),
    .Y(_03123_));
 sky130_fd_sc_hd__nand2_1 _10037_ (.A(reg1_val[5]),
    .B(curr_PC[5]),
    .Y(_03124_));
 sky130_fd_sc_hd__and2b_1 _10038_ (.A_N(_03123_),
    .B(_03124_),
    .X(_03125_));
 sky130_fd_sc_hd__xnor2_1 _10039_ (.A(_03122_),
    .B(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__a31o_1 _10040_ (.A1(net250),
    .A2(net210),
    .A3(_03126_),
    .B1(_03121_),
    .X(_03127_));
 sky130_fd_sc_hd__a221o_1 _10041_ (.A1(_02975_),
    .A2(_03113_),
    .B1(_03115_),
    .B2(_02328_),
    .C1(_03127_),
    .X(_03128_));
 sky130_fd_sc_hd__a221o_1 _10042_ (.A1(_02317_),
    .A2(_03101_),
    .B1(_03103_),
    .B2(net179),
    .C1(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__a311o_1 _10043_ (.A1(_02323_),
    .A2(_03096_),
    .A3(_03097_),
    .B1(_03129_),
    .C1(_03095_),
    .X(_03130_));
 sky130_fd_sc_hd__a31o_1 _10044_ (.A1(curr_PC[3]),
    .A2(curr_PC[4]),
    .A3(_02532_),
    .B1(curr_PC[5]),
    .X(_03131_));
 sky130_fd_sc_hd__and3_1 _10045_ (.A(curr_PC[4]),
    .B(curr_PC[5]),
    .C(_02851_),
    .X(_03132_));
 sky130_fd_sc_hd__nor2_1 _10046_ (.A(net242),
    .B(_03132_),
    .Y(_03133_));
 sky130_fd_sc_hd__a22o_4 _10047_ (.A1(net242),
    .A2(_03130_),
    .B1(_03131_),
    .B2(_03133_),
    .X(dest_val[5]));
 sky130_fd_sc_hd__nand2b_1 _10048_ (.A_N(_02996_),
    .B(_03093_),
    .Y(_03134_));
 sky130_fd_sc_hd__nand2_1 _10049_ (.A(net163),
    .B(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__a21oi_4 _10050_ (.A1(_02999_),
    .A2(_03084_),
    .B1(_03083_),
    .Y(_03136_));
 sky130_fd_sc_hd__a21bo_2 _10051_ (.A1(_03073_),
    .A2(_03079_),
    .B1_N(_03081_),
    .X(_03137_));
 sky130_fd_sc_hd__o21ai_2 _10052_ (.A1(_06532_),
    .A2(_03033_),
    .B1(_03035_),
    .Y(_03138_));
 sky130_fd_sc_hd__o211a_1 _10053_ (.A1(_03043_),
    .A2(_03045_),
    .B1(_00374_),
    .C1(net22),
    .X(_03139_));
 sky130_fd_sc_hd__a211o_1 _10054_ (.A1(_00374_),
    .A2(net22),
    .B1(_03043_),
    .C1(_03045_),
    .X(_03140_));
 sky130_fd_sc_hd__and2b_1 _10055_ (.A_N(_03139_),
    .B(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__xnor2_2 _10056_ (.A(_03138_),
    .B(_03141_),
    .Y(_03142_));
 sky130_fd_sc_hd__o22a_1 _10057_ (.A1(net67),
    .A2(net86),
    .B1(net82),
    .B2(net66),
    .X(_03143_));
 sky130_fd_sc_hd__xnor2_2 _10058_ (.A(_00339_),
    .B(_03143_),
    .Y(_03144_));
 sky130_fd_sc_hd__o32a_1 _10059_ (.A1(_00390_),
    .A2(_00405_),
    .A3(_00407_),
    .B1(net104),
    .B2(net55),
    .X(_03145_));
 sky130_fd_sc_hd__xnor2_2 _10060_ (.A(_00341_),
    .B(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__o22a_1 _10061_ (.A1(net60),
    .A2(net78),
    .B1(net74),
    .B2(net58),
    .X(_03147_));
 sky130_fd_sc_hd__xnor2_2 _10062_ (.A(net122),
    .B(_03147_),
    .Y(_03148_));
 sky130_fd_sc_hd__nor2_1 _10063_ (.A(_03146_),
    .B(_03148_),
    .Y(_03149_));
 sky130_fd_sc_hd__nand2_1 _10064_ (.A(_03146_),
    .B(_03148_),
    .Y(_03150_));
 sky130_fd_sc_hd__xnor2_1 _10065_ (.A(_03146_),
    .B(_03148_),
    .Y(_03151_));
 sky130_fd_sc_hd__xnor2_2 _10066_ (.A(_03144_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__a21o_1 _10067_ (.A1(_03060_),
    .A2(_03062_),
    .B1(_03059_),
    .X(_03153_));
 sky130_fd_sc_hd__nand2_1 _10068_ (.A(_03152_),
    .B(_03153_),
    .Y(_03154_));
 sky130_fd_sc_hd__xor2_2 _10069_ (.A(_03152_),
    .B(_03153_),
    .X(_03155_));
 sky130_fd_sc_hd__o22a_1 _10070_ (.A1(net132),
    .A2(net14),
    .B1(net13),
    .B2(net134),
    .X(_03156_));
 sky130_fd_sc_hd__xnor2_1 _10071_ (.A(net182),
    .B(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__nor2_1 _10072_ (.A(_00158_),
    .B(net8),
    .Y(_03158_));
 sky130_fd_sc_hd__o22a_1 _10073_ (.A1(_00165_),
    .A2(net8),
    .B1(_03158_),
    .B2(net203),
    .X(_03159_));
 sky130_fd_sc_hd__and2_1 _10074_ (.A(_03157_),
    .B(_03159_),
    .X(_03160_));
 sky130_fd_sc_hd__nor2_1 _10075_ (.A(_03157_),
    .B(_03159_),
    .Y(_03161_));
 sky130_fd_sc_hd__or2_1 _10076_ (.A(_03160_),
    .B(_03161_),
    .X(_03162_));
 sky130_fd_sc_hd__xor2_2 _10077_ (.A(_03155_),
    .B(_03162_),
    .X(_03163_));
 sky130_fd_sc_hd__o22a_1 _10078_ (.A1(net112),
    .A2(net23),
    .B1(net15),
    .B2(net110),
    .X(_03164_));
 sky130_fd_sc_hd__xnor2_2 _10079_ (.A(net70),
    .B(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__a22o_1 _10080_ (.A1(_00308_),
    .A2(_01967_),
    .B1(_02082_),
    .B2(_00314_),
    .X(_03166_));
 sky130_fd_sc_hd__xnor2_2 _10081_ (.A(net21),
    .B(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__a22o_1 _10082_ (.A1(net43),
    .A2(net118),
    .B1(net116),
    .B2(net41),
    .X(_03168_));
 sky130_fd_sc_hd__xor2_2 _10083_ (.A(net92),
    .B(_03168_),
    .X(_03169_));
 sky130_fd_sc_hd__nand2_1 _10084_ (.A(_03167_),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__xnor2_2 _10085_ (.A(_03167_),
    .B(_03169_),
    .Y(_03171_));
 sky130_fd_sc_hd__xor2_2 _10086_ (.A(_03165_),
    .B(_03171_),
    .X(_03172_));
 sky130_fd_sc_hd__nand2_1 _10087_ (.A(_03163_),
    .B(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__xnor2_2 _10088_ (.A(_03163_),
    .B(_03172_),
    .Y(_03174_));
 sky130_fd_sc_hd__xor2_1 _10089_ (.A(_03142_),
    .B(_03174_),
    .X(_03175_));
 sky130_fd_sc_hd__a21o_1 _10090_ (.A1(_03007_),
    .A2(_03009_),
    .B1(_03005_),
    .X(_03176_));
 sky130_fd_sc_hd__o22a_1 _10091_ (.A1(net64),
    .A2(net36),
    .B1(net33),
    .B2(net61),
    .X(_03177_));
 sky130_fd_sc_hd__xnor2_1 _10092_ (.A(net125),
    .B(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__o22a_1 _10093_ (.A1(net54),
    .A2(net28),
    .B1(net26),
    .B2(net52),
    .X(_03179_));
 sky130_fd_sc_hd__xnor2_1 _10094_ (.A(net89),
    .B(_03179_),
    .Y(_03180_));
 sky130_fd_sc_hd__nand2_1 _10095_ (.A(_03178_),
    .B(_03180_),
    .Y(_03181_));
 sky130_fd_sc_hd__or2_1 _10096_ (.A(_03178_),
    .B(_03180_),
    .X(_03182_));
 sky130_fd_sc_hd__and2_1 _10097_ (.A(_03181_),
    .B(_03182_),
    .X(_03183_));
 sky130_fd_sc_hd__o21ai_2 _10098_ (.A1(_03026_),
    .A2(_03028_),
    .B1(_03024_),
    .Y(_03184_));
 sky130_fd_sc_hd__and2_1 _10099_ (.A(_03183_),
    .B(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__xnor2_1 _10100_ (.A(_03183_),
    .B(_03184_),
    .Y(_03186_));
 sky130_fd_sc_hd__and2b_1 _10101_ (.A_N(_03186_),
    .B(_03176_),
    .X(_03187_));
 sky130_fd_sc_hd__xnor2_1 _10102_ (.A(_03176_),
    .B(_03186_),
    .Y(_03188_));
 sky130_fd_sc_hd__nand2_1 _10103_ (.A(_03175_),
    .B(_03188_),
    .Y(_03189_));
 sky130_fd_sc_hd__or2_1 _10104_ (.A(_03175_),
    .B(_03188_),
    .X(_03190_));
 sky130_fd_sc_hd__and2_2 _10105_ (.A(_03189_),
    .B(_03190_),
    .X(_03191_));
 sky130_fd_sc_hd__a32oi_4 _10106_ (.A1(_02922_),
    .A2(_02924_),
    .A3(_03046_),
    .B1(_03047_),
    .B2(_03036_),
    .Y(_03192_));
 sky130_fd_sc_hd__a22o_1 _10107_ (.A1(net40),
    .A2(_00361_),
    .B1(_00366_),
    .B2(net38),
    .X(_03193_));
 sky130_fd_sc_hd__xor2_1 _10108_ (.A(_00245_),
    .B(_03193_),
    .X(_03194_));
 sky130_fd_sc_hd__a22o_1 _10109_ (.A1(net102),
    .A2(net32),
    .B1(net30),
    .B2(_00189_),
    .X(_03195_));
 sky130_fd_sc_hd__xnor2_1 _10110_ (.A(_00217_),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__and2_1 _10111_ (.A(_03194_),
    .B(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__nor2_1 _10112_ (.A(_03194_),
    .B(_03196_),
    .Y(_03198_));
 sky130_fd_sc_hd__nor2_2 _10113_ (.A(_03197_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__o22a_1 _10114_ (.A1(net47),
    .A2(net85),
    .B1(net81),
    .B2(net45),
    .X(_03200_));
 sky130_fd_sc_hd__xnor2_2 _10115_ (.A(net96),
    .B(_03200_),
    .Y(_03201_));
 sky130_fd_sc_hd__xor2_4 _10116_ (.A(_03199_),
    .B(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__a21o_1 _10117_ (.A1(_03016_),
    .A2(_03018_),
    .B1(_03017_),
    .X(_03203_));
 sky130_fd_sc_hd__xor2_4 _10118_ (.A(_03202_),
    .B(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__nand2b_1 _10119_ (.A_N(_03192_),
    .B(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__xnor2_4 _10120_ (.A(_03192_),
    .B(_03204_),
    .Y(_03206_));
 sky130_fd_sc_hd__xor2_4 _10121_ (.A(_03191_),
    .B(_03206_),
    .X(_03207_));
 sky130_fd_sc_hd__a21o_1 _10122_ (.A1(_03015_),
    .A2(_03069_),
    .B1(_03068_),
    .X(_03208_));
 sky130_fd_sc_hd__a21o_2 _10123_ (.A1(_03010_),
    .A2(_03011_),
    .B1(_03013_),
    .X(_03209_));
 sky130_fd_sc_hd__or2_2 _10124_ (.A(_03049_),
    .B(_03051_),
    .X(_03210_));
 sky130_fd_sc_hd__a21oi_4 _10125_ (.A1(_03054_),
    .A2(_03066_),
    .B1(_03065_),
    .Y(_03211_));
 sky130_fd_sc_hd__o21ba_1 _10126_ (.A1(_03049_),
    .A2(_03051_),
    .B1_N(_03211_),
    .X(_03212_));
 sky130_fd_sc_hd__xnor2_4 _10127_ (.A(_03210_),
    .B(_03211_),
    .Y(_03213_));
 sky130_fd_sc_hd__xnor2_4 _10128_ (.A(_03209_),
    .B(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__a21oi_4 _10129_ (.A1(_03074_),
    .A2(_03078_),
    .B1(_03077_),
    .Y(_03215_));
 sky130_fd_sc_hd__xnor2_2 _10130_ (.A(_03214_),
    .B(_03215_),
    .Y(_03216_));
 sky130_fd_sc_hd__and2b_1 _10131_ (.A_N(_03216_),
    .B(_03208_),
    .X(_03217_));
 sky130_fd_sc_hd__xnor2_2 _10132_ (.A(_03208_),
    .B(_03216_),
    .Y(_03218_));
 sky130_fd_sc_hd__and2_1 _10133_ (.A(_03207_),
    .B(_03218_),
    .X(_03219_));
 sky130_fd_sc_hd__xor2_4 _10134_ (.A(_03207_),
    .B(_03218_),
    .X(_03220_));
 sky130_fd_sc_hd__xnor2_4 _10135_ (.A(_03137_),
    .B(_03220_),
    .Y(_03221_));
 sky130_fd_sc_hd__xnor2_4 _10136_ (.A(_03136_),
    .B(_03221_),
    .Y(_03222_));
 sky130_fd_sc_hd__or4_4 _10137_ (.A(_02638_),
    .B(_02796_),
    .C(_02950_),
    .D(_03086_),
    .X(_03223_));
 sky130_fd_sc_hd__or3_1 _10138_ (.A(_02014_),
    .B(_02639_),
    .C(_03223_),
    .X(_03224_));
 sky130_fd_sc_hd__a21o_1 _10139_ (.A1(_02641_),
    .A2(_02642_),
    .B1(_03223_),
    .X(_03225_));
 sky130_fd_sc_hd__o22a_1 _10140_ (.A1(_02855_),
    .A2(_02949_),
    .B1(_02998_),
    .B2(_03085_),
    .X(_03226_));
 sky130_fd_sc_hd__a21oi_2 _10141_ (.A1(_02998_),
    .A2(_03085_),
    .B1(_03226_),
    .Y(_03227_));
 sky130_fd_sc_hd__a2111oi_2 _10142_ (.A1(_02636_),
    .A2(_02794_),
    .B1(_02795_),
    .C1(_02950_),
    .D1(_03086_),
    .Y(_03228_));
 sky130_fd_sc_hd__nor2_1 _10143_ (.A(_03227_),
    .B(_03228_),
    .Y(_03229_));
 sky130_fd_sc_hd__a31o_1 _10144_ (.A1(_03224_),
    .A2(_03225_),
    .A3(_03229_),
    .B1(_03222_),
    .X(_03230_));
 sky130_fd_sc_hd__o211ai_2 _10145_ (.A1(_02643_),
    .A2(_03223_),
    .B1(_03229_),
    .C1(_03222_),
    .Y(_03231_));
 sky130_fd_sc_hd__nand2_2 _10146_ (.A(_03230_),
    .B(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__inv_2 _10147_ (.A(_03232_),
    .Y(_03233_));
 sky130_fd_sc_hd__a21oi_1 _10148_ (.A1(_03135_),
    .A2(_03232_),
    .B1(_02242_),
    .Y(_03234_));
 sky130_fd_sc_hd__o21ai_1 _10149_ (.A1(_03135_),
    .A2(_03232_),
    .B1(_03234_),
    .Y(_03235_));
 sky130_fd_sc_hd__o21a_1 _10150_ (.A1(net157),
    .A2(_01814_),
    .B1(_01815_),
    .X(_03236_));
 sky130_fd_sc_hd__or3_1 _10151_ (.A(net157),
    .B(_01814_),
    .C(_01815_),
    .X(_03237_));
 sky130_fd_sc_hd__or3b_1 _10152_ (.A(_02324_),
    .B(_03236_),
    .C_N(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__o21ai_1 _10153_ (.A1(_06334_),
    .A2(_03098_),
    .B1(_06336_),
    .Y(_03239_));
 sky130_fd_sc_hd__mux2_1 _10154_ (.A0(_06376_),
    .A1(_03239_),
    .S(net285),
    .X(_03240_));
 sky130_fd_sc_hd__nand2_1 _10155_ (.A(_06329_),
    .B(_03240_),
    .Y(_03241_));
 sky130_fd_sc_hd__o21a_1 _10156_ (.A1(_06329_),
    .A2(_03240_),
    .B1(_02317_),
    .X(_03242_));
 sky130_fd_sc_hd__o21a_1 _10157_ (.A1(net223),
    .A2(_02490_),
    .B1(_02342_),
    .X(_03243_));
 sky130_fd_sc_hd__o21ai_2 _10158_ (.A1(net226),
    .A2(_03243_),
    .B1(_02335_),
    .Y(_03244_));
 sky130_fd_sc_hd__nor2_1 _10159_ (.A(net177),
    .B(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__mux2_1 _10160_ (.A0(_02654_),
    .A1(_02656_),
    .S(net219),
    .X(_03246_));
 sky130_fd_sc_hd__mux2_1 _10161_ (.A0(_02657_),
    .A1(_02662_),
    .S(net219),
    .X(_03247_));
 sky130_fd_sc_hd__mux2_1 _10162_ (.A0(_03246_),
    .A1(_03247_),
    .S(net222),
    .X(_03248_));
 sky130_fd_sc_hd__mux2_1 _10163_ (.A0(_02660_),
    .A1(_02663_),
    .S(_06352_),
    .X(_03249_));
 sky130_fd_sc_hd__mux2_1 _10164_ (.A0(_02527_),
    .A1(_03249_),
    .S(net224),
    .X(_03250_));
 sky130_fd_sc_hd__mux2_2 _10165_ (.A0(_03248_),
    .A1(_03250_),
    .S(net227),
    .X(_03251_));
 sky130_fd_sc_hd__or3_1 _10166_ (.A(\div_res[5] ),
    .B(\div_res[4] ),
    .C(_02976_),
    .X(_03252_));
 sky130_fd_sc_hd__a21oi_1 _10167_ (.A1(net162),
    .A2(_03252_),
    .B1(\div_res[6] ),
    .Y(_03253_));
 sky130_fd_sc_hd__a31o_1 _10168_ (.A1(\div_res[6] ),
    .A2(net162),
    .A3(_03252_),
    .B1(net195),
    .X(_03254_));
 sky130_fd_sc_hd__nor2_1 _10169_ (.A(_03253_),
    .B(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hd__or3_1 _10170_ (.A(\div_shifter[37] ),
    .B(\div_shifter[36] ),
    .C(_02979_),
    .X(_03256_));
 sky130_fd_sc_hd__a21oi_1 _10171_ (.A1(net235),
    .A2(_03256_),
    .B1(\div_shifter[38] ),
    .Y(_03257_));
 sky130_fd_sc_hd__a311oi_1 _10172_ (.A1(\div_shifter[38] ),
    .A2(net235),
    .A3(_03256_),
    .B1(_03257_),
    .C1(net193),
    .Y(_03258_));
 sky130_fd_sc_hd__a221o_1 _10173_ (.A1(_06325_),
    .A2(net241),
    .B1(_02325_),
    .B2(_06327_),
    .C1(_03258_),
    .X(_03259_));
 sky130_fd_sc_hd__a221o_1 _10174_ (.A1(_06326_),
    .A2(_02315_),
    .B1(_02319_),
    .B2(_06329_),
    .C1(_03259_),
    .X(_03260_));
 sky130_fd_sc_hd__o21a_1 _10175_ (.A1(_03122_),
    .A2(_03123_),
    .B1(_03124_),
    .X(_03261_));
 sky130_fd_sc_hd__nor2_1 _10176_ (.A(reg1_val[6]),
    .B(curr_PC[6]),
    .Y(_03262_));
 sky130_fd_sc_hd__nand2_1 _10177_ (.A(reg1_val[6]),
    .B(curr_PC[6]),
    .Y(_03263_));
 sky130_fd_sc_hd__and2b_1 _10178_ (.A_N(_03262_),
    .B(_03263_),
    .X(_03264_));
 sky130_fd_sc_hd__xnor2_1 _10179_ (.A(_03261_),
    .B(_03264_),
    .Y(_03265_));
 sky130_fd_sc_hd__a311o_1 _10180_ (.A1(_06330_),
    .A2(net210),
    .A3(_03265_),
    .B1(_03260_),
    .C1(_03255_),
    .X(_03266_));
 sky130_fd_sc_hd__a211o_1 _10181_ (.A1(_02975_),
    .A2(_03251_),
    .B1(_03266_),
    .C1(_03245_),
    .X(_03267_));
 sky130_fd_sc_hd__a21oi_1 _10182_ (.A1(_03241_),
    .A2(_03242_),
    .B1(_03267_),
    .Y(_03268_));
 sky130_fd_sc_hd__a31o_1 _10183_ (.A1(_03235_),
    .A2(_03238_),
    .A3(_03268_),
    .B1(net248),
    .X(_03269_));
 sky130_fd_sc_hd__and2_2 _10184_ (.A(curr_PC[6]),
    .B(_03132_),
    .X(_03270_));
 sky130_fd_sc_hd__o21ai_2 _10185_ (.A1(curr_PC[6]),
    .A2(_03132_),
    .B1(net248),
    .Y(_03271_));
 sky130_fd_sc_hd__o21ai_4 _10186_ (.A1(_03270_),
    .A2(_03271_),
    .B1(_03269_),
    .Y(dest_val[6]));
 sky130_fd_sc_hd__o21a_1 _10187_ (.A1(_03134_),
    .A2(_03233_),
    .B1(net163),
    .X(_03272_));
 sky130_fd_sc_hd__a21oi_4 _10188_ (.A1(_03137_),
    .A2(_03220_),
    .B1(_03219_),
    .Y(_03273_));
 sky130_fd_sc_hd__o21bai_4 _10189_ (.A1(_03214_),
    .A2(_03215_),
    .B1_N(_03217_),
    .Y(_03274_));
 sky130_fd_sc_hd__a21bo_2 _10190_ (.A1(_03155_),
    .A2(_03162_),
    .B1_N(_03154_),
    .X(_03275_));
 sky130_fd_sc_hd__a21o_2 _10191_ (.A1(_03138_),
    .A2(_03140_),
    .B1(_03139_),
    .X(_03276_));
 sky130_fd_sc_hd__o22a_1 _10192_ (.A1(net99),
    .A2(net47),
    .B1(net45),
    .B2(net85),
    .X(_03277_));
 sky130_fd_sc_hd__xnor2_1 _10193_ (.A(net96),
    .B(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__o22a_1 _10194_ (.A1(net62),
    .A2(net28),
    .B1(net26),
    .B2(net54),
    .X(_03279_));
 sky130_fd_sc_hd__xnor2_1 _10195_ (.A(net89),
    .B(_03279_),
    .Y(_03280_));
 sky130_fd_sc_hd__and2_1 _10196_ (.A(_03278_),
    .B(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__nor2_1 _10197_ (.A(_03278_),
    .B(_03280_),
    .Y(_03282_));
 sky130_fd_sc_hd__nor2_2 _10198_ (.A(_03281_),
    .B(_03282_),
    .Y(_03283_));
 sky130_fd_sc_hd__a22o_2 _10199_ (.A1(_00172_),
    .A2(_00305_),
    .B1(net30),
    .B2(net102),
    .X(_03284_));
 sky130_fd_sc_hd__xnor2_4 _10200_ (.A(_00217_),
    .B(_03284_),
    .Y(_03285_));
 sky130_fd_sc_hd__xnor2_4 _10201_ (.A(_03283_),
    .B(_03285_),
    .Y(_03286_));
 sky130_fd_sc_hd__and2b_1 _10202_ (.A_N(_03286_),
    .B(_03276_),
    .X(_03287_));
 sky130_fd_sc_hd__xnor2_4 _10203_ (.A(_03276_),
    .B(_03286_),
    .Y(_03288_));
 sky130_fd_sc_hd__xnor2_4 _10204_ (.A(_03275_),
    .B(_03288_),
    .Y(_03289_));
 sky130_fd_sc_hd__a21oi_1 _10205_ (.A1(_03199_),
    .A2(_03201_),
    .B1(_03197_),
    .Y(_03290_));
 sky130_fd_sc_hd__o22a_1 _10206_ (.A1(net56),
    .A2(net86),
    .B1(net82),
    .B2(net67),
    .X(_03291_));
 sky130_fd_sc_hd__xnor2_1 _10207_ (.A(net138),
    .B(_03291_),
    .Y(_03292_));
 sky130_fd_sc_hd__o22a_1 _10208_ (.A1(net57),
    .A2(net36),
    .B1(net34),
    .B2(net63),
    .X(_03293_));
 sky130_fd_sc_hd__xnor2_1 _10209_ (.A(_00276_),
    .B(_03293_),
    .Y(_03294_));
 sky130_fd_sc_hd__nor2_1 _10210_ (.A(_03292_),
    .B(_03294_),
    .Y(_03295_));
 sky130_fd_sc_hd__and2_1 _10211_ (.A(_03292_),
    .B(_03294_),
    .X(_03296_));
 sky130_fd_sc_hd__or2_1 _10212_ (.A(_03295_),
    .B(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__o22a_1 _10213_ (.A1(net65),
    .A2(net78),
    .B1(net74),
    .B2(net59),
    .X(_03298_));
 sky130_fd_sc_hd__xnor2_1 _10214_ (.A(net122),
    .B(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__xnor2_1 _10215_ (.A(_03297_),
    .B(_03299_),
    .Y(_03300_));
 sky130_fd_sc_hd__o21a_1 _10216_ (.A1(_03165_),
    .A2(_03171_),
    .B1(_03170_),
    .X(_03301_));
 sky130_fd_sc_hd__nor2_1 _10217_ (.A(_03300_),
    .B(_03301_),
    .Y(_03302_));
 sky130_fd_sc_hd__xor2_1 _10218_ (.A(_03300_),
    .B(_03301_),
    .X(_03303_));
 sky130_fd_sc_hd__and2b_1 _10219_ (.A_N(_03290_),
    .B(_03303_),
    .X(_03304_));
 sky130_fd_sc_hd__xnor2_1 _10220_ (.A(_03290_),
    .B(_03303_),
    .Y(_03305_));
 sky130_fd_sc_hd__o22a_1 _10221_ (.A1(net110),
    .A2(net11),
    .B1(net6),
    .B2(net115),
    .X(_03306_));
 sky130_fd_sc_hd__xnor2_1 _10222_ (.A(net21),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__nor2_1 _10223_ (.A(_03160_),
    .B(_03307_),
    .Y(_03308_));
 sky130_fd_sc_hd__xor2_1 _10224_ (.A(_03160_),
    .B(_03307_),
    .X(_03309_));
 sky130_fd_sc_hd__and3_1 _10225_ (.A(_00314_),
    .B(net22),
    .C(_03309_),
    .X(_03310_));
 sky130_fd_sc_hd__a21oi_1 _10226_ (.A1(_00314_),
    .A2(net22),
    .B1(_03309_),
    .Y(_03311_));
 sky130_fd_sc_hd__or2_1 _10227_ (.A(_03310_),
    .B(_03311_),
    .X(_03312_));
 sky130_fd_sc_hd__a32o_1 _10228_ (.A1(_00324_),
    .A2(_00686_),
    .A3(_00687_),
    .B1(_00452_),
    .B2(net116),
    .X(_03313_));
 sky130_fd_sc_hd__xnor2_1 _10229_ (.A(_00678_),
    .B(_03313_),
    .Y(_03314_));
 sky130_fd_sc_hd__a22o_1 _10230_ (.A1(net40),
    .A2(_00354_),
    .B1(_00361_),
    .B2(net38),
    .X(_03315_));
 sky130_fd_sc_hd__xor2_1 _10231_ (.A(_00245_),
    .B(_03315_),
    .X(_03316_));
 sky130_fd_sc_hd__nand2b_1 _10232_ (.A_N(_03314_),
    .B(_03316_),
    .Y(_03317_));
 sky130_fd_sc_hd__xor2_1 _10233_ (.A(_03314_),
    .B(_03316_),
    .X(_03318_));
 sky130_fd_sc_hd__a22o_1 _10234_ (.A1(net41),
    .A2(net118),
    .B1(_00366_),
    .B2(net43),
    .X(_03319_));
 sky130_fd_sc_hd__xor2_1 _10235_ (.A(net92),
    .B(_03319_),
    .X(_03320_));
 sky130_fd_sc_hd__nand2b_1 _10236_ (.A_N(_03318_),
    .B(_03320_),
    .Y(_03321_));
 sky130_fd_sc_hd__xnor2_1 _10237_ (.A(_03318_),
    .B(_03320_),
    .Y(_03322_));
 sky130_fd_sc_hd__a21o_1 _10238_ (.A1(_03144_),
    .A2(_03150_),
    .B1(_03149_),
    .X(_03323_));
 sky130_fd_sc_hd__a21o_1 _10239_ (.A1(_00697_),
    .A2(_00698_),
    .B1(net106),
    .X(_03324_));
 sky130_fd_sc_hd__or3_1 _10240_ (.A(net104),
    .B(_00405_),
    .C(_00407_),
    .X(_03325_));
 sky130_fd_sc_hd__a21o_1 _10241_ (.A1(_03324_),
    .A2(_03325_),
    .B1(net136),
    .X(_03326_));
 sky130_fd_sc_hd__nand3_1 _10242_ (.A(net135),
    .B(_03324_),
    .C(_03325_),
    .Y(_03327_));
 sky130_fd_sc_hd__nand3_2 _10243_ (.A(net203),
    .B(_03326_),
    .C(_03327_),
    .Y(_03328_));
 sky130_fd_sc_hd__a21o_1 _10244_ (.A1(_03326_),
    .A2(_03327_),
    .B1(net203),
    .X(_03329_));
 sky130_fd_sc_hd__o22a_1 _10245_ (.A1(net132),
    .A2(net13),
    .B1(net8),
    .B2(net134),
    .X(_03330_));
 sky130_fd_sc_hd__xor2_2 _10246_ (.A(net182),
    .B(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__nand3_2 _10247_ (.A(_03328_),
    .B(_03329_),
    .C(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__a21o_1 _10248_ (.A1(_03328_),
    .A2(_03329_),
    .B1(_03331_),
    .X(_03333_));
 sky130_fd_sc_hd__nand3_2 _10249_ (.A(_03323_),
    .B(_03332_),
    .C(_03333_),
    .Y(_03334_));
 sky130_fd_sc_hd__a21o_1 _10250_ (.A1(_03332_),
    .A2(_03333_),
    .B1(_03323_),
    .X(_03335_));
 sky130_fd_sc_hd__nand3b_1 _10251_ (.A_N(_03181_),
    .B(_03334_),
    .C(_03335_),
    .Y(_03336_));
 sky130_fd_sc_hd__a21bo_1 _10252_ (.A1(_03334_),
    .A2(_03335_),
    .B1_N(_03181_),
    .X(_03337_));
 sky130_fd_sc_hd__and3_1 _10253_ (.A(_03322_),
    .B(_03336_),
    .C(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__a21oi_1 _10254_ (.A1(_03336_),
    .A2(_03337_),
    .B1(_03322_),
    .Y(_03339_));
 sky130_fd_sc_hd__or3_1 _10255_ (.A(_03312_),
    .B(_03338_),
    .C(_03339_),
    .X(_03340_));
 sky130_fd_sc_hd__o21ai_1 _10256_ (.A1(_03338_),
    .A2(_03339_),
    .B1(_03312_),
    .Y(_03341_));
 sky130_fd_sc_hd__and3_1 _10257_ (.A(_03305_),
    .B(_03340_),
    .C(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__a21oi_1 _10258_ (.A1(_03340_),
    .A2(_03341_),
    .B1(_03305_),
    .Y(_03343_));
 sky130_fd_sc_hd__nor2_2 _10259_ (.A(_03342_),
    .B(_03343_),
    .Y(_03344_));
 sky130_fd_sc_hd__xnor2_4 _10260_ (.A(_03289_),
    .B(_03344_),
    .Y(_03345_));
 sky130_fd_sc_hd__a21bo_2 _10261_ (.A1(_03191_),
    .A2(_03206_),
    .B1_N(_03189_),
    .X(_03346_));
 sky130_fd_sc_hd__a21oi_2 _10262_ (.A1(_03209_),
    .A2(_03213_),
    .B1(_03212_),
    .Y(_03347_));
 sky130_fd_sc_hd__a21bo_1 _10263_ (.A1(_03202_),
    .A2(_03203_),
    .B1_N(_03205_),
    .X(_03348_));
 sky130_fd_sc_hd__o21ai_2 _10264_ (.A1(_03142_),
    .A2(_03174_),
    .B1(_03173_),
    .Y(_03349_));
 sky130_fd_sc_hd__nor2_1 _10265_ (.A(_03185_),
    .B(_03187_),
    .Y(_03350_));
 sky130_fd_sc_hd__o21ai_1 _10266_ (.A1(_03185_),
    .A2(_03187_),
    .B1(_03349_),
    .Y(_03351_));
 sky130_fd_sc_hd__xnor2_2 _10267_ (.A(_03349_),
    .B(_03350_),
    .Y(_03352_));
 sky130_fd_sc_hd__xnor2_2 _10268_ (.A(_03348_),
    .B(_03352_),
    .Y(_03353_));
 sky130_fd_sc_hd__nor2_1 _10269_ (.A(_03347_),
    .B(_03353_),
    .Y(_03354_));
 sky130_fd_sc_hd__xnor2_2 _10270_ (.A(_03347_),
    .B(_03353_),
    .Y(_03355_));
 sky130_fd_sc_hd__and2b_1 _10271_ (.A_N(_03355_),
    .B(_03346_),
    .X(_03356_));
 sky130_fd_sc_hd__xnor2_4 _10272_ (.A(_03346_),
    .B(_03355_),
    .Y(_03357_));
 sky130_fd_sc_hd__nand2_1 _10273_ (.A(_03345_),
    .B(_03357_),
    .Y(_03358_));
 sky130_fd_sc_hd__xor2_4 _10274_ (.A(_03345_),
    .B(_03357_),
    .X(_03359_));
 sky130_fd_sc_hd__xnor2_4 _10275_ (.A(_03274_),
    .B(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__xnor2_4 _10276_ (.A(_03273_),
    .B(_03360_),
    .Y(_03361_));
 sky130_fd_sc_hd__nor2_1 _10277_ (.A(_03086_),
    .B(_03222_),
    .Y(_03362_));
 sky130_fd_sc_hd__nand2_1 _10278_ (.A(_03089_),
    .B(_03362_),
    .Y(_03363_));
 sky130_fd_sc_hd__o22a_1 _10279_ (.A1(_02998_),
    .A2(_03085_),
    .B1(_03136_),
    .B2(_03221_),
    .X(_03364_));
 sky130_fd_sc_hd__a21oi_1 _10280_ (.A1(_03136_),
    .A2(_03221_),
    .B1(_03364_),
    .Y(_03365_));
 sky130_fd_sc_hd__a21oi_1 _10281_ (.A1(_03088_),
    .A2(_03362_),
    .B1(_03365_),
    .Y(_03366_));
 sky130_fd_sc_hd__o21ai_4 _10282_ (.A1(_02801_),
    .A2(_03363_),
    .B1(_03366_),
    .Y(_03367_));
 sky130_fd_sc_hd__xnor2_4 _10283_ (.A(_03361_),
    .B(_03367_),
    .Y(_03368_));
 sky130_fd_sc_hd__o21ai_1 _10284_ (.A1(_03272_),
    .A2(_03368_),
    .B1(net200),
    .Y(_03369_));
 sky130_fd_sc_hd__a21oi_1 _10285_ (.A1(_03272_),
    .A2(_03368_),
    .B1(_03369_),
    .Y(_03370_));
 sky130_fd_sc_hd__o21ai_1 _10286_ (.A1(net158),
    .A2(_01816_),
    .B1(_01817_),
    .Y(_03371_));
 sky130_fd_sc_hd__or3_1 _10287_ (.A(net158),
    .B(_01816_),
    .C(_01817_),
    .X(_03372_));
 sky130_fd_sc_hd__a21oi_1 _10288_ (.A1(_06326_),
    .A2(_03239_),
    .B1(_06327_),
    .Y(_03373_));
 sky130_fd_sc_hd__mux2_1 _10289_ (.A0(_06378_),
    .A1(_03373_),
    .S(net285),
    .X(_03374_));
 sky130_fd_sc_hd__or2_1 _10290_ (.A(_06323_),
    .B(_03374_),
    .X(_03375_));
 sky130_fd_sc_hd__nand2_1 _10291_ (.A(_06323_),
    .B(_03374_),
    .Y(_03376_));
 sky130_fd_sc_hd__o21a_1 _10292_ (.A1(net222),
    .A2(_02291_),
    .B1(_02342_),
    .X(_03377_));
 sky130_fd_sc_hd__o21a_1 _10293_ (.A1(net226),
    .A2(_03377_),
    .B1(_02335_),
    .X(_03378_));
 sky130_fd_sc_hd__mux2_1 _10294_ (.A0(_02808_),
    .A1(_02810_),
    .S(net220),
    .X(_03379_));
 sky130_fd_sc_hd__mux2_1 _10295_ (.A0(_02811_),
    .A1(_02816_),
    .S(net219),
    .X(_03380_));
 sky130_fd_sc_hd__mux2_1 _10296_ (.A0(_03379_),
    .A1(_03380_),
    .S(net222),
    .X(_03381_));
 sky130_fd_sc_hd__mux2_1 _10297_ (.A0(_02814_),
    .A1(_02817_),
    .S(_06352_),
    .X(_03382_));
 sky130_fd_sc_hd__mux2_1 _10298_ (.A0(_02340_),
    .A1(_03382_),
    .S(net224),
    .X(_03383_));
 sky130_fd_sc_hd__mux2_1 _10299_ (.A0(_03381_),
    .A1(_03383_),
    .S(net226),
    .X(_03384_));
 sky130_fd_sc_hd__or2_1 _10300_ (.A(\div_res[6] ),
    .B(_03252_),
    .X(_03385_));
 sky130_fd_sc_hd__a21oi_1 _10301_ (.A1(net165),
    .A2(_03385_),
    .B1(\div_res[7] ),
    .Y(_03386_));
 sky130_fd_sc_hd__a31o_1 _10302_ (.A1(\div_res[7] ),
    .A2(net165),
    .A3(_03385_),
    .B1(net195),
    .X(_03387_));
 sky130_fd_sc_hd__or2_1 _10303_ (.A(\div_shifter[38] ),
    .B(_03256_),
    .X(_03388_));
 sky130_fd_sc_hd__a21oi_1 _10304_ (.A1(net235),
    .A2(_03388_),
    .B1(\div_shifter[39] ),
    .Y(_03389_));
 sky130_fd_sc_hd__a31o_1 _10305_ (.A1(\div_shifter[39] ),
    .A2(net235),
    .A3(_03388_),
    .B1(net193),
    .X(_03390_));
 sky130_fd_sc_hd__o2bb2a_1 _10306_ (.A1_N(_06320_),
    .A2_N(net241),
    .B1(_03389_),
    .B2(_03390_),
    .X(_03391_));
 sky130_fd_sc_hd__o221a_1 _10307_ (.A1(_06321_),
    .A2(net199),
    .B1(net196),
    .B2(_06322_),
    .C1(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__o221ai_1 _10308_ (.A1(_06323_),
    .A2(net197),
    .B1(_03386_),
    .B2(_03387_),
    .C1(_03392_),
    .Y(_03393_));
 sky130_fd_sc_hd__o21a_1 _10309_ (.A1(_03261_),
    .A2(_03262_),
    .B1(_03263_),
    .X(_03394_));
 sky130_fd_sc_hd__nor2_1 _10310_ (.A(reg1_val[7]),
    .B(curr_PC[7]),
    .Y(_03395_));
 sky130_fd_sc_hd__nand2_1 _10311_ (.A(reg1_val[7]),
    .B(curr_PC[7]),
    .Y(_03396_));
 sky130_fd_sc_hd__and2b_1 _10312_ (.A_N(_03395_),
    .B(_03396_),
    .X(_03397_));
 sky130_fd_sc_hd__xnor2_1 _10313_ (.A(_03394_),
    .B(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__a31o_1 _10314_ (.A1(net249),
    .A2(net210),
    .A3(_03398_),
    .B1(_03393_),
    .X(_03399_));
 sky130_fd_sc_hd__a221o_1 _10315_ (.A1(net179),
    .A2(_03378_),
    .B1(_03384_),
    .B2(_02975_),
    .C1(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__a31o_1 _10316_ (.A1(_02317_),
    .A2(_03375_),
    .A3(_03376_),
    .B1(_03400_),
    .X(_03401_));
 sky130_fd_sc_hd__a311o_1 _10317_ (.A1(_02323_),
    .A2(_03371_),
    .A3(_03372_),
    .B1(_03401_),
    .C1(_03370_),
    .X(_03402_));
 sky130_fd_sc_hd__or2_1 _10318_ (.A(curr_PC[7]),
    .B(_03270_),
    .X(_03403_));
 sky130_fd_sc_hd__a21oi_1 _10319_ (.A1(curr_PC[7]),
    .A2(_03270_),
    .B1(net242),
    .Y(_03404_));
 sky130_fd_sc_hd__a22o_4 _10320_ (.A1(net242),
    .A2(_03402_),
    .B1(_03403_),
    .B2(_03404_),
    .X(dest_val[7]));
 sky130_fd_sc_hd__nor3_1 _10321_ (.A(_02132_),
    .B(_02239_),
    .C(_02644_),
    .Y(_03405_));
 sky130_fd_sc_hd__o21ba_1 _10322_ (.A1(_02955_),
    .A2(_02956_),
    .B1_N(_02467_),
    .X(_03406_));
 sky130_fd_sc_hd__a21boi_1 _10323_ (.A1(_03230_),
    .A2(_03231_),
    .B1_N(_02802_),
    .Y(_03407_));
 sky130_fd_sc_hd__nand4_2 _10324_ (.A(_03093_),
    .B(_03405_),
    .C(_03406_),
    .D(_03407_),
    .Y(_03408_));
 sky130_fd_sc_hd__nor2_1 _10325_ (.A(_03368_),
    .B(_03408_),
    .Y(_03409_));
 sky130_fd_sc_hd__or2_1 _10326_ (.A(net158),
    .B(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__o22a_1 _10327_ (.A1(_03136_),
    .A2(_03221_),
    .B1(_03273_),
    .B2(_03360_),
    .X(_03411_));
 sky130_fd_sc_hd__a21oi_1 _10328_ (.A1(_03273_),
    .A2(_03360_),
    .B1(_03411_),
    .Y(_03412_));
 sky130_fd_sc_hd__nor2_1 _10329_ (.A(_03222_),
    .B(_03361_),
    .Y(_03413_));
 sky130_fd_sc_hd__a21oi_2 _10330_ (.A1(_03227_),
    .A2(_03413_),
    .B1(_03412_),
    .Y(_03414_));
 sky130_fd_sc_hd__or4_2 _10331_ (.A(_02950_),
    .B(_03086_),
    .C(_03222_),
    .D(_03361_),
    .X(_03415_));
 sky130_fd_sc_hd__a211o_1 _10332_ (.A1(_02133_),
    .A2(_02135_),
    .B1(_02951_),
    .C1(_03415_),
    .X(_03416_));
 sky130_fd_sc_hd__o211ai_4 _10333_ (.A1(_02954_),
    .A2(_03415_),
    .B1(_03416_),
    .C1(_03414_),
    .Y(_03417_));
 sky130_fd_sc_hd__a21boi_4 _10334_ (.A1(_03274_),
    .A2(_03359_),
    .B1_N(_03358_),
    .Y(_03418_));
 sky130_fd_sc_hd__o22a_1 _10335_ (.A1(net112),
    .A2(net11),
    .B1(net6),
    .B2(net110),
    .X(_03419_));
 sky130_fd_sc_hd__xnor2_1 _10336_ (.A(net19),
    .B(_03419_),
    .Y(_03420_));
 sky130_fd_sc_hd__nand2_1 _10337_ (.A(_00308_),
    .B(_02078_),
    .Y(_03421_));
 sky130_fd_sc_hd__o22a_1 _10338_ (.A1(net119),
    .A2(net23),
    .B1(net15),
    .B2(net117),
    .X(_03422_));
 sky130_fd_sc_hd__xnor2_1 _10339_ (.A(net70),
    .B(_03422_),
    .Y(_03423_));
 sky130_fd_sc_hd__or2_1 _10340_ (.A(_03421_),
    .B(_03423_),
    .X(_03424_));
 sky130_fd_sc_hd__xnor2_1 _10341_ (.A(_03421_),
    .B(_03423_),
    .Y(_03425_));
 sky130_fd_sc_hd__or2_1 _10342_ (.A(_03420_),
    .B(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__nand2_1 _10343_ (.A(_03420_),
    .B(_03425_),
    .Y(_03427_));
 sky130_fd_sc_hd__and2_1 _10344_ (.A(_03426_),
    .B(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__o21bai_1 _10345_ (.A1(_03297_),
    .A2(_03299_),
    .B1_N(_03295_),
    .Y(_03429_));
 sky130_fd_sc_hd__a21bo_1 _10346_ (.A1(_03329_),
    .A2(_03331_),
    .B1_N(_03328_),
    .X(_03430_));
 sky130_fd_sc_hd__o22a_1 _10347_ (.A1(_00391_),
    .A2(net14),
    .B1(net13),
    .B2(net106),
    .X(_03431_));
 sky130_fd_sc_hd__xnor2_2 _10348_ (.A(_00342_),
    .B(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__o21ba_1 _10349_ (.A1(_00183_),
    .A2(net8),
    .B1_N(net181),
    .X(_03433_));
 sky130_fd_sc_hd__nor2_1 _10350_ (.A(_00182_),
    .B(net8),
    .Y(_03434_));
 sky130_fd_sc_hd__a21o_1 _10351_ (.A1(net181),
    .A2(_03434_),
    .B1(_03433_),
    .X(_03435_));
 sky130_fd_sc_hd__nor2_1 _10352_ (.A(_03432_),
    .B(_03435_),
    .Y(_03436_));
 sky130_fd_sc_hd__xor2_2 _10353_ (.A(_03432_),
    .B(_03435_),
    .X(_03437_));
 sky130_fd_sc_hd__a21oi_1 _10354_ (.A1(_03328_),
    .A2(_03332_),
    .B1(_03437_),
    .Y(_03438_));
 sky130_fd_sc_hd__xnor2_2 _10355_ (.A(_03430_),
    .B(_03437_),
    .Y(_03439_));
 sky130_fd_sc_hd__xor2_1 _10356_ (.A(_03429_),
    .B(_03439_),
    .X(_03440_));
 sky130_fd_sc_hd__o22a_1 _10357_ (.A1(net101),
    .A2(net47),
    .B1(net45),
    .B2(net99),
    .X(_03441_));
 sky130_fd_sc_hd__xnor2_1 _10358_ (.A(net96),
    .B(_03441_),
    .Y(_03442_));
 sky130_fd_sc_hd__a22o_1 _10359_ (.A1(net43),
    .A2(_00361_),
    .B1(_00366_),
    .B2(net41),
    .X(_03443_));
 sky130_fd_sc_hd__xor2_1 _10360_ (.A(net92),
    .B(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__and2_1 _10361_ (.A(_03442_),
    .B(_03444_),
    .X(_03445_));
 sky130_fd_sc_hd__nor2_1 _10362_ (.A(_03442_),
    .B(_03444_),
    .Y(_03446_));
 sky130_fd_sc_hd__nor2_1 _10363_ (.A(_03445_),
    .B(_03446_),
    .Y(_03447_));
 sky130_fd_sc_hd__a22o_1 _10364_ (.A1(net40),
    .A2(_00348_),
    .B1(_00354_),
    .B2(net38),
    .X(_03448_));
 sky130_fd_sc_hd__xor2_1 _10365_ (.A(_00245_),
    .B(_03448_),
    .X(_03449_));
 sky130_fd_sc_hd__xor2_1 _10366_ (.A(_03447_),
    .B(_03449_),
    .X(_03450_));
 sky130_fd_sc_hd__xor2_1 _10367_ (.A(_03440_),
    .B(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__xnor2_1 _10368_ (.A(_03428_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__a21o_1 _10369_ (.A1(_03283_),
    .A2(_03285_),
    .B1(_03281_),
    .X(_03453_));
 sky130_fd_sc_hd__o32a_1 _10370_ (.A1(_00347_),
    .A2(_00405_),
    .A3(_00407_),
    .B1(net83),
    .B2(net55),
    .X(_03454_));
 sky130_fd_sc_hd__xnor2_2 _10371_ (.A(_00339_),
    .B(_03454_),
    .Y(_03455_));
 sky130_fd_sc_hd__o22a_1 _10372_ (.A1(net67),
    .A2(net79),
    .B1(net74),
    .B2(net65),
    .X(_03456_));
 sky130_fd_sc_hd__xor2_2 _10373_ (.A(net122),
    .B(_03456_),
    .X(_03457_));
 sky130_fd_sc_hd__xnor2_1 _10374_ (.A(_03455_),
    .B(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__a21oi_1 _10375_ (.A1(_03317_),
    .A2(_03321_),
    .B1(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__and3_1 _10376_ (.A(_03317_),
    .B(_03321_),
    .C(_03458_),
    .X(_03460_));
 sky130_fd_sc_hd__or2_1 _10377_ (.A(_03459_),
    .B(_03460_),
    .X(_03461_));
 sky130_fd_sc_hd__and2b_1 _10378_ (.A_N(_03461_),
    .B(_03453_),
    .X(_03462_));
 sky130_fd_sc_hd__xor2_1 _10379_ (.A(_03453_),
    .B(_03461_),
    .X(_03463_));
 sky130_fd_sc_hd__nor2_1 _10380_ (.A(_03452_),
    .B(_03463_),
    .Y(_03464_));
 sky130_fd_sc_hd__nand2_1 _10381_ (.A(_03452_),
    .B(_03463_),
    .Y(_03465_));
 sky130_fd_sc_hd__and2b_1 _10382_ (.A_N(_03464_),
    .B(_03465_),
    .X(_03466_));
 sky130_fd_sc_hd__nand2_1 _10383_ (.A(_03334_),
    .B(_03336_),
    .Y(_03467_));
 sky130_fd_sc_hd__o22a_1 _10384_ (.A1(net59),
    .A2(net36),
    .B1(net34),
    .B2(net57),
    .X(_03468_));
 sky130_fd_sc_hd__xnor2_1 _10385_ (.A(net126),
    .B(_03468_),
    .Y(_03469_));
 sky130_fd_sc_hd__a22o_1 _10386_ (.A1(_00163_),
    .A2(net32),
    .B1(net30),
    .B2(_00172_),
    .X(_03470_));
 sky130_fd_sc_hd__xnor2_1 _10387_ (.A(net50),
    .B(_03470_),
    .Y(_03471_));
 sky130_fd_sc_hd__and2_1 _10388_ (.A(_03469_),
    .B(_03471_),
    .X(_03472_));
 sky130_fd_sc_hd__nor2_1 _10389_ (.A(_03469_),
    .B(_03471_),
    .Y(_03473_));
 sky130_fd_sc_hd__nor2_1 _10390_ (.A(_03472_),
    .B(_03473_),
    .Y(_03474_));
 sky130_fd_sc_hd__o22a_1 _10391_ (.A1(net64),
    .A2(net28),
    .B1(net26),
    .B2(net62),
    .X(_03475_));
 sky130_fd_sc_hd__xnor2_1 _10392_ (.A(_00301_),
    .B(_03475_),
    .Y(_03476_));
 sky130_fd_sc_hd__xor2_1 _10393_ (.A(_03474_),
    .B(_03476_),
    .X(_03477_));
 sky130_fd_sc_hd__o21a_1 _10394_ (.A1(_03308_),
    .A2(_03310_),
    .B1(_03477_),
    .X(_03478_));
 sky130_fd_sc_hd__or3_1 _10395_ (.A(_03308_),
    .B(_03310_),
    .C(_03477_),
    .X(_03479_));
 sky130_fd_sc_hd__and2b_1 _10396_ (.A_N(_03478_),
    .B(_03479_),
    .X(_03480_));
 sky130_fd_sc_hd__xor2_1 _10397_ (.A(_03467_),
    .B(_03480_),
    .X(_03481_));
 sky130_fd_sc_hd__xnor2_1 _10398_ (.A(_03466_),
    .B(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__o21bai_1 _10399_ (.A1(_03289_),
    .A2(_03343_),
    .B1_N(_03342_),
    .Y(_03483_));
 sky130_fd_sc_hd__a21o_1 _10400_ (.A1(_03275_),
    .A2(_03288_),
    .B1(_03287_),
    .X(_03484_));
 sky130_fd_sc_hd__or2_1 _10401_ (.A(_03302_),
    .B(_03304_),
    .X(_03485_));
 sky130_fd_sc_hd__o21ba_1 _10402_ (.A1(_03312_),
    .A2(_03339_),
    .B1_N(_03338_),
    .X(_03486_));
 sky130_fd_sc_hd__o21ba_1 _10403_ (.A1(_03302_),
    .A2(_03304_),
    .B1_N(_03486_),
    .X(_03487_));
 sky130_fd_sc_hd__xnor2_1 _10404_ (.A(_03485_),
    .B(_03486_),
    .Y(_03488_));
 sky130_fd_sc_hd__xnor2_1 _10405_ (.A(_03484_),
    .B(_03488_),
    .Y(_03489_));
 sky130_fd_sc_hd__a21boi_1 _10406_ (.A1(_03348_),
    .A2(_03352_),
    .B1_N(_03351_),
    .Y(_03490_));
 sky130_fd_sc_hd__nor2_1 _10407_ (.A(_03489_),
    .B(_03490_),
    .Y(_03491_));
 sky130_fd_sc_hd__xor2_1 _10408_ (.A(_03489_),
    .B(_03490_),
    .X(_03492_));
 sky130_fd_sc_hd__xnor2_1 _10409_ (.A(_03483_),
    .B(_03492_),
    .Y(_03493_));
 sky130_fd_sc_hd__nor2_1 _10410_ (.A(_03482_),
    .B(_03493_),
    .Y(_03494_));
 sky130_fd_sc_hd__xor2_1 _10411_ (.A(_03482_),
    .B(_03493_),
    .X(_03495_));
 sky130_fd_sc_hd__o21a_1 _10412_ (.A1(_03354_),
    .A2(_03356_),
    .B1(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__nor3_1 _10413_ (.A(_03354_),
    .B(_03356_),
    .C(_03495_),
    .Y(_03497_));
 sky130_fd_sc_hd__or2_4 _10414_ (.A(_03496_),
    .B(_03497_),
    .X(_03498_));
 sky130_fd_sc_hd__xnor2_4 _10415_ (.A(_03418_),
    .B(_03498_),
    .Y(_03499_));
 sky130_fd_sc_hd__xor2_4 _10416_ (.A(_03417_),
    .B(_03499_),
    .X(_03500_));
 sky130_fd_sc_hd__o21ai_1 _10417_ (.A1(_03410_),
    .A2(_03500_),
    .B1(net200),
    .Y(_03501_));
 sky130_fd_sc_hd__a21o_1 _10418_ (.A1(_03410_),
    .A2(_03500_),
    .B1(_03501_),
    .X(_03502_));
 sky130_fd_sc_hd__o21a_1 _10419_ (.A1(net157),
    .A2(_01818_),
    .B1(_01819_),
    .X(_03503_));
 sky130_fd_sc_hd__nor3_1 _10420_ (.A(net157),
    .B(_01818_),
    .C(_01819_),
    .Y(_03504_));
 sky130_fd_sc_hd__o21a_1 _10421_ (.A1(_06321_),
    .A2(_03373_),
    .B1(_06322_),
    .X(_03505_));
 sky130_fd_sc_hd__mux2_1 _10422_ (.A0(_06380_),
    .A1(_03505_),
    .S(net285),
    .X(_03506_));
 sky130_fd_sc_hd__nor2_1 _10423_ (.A(_06318_),
    .B(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__a211o_1 _10424_ (.A1(_06318_),
    .A2(_03506_),
    .B1(_03507_),
    .C1(net236),
    .X(_03508_));
 sky130_fd_sc_hd__o21a_1 _10425_ (.A1(_03394_),
    .A2(_03395_),
    .B1(_03396_),
    .X(_03509_));
 sky130_fd_sc_hd__nor2_1 _10426_ (.A(reg1_val[8]),
    .B(curr_PC[8]),
    .Y(_03510_));
 sky130_fd_sc_hd__nand2_1 _10427_ (.A(reg1_val[8]),
    .B(curr_PC[8]),
    .Y(_03511_));
 sky130_fd_sc_hd__nand2b_1 _10428_ (.A_N(_03510_),
    .B(_03511_),
    .Y(_03512_));
 sky130_fd_sc_hd__xnor2_1 _10429_ (.A(_03509_),
    .B(_03512_),
    .Y(_03513_));
 sky130_fd_sc_hd__mux2_1 _10430_ (.A0(_02275_),
    .A1(_02306_),
    .S(net222),
    .X(_03514_));
 sky130_fd_sc_hd__or2_1 _10431_ (.A(net226),
    .B(_03514_),
    .X(_03515_));
 sky130_fd_sc_hd__o21ai_2 _10432_ (.A1(net225),
    .A2(_03377_),
    .B1(_03515_),
    .Y(_03516_));
 sky130_fd_sc_hd__mux2_1 _10433_ (.A0(_03513_),
    .A1(_03516_),
    .S(net229),
    .X(_03517_));
 sky130_fd_sc_hd__or2_1 _10434_ (.A(\div_res[7] ),
    .B(_03385_),
    .X(_03518_));
 sky130_fd_sc_hd__a21oi_1 _10435_ (.A1(net165),
    .A2(_03518_),
    .B1(\div_res[8] ),
    .Y(_03519_));
 sky130_fd_sc_hd__a31o_1 _10436_ (.A1(\div_res[8] ),
    .A2(net165),
    .A3(_03518_),
    .B1(net195),
    .X(_03520_));
 sky130_fd_sc_hd__a21oi_1 _10437_ (.A1(_06317_),
    .A2(_02319_),
    .B1(_02315_),
    .Y(_03521_));
 sky130_fd_sc_hd__or2_1 _10438_ (.A(\div_shifter[39] ),
    .B(_03388_),
    .X(_03522_));
 sky130_fd_sc_hd__a21oi_1 _10439_ (.A1(net235),
    .A2(_03522_),
    .B1(\div_shifter[40] ),
    .Y(_03523_));
 sky130_fd_sc_hd__a31o_1 _10440_ (.A1(\div_shifter[40] ),
    .A2(net235),
    .A3(_03522_),
    .B1(net193),
    .X(_03524_));
 sky130_fd_sc_hd__o2bb2a_1 _10441_ (.A1_N(_06315_),
    .A2_N(_06487_),
    .B1(_03523_),
    .B2(_03524_),
    .X(_03525_));
 sky130_fd_sc_hd__o221a_1 _10442_ (.A1(_06317_),
    .A2(net196),
    .B1(_03521_),
    .B2(_06316_),
    .C1(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__o21a_1 _10443_ (.A1(_03519_),
    .A2(_03520_),
    .B1(_03526_),
    .X(_03527_));
 sky130_fd_sc_hd__o21ai_2 _10444_ (.A1(net226),
    .A2(_03383_),
    .B1(_02335_),
    .Y(_03528_));
 sky130_fd_sc_hd__o221a_1 _10445_ (.A1(_02314_),
    .A2(_03516_),
    .B1(_03528_),
    .B2(net177),
    .C1(_03527_),
    .X(_03529_));
 sky130_fd_sc_hd__o211a_1 _10446_ (.A1(_06476_),
    .A2(_03517_),
    .B1(_03529_),
    .C1(_03508_),
    .X(_03530_));
 sky130_fd_sc_hd__o311a_1 _10447_ (.A1(_02324_),
    .A2(_03503_),
    .A3(_03504_),
    .B1(_03530_),
    .C1(_03502_),
    .X(_03531_));
 sky130_fd_sc_hd__and3_1 _10448_ (.A(curr_PC[7]),
    .B(curr_PC[8]),
    .C(_03270_),
    .X(_03532_));
 sky130_fd_sc_hd__a21oi_1 _10449_ (.A1(curr_PC[7]),
    .A2(_03270_),
    .B1(curr_PC[8]),
    .Y(_03533_));
 sky130_fd_sc_hd__or3_1 _10450_ (.A(net242),
    .B(_03532_),
    .C(_03533_),
    .X(_03534_));
 sky130_fd_sc_hd__o21ai_4 _10451_ (.A1(net248),
    .A2(_03531_),
    .B1(_03534_),
    .Y(dest_val[8]));
 sky130_fd_sc_hd__xor2_1 _10452_ (.A(curr_PC[9]),
    .B(_03532_),
    .X(_03535_));
 sky130_fd_sc_hd__nand2_1 _10453_ (.A(_03409_),
    .B(_03500_),
    .Y(_03536_));
 sky130_fd_sc_hd__a21o_1 _10454_ (.A1(_03483_),
    .A2(_03492_),
    .B1(_03491_),
    .X(_03537_));
 sky130_fd_sc_hd__a21o_1 _10455_ (.A1(_03429_),
    .A2(_03439_),
    .B1(_03438_),
    .X(_03538_));
 sky130_fd_sc_hd__o22a_1 _10456_ (.A1(net55),
    .A2(net79),
    .B1(net74),
    .B2(net67),
    .X(_03539_));
 sky130_fd_sc_hd__xnor2_1 _10457_ (.A(net122),
    .B(_03539_),
    .Y(_03540_));
 sky130_fd_sc_hd__o22a_1 _10458_ (.A1(net58),
    .A2(net28),
    .B1(net26),
    .B2(net64),
    .X(_03541_));
 sky130_fd_sc_hd__xnor2_1 _10459_ (.A(_00301_),
    .B(_03541_),
    .Y(_03542_));
 sky130_fd_sc_hd__nand2b_1 _10460_ (.A_N(_03540_),
    .B(_03542_),
    .Y(_03543_));
 sky130_fd_sc_hd__xor2_1 _10461_ (.A(_03540_),
    .B(_03542_),
    .X(_03544_));
 sky130_fd_sc_hd__o22a_1 _10462_ (.A1(net65),
    .A2(net36),
    .B1(net34),
    .B2(net60),
    .X(_03545_));
 sky130_fd_sc_hd__xnor2_1 _10463_ (.A(net126),
    .B(_03545_),
    .Y(_03546_));
 sky130_fd_sc_hd__nand2b_1 _10464_ (.A_N(_03544_),
    .B(_03546_),
    .Y(_03547_));
 sky130_fd_sc_hd__nand2b_1 _10465_ (.A_N(_03546_),
    .B(_03544_),
    .Y(_03548_));
 sky130_fd_sc_hd__nand2_1 _10466_ (.A(_03547_),
    .B(_03548_),
    .Y(_03549_));
 sky130_fd_sc_hd__a21oi_1 _10467_ (.A1(_03424_),
    .A2(_03426_),
    .B1(_03549_),
    .Y(_03550_));
 sky130_fd_sc_hd__and3_1 _10468_ (.A(_03424_),
    .B(_03426_),
    .C(_03549_),
    .X(_03551_));
 sky130_fd_sc_hd__or2_1 _10469_ (.A(_03550_),
    .B(_03551_),
    .X(_03552_));
 sky130_fd_sc_hd__and2b_1 _10470_ (.A_N(_03552_),
    .B(_03538_),
    .X(_03553_));
 sky130_fd_sc_hd__xnor2_1 _10471_ (.A(_03538_),
    .B(_03552_),
    .Y(_03554_));
 sky130_fd_sc_hd__a21oi_1 _10472_ (.A1(_03474_),
    .A2(_03476_),
    .B1(_03472_),
    .Y(_03555_));
 sky130_fd_sc_hd__o22a_1 _10473_ (.A1(net104),
    .A2(net12),
    .B1(net7),
    .B2(net106),
    .X(_03556_));
 sky130_fd_sc_hd__xnor2_2 _10474_ (.A(_00342_),
    .B(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__a21o_1 _10475_ (.A1(_00697_),
    .A2(_00698_),
    .B1(net87),
    .X(_03558_));
 sky130_fd_sc_hd__or3_1 _10476_ (.A(net83),
    .B(_00405_),
    .C(_00407_),
    .X(_03559_));
 sky130_fd_sc_hd__a21o_1 _10477_ (.A1(_03558_),
    .A2(_03559_),
    .B1(net138),
    .X(_03560_));
 sky130_fd_sc_hd__nand3_1 _10478_ (.A(net137),
    .B(_03558_),
    .C(_03559_),
    .Y(_03561_));
 sky130_fd_sc_hd__nand3_1 _10479_ (.A(net181),
    .B(_03560_),
    .C(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__a21o_1 _10480_ (.A1(_03560_),
    .A2(_03561_),
    .B1(net181),
    .X(_03563_));
 sky130_fd_sc_hd__nand2_1 _10481_ (.A(_03562_),
    .B(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__xnor2_2 _10482_ (.A(_03557_),
    .B(_03564_),
    .Y(_03565_));
 sky130_fd_sc_hd__a21o_1 _10483_ (.A1(_03447_),
    .A2(_03449_),
    .B1(_03445_),
    .X(_03566_));
 sky130_fd_sc_hd__nand2_1 _10484_ (.A(_03565_),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__xnor2_1 _10485_ (.A(_03565_),
    .B(_03566_),
    .Y(_03568_));
 sky130_fd_sc_hd__nor2_1 _10486_ (.A(_03555_),
    .B(_03568_),
    .Y(_03569_));
 sky130_fd_sc_hd__and2_1 _10487_ (.A(_03555_),
    .B(_03568_),
    .X(_03570_));
 sky130_fd_sc_hd__o22a_1 _10488_ (.A1(net73),
    .A2(net23),
    .B1(net15),
    .B2(net119),
    .X(_03571_));
 sky130_fd_sc_hd__xnor2_1 _10489_ (.A(net70),
    .B(_03571_),
    .Y(_03572_));
 sky130_fd_sc_hd__o22a_1 _10490_ (.A1(_00290_),
    .A2(net11),
    .B1(net6),
    .B2(net112),
    .X(_03573_));
 sky130_fd_sc_hd__xnor2_1 _10491_ (.A(net19),
    .B(_03573_),
    .Y(_03574_));
 sky130_fd_sc_hd__a22o_1 _10492_ (.A1(net43),
    .A2(_00354_),
    .B1(_00361_),
    .B2(net41),
    .X(_03575_));
 sky130_fd_sc_hd__xor2_1 _10493_ (.A(net92),
    .B(_03575_),
    .X(_03576_));
 sky130_fd_sc_hd__nand2b_1 _10494_ (.A_N(_03574_),
    .B(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__nand2b_1 _10495_ (.A_N(_03576_),
    .B(_03574_),
    .Y(_03578_));
 sky130_fd_sc_hd__nand2_1 _10496_ (.A(_03577_),
    .B(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__or2_1 _10497_ (.A(_03572_),
    .B(_03579_),
    .X(_03580_));
 sky130_fd_sc_hd__nand2_1 _10498_ (.A(_03572_),
    .B(_03579_),
    .Y(_03581_));
 sky130_fd_sc_hd__and2_1 _10499_ (.A(_03580_),
    .B(_03581_),
    .X(_03582_));
 sky130_fd_sc_hd__nor2_1 _10500_ (.A(net110),
    .B(net19),
    .Y(_03583_));
 sky130_fd_sc_hd__and3_1 _10501_ (.A(_03455_),
    .B(_03457_),
    .C(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__a21oi_1 _10502_ (.A1(_03455_),
    .A2(_03457_),
    .B1(_03583_),
    .Y(_03585_));
 sky130_fd_sc_hd__or2_1 _10503_ (.A(_03584_),
    .B(_03585_),
    .X(_03586_));
 sky130_fd_sc_hd__xor2_2 _10504_ (.A(_03436_),
    .B(_03586_),
    .X(_03587_));
 sky130_fd_sc_hd__a22o_1 _10505_ (.A1(_00189_),
    .A2(net40),
    .B1(net37),
    .B2(_00348_),
    .X(_03588_));
 sky130_fd_sc_hd__xor2_1 _10506_ (.A(_00245_),
    .B(_03588_),
    .X(_03589_));
 sky130_fd_sc_hd__a22o_1 _10507_ (.A1(_06547_),
    .A2(net32),
    .B1(net30),
    .B2(_00163_),
    .X(_03590_));
 sky130_fd_sc_hd__xnor2_1 _10508_ (.A(net50),
    .B(_03590_),
    .Y(_03591_));
 sky130_fd_sc_hd__and2_1 _10509_ (.A(_03589_),
    .B(_03591_),
    .X(_03592_));
 sky130_fd_sc_hd__nor2_1 _10510_ (.A(_03589_),
    .B(_03591_),
    .Y(_03593_));
 sky130_fd_sc_hd__nor2_1 _10511_ (.A(_03592_),
    .B(_03593_),
    .Y(_03594_));
 sky130_fd_sc_hd__o22a_1 _10512_ (.A1(net52),
    .A2(net47),
    .B1(net45),
    .B2(net101),
    .X(_03595_));
 sky130_fd_sc_hd__xnor2_1 _10513_ (.A(net95),
    .B(_03595_),
    .Y(_03596_));
 sky130_fd_sc_hd__xor2_1 _10514_ (.A(_03594_),
    .B(_03596_),
    .X(_03597_));
 sky130_fd_sc_hd__xor2_1 _10515_ (.A(_03587_),
    .B(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__xnor2_1 _10516_ (.A(_03582_),
    .B(_03598_),
    .Y(_03599_));
 sky130_fd_sc_hd__or3_1 _10517_ (.A(_03569_),
    .B(_03570_),
    .C(_03599_),
    .X(_03600_));
 sky130_fd_sc_hd__o21ai_1 _10518_ (.A1(_03569_),
    .A2(_03570_),
    .B1(_03599_),
    .Y(_03601_));
 sky130_fd_sc_hd__and3_1 _10519_ (.A(_03554_),
    .B(_03600_),
    .C(_03601_),
    .X(_03602_));
 sky130_fd_sc_hd__a21oi_1 _10520_ (.A1(_03600_),
    .A2(_03601_),
    .B1(_03554_),
    .Y(_03603_));
 sky130_fd_sc_hd__nor2_1 _10521_ (.A(_03602_),
    .B(_03603_),
    .Y(_03604_));
 sky130_fd_sc_hd__a21o_1 _10522_ (.A1(_03465_),
    .A2(_03481_),
    .B1(_03464_),
    .X(_03605_));
 sky130_fd_sc_hd__a21o_1 _10523_ (.A1(_03467_),
    .A2(_03479_),
    .B1(_03478_),
    .X(_03606_));
 sky130_fd_sc_hd__a32o_1 _10524_ (.A1(_03426_),
    .A2(_03427_),
    .A3(_03451_),
    .B1(_03450_),
    .B2(_03440_),
    .X(_03607_));
 sky130_fd_sc_hd__nor2_1 _10525_ (.A(_03459_),
    .B(_03462_),
    .Y(_03608_));
 sky130_fd_sc_hd__o21a_1 _10526_ (.A1(_03459_),
    .A2(_03462_),
    .B1(_03607_),
    .X(_03609_));
 sky130_fd_sc_hd__xnor2_1 _10527_ (.A(_03607_),
    .B(_03608_),
    .Y(_03610_));
 sky130_fd_sc_hd__xnor2_1 _10528_ (.A(_03606_),
    .B(_03610_),
    .Y(_03611_));
 sky130_fd_sc_hd__a21oi_1 _10529_ (.A1(_03484_),
    .A2(_03488_),
    .B1(_03487_),
    .Y(_03612_));
 sky130_fd_sc_hd__xnor2_1 _10530_ (.A(_03611_),
    .B(_03612_),
    .Y(_03613_));
 sky130_fd_sc_hd__nand2b_1 _10531_ (.A_N(_03613_),
    .B(_03605_),
    .Y(_03614_));
 sky130_fd_sc_hd__xnor2_2 _10532_ (.A(_03605_),
    .B(_03613_),
    .Y(_03615_));
 sky130_fd_sc_hd__nand2_1 _10533_ (.A(_03604_),
    .B(_03615_),
    .Y(_03616_));
 sky130_fd_sc_hd__xnor2_2 _10534_ (.A(_03604_),
    .B(_03615_),
    .Y(_03617_));
 sky130_fd_sc_hd__nand2b_1 _10535_ (.A_N(_03617_),
    .B(_03537_),
    .Y(_03618_));
 sky130_fd_sc_hd__xnor2_2 _10536_ (.A(_03537_),
    .B(_03617_),
    .Y(_03619_));
 sky130_fd_sc_hd__o21ai_4 _10537_ (.A1(_03494_),
    .A2(_03496_),
    .B1(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__or3_2 _10538_ (.A(_03494_),
    .B(_03496_),
    .C(_03619_),
    .X(_03621_));
 sky130_fd_sc_hd__nand2_4 _10539_ (.A(_03620_),
    .B(_03621_),
    .Y(_03622_));
 sky130_fd_sc_hd__nor2_1 _10540_ (.A(_03361_),
    .B(_03499_),
    .Y(_03623_));
 sky130_fd_sc_hd__and2_1 _10541_ (.A(_03362_),
    .B(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__or4_2 _10542_ (.A(_03086_),
    .B(_03222_),
    .C(_03361_),
    .D(_03499_),
    .X(_03625_));
 sky130_fd_sc_hd__a21oi_2 _10543_ (.A1(_02463_),
    .A2(_02465_),
    .B1(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__o22a_1 _10544_ (.A1(_03273_),
    .A2(_03360_),
    .B1(_03418_),
    .B2(_03498_),
    .X(_03627_));
 sky130_fd_sc_hd__a21oi_2 _10545_ (.A1(_03418_),
    .A2(_03498_),
    .B1(_03627_),
    .Y(_03628_));
 sky130_fd_sc_hd__a21o_2 _10546_ (.A1(_03365_),
    .A2(_03623_),
    .B1(_03628_),
    .X(_03629_));
 sky130_fd_sc_hd__a221oi_4 _10547_ (.A1(_03090_),
    .A2(_03624_),
    .B1(_03626_),
    .B2(net4),
    .C1(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__xor2_4 _10548_ (.A(_03622_),
    .B(_03630_),
    .X(_03631_));
 sky130_fd_sc_hd__nand3_1 _10549_ (.A(net161),
    .B(_03536_),
    .C(_03631_),
    .Y(_03632_));
 sky130_fd_sc_hd__a21o_1 _10550_ (.A1(net162),
    .A2(_03536_),
    .B1(_03631_),
    .X(_03633_));
 sky130_fd_sc_hd__o21ai_1 _10551_ (.A1(net157),
    .A2(_01820_),
    .B1(_01822_),
    .Y(_03634_));
 sky130_fd_sc_hd__or3_1 _10552_ (.A(net157),
    .B(_01820_),
    .C(_01822_),
    .X(_03635_));
 sky130_fd_sc_hd__o21a_1 _10553_ (.A1(_06316_),
    .A2(_03505_),
    .B1(_06317_),
    .X(_03636_));
 sky130_fd_sc_hd__mux2_1 _10554_ (.A0(_06382_),
    .A1(_03636_),
    .S(net285),
    .X(_03637_));
 sky130_fd_sc_hd__a21oi_1 _10555_ (.A1(_06313_),
    .A2(_03637_),
    .B1(net236),
    .Y(_03638_));
 sky130_fd_sc_hd__o21a_1 _10556_ (.A1(_06313_),
    .A2(_03637_),
    .B1(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__o21a_1 _10557_ (.A1(_03509_),
    .A2(_03510_),
    .B1(_03511_),
    .X(_03640_));
 sky130_fd_sc_hd__nor2_1 _10558_ (.A(reg1_val[9]),
    .B(curr_PC[9]),
    .Y(_03641_));
 sky130_fd_sc_hd__nand2_1 _10559_ (.A(reg1_val[9]),
    .B(curr_PC[9]),
    .Y(_03642_));
 sky130_fd_sc_hd__nand2b_1 _10560_ (.A_N(_03641_),
    .B(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__xor2_1 _10561_ (.A(_03640_),
    .B(_03643_),
    .X(_03644_));
 sky130_fd_sc_hd__mux2_1 _10562_ (.A0(_02483_),
    .A1(_02497_),
    .S(net223),
    .X(_03645_));
 sky130_fd_sc_hd__mux2_1 _10563_ (.A0(_03243_),
    .A1(_03645_),
    .S(net225),
    .X(_03646_));
 sky130_fd_sc_hd__mux2_1 _10564_ (.A0(_03644_),
    .A1(_03646_),
    .S(net229),
    .X(_03647_));
 sky130_fd_sc_hd__or2_1 _10565_ (.A(\div_res[8] ),
    .B(_03518_),
    .X(_03648_));
 sky130_fd_sc_hd__a21oi_1 _10566_ (.A1(net165),
    .A2(_03648_),
    .B1(\div_res[9] ),
    .Y(_03649_));
 sky130_fd_sc_hd__a31o_1 _10567_ (.A1(\div_res[9] ),
    .A2(net165),
    .A3(_03648_),
    .B1(net195),
    .X(_03650_));
 sky130_fd_sc_hd__a21oi_1 _10568_ (.A1(_06307_),
    .A2(_02319_),
    .B1(_02315_),
    .Y(_03651_));
 sky130_fd_sc_hd__or3_1 _10569_ (.A(\div_shifter[40] ),
    .B(\div_shifter[39] ),
    .C(_03388_),
    .X(_03652_));
 sky130_fd_sc_hd__a21oi_1 _10570_ (.A1(net235),
    .A2(_03652_),
    .B1(\div_shifter[41] ),
    .Y(_03653_));
 sky130_fd_sc_hd__a31o_1 _10571_ (.A1(\div_shifter[41] ),
    .A2(net235),
    .A3(_03652_),
    .B1(net193),
    .X(_03654_));
 sky130_fd_sc_hd__o221a_1 _10572_ (.A1(_06291_),
    .A2(net209),
    .B1(_02326_),
    .B2(_06307_),
    .C1(net247),
    .X(_03655_));
 sky130_fd_sc_hd__o221a_1 _10573_ (.A1(_06300_),
    .A2(_03651_),
    .B1(_03653_),
    .B2(_03654_),
    .C1(_03655_),
    .X(_03656_));
 sky130_fd_sc_hd__o21ai_1 _10574_ (.A1(_03649_),
    .A2(_03650_),
    .B1(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__o21a_1 _10575_ (.A1(net227),
    .A2(_03250_),
    .B1(_02335_),
    .X(_03658_));
 sky130_fd_sc_hd__a221o_1 _10576_ (.A1(_02313_),
    .A2(_03646_),
    .B1(_03658_),
    .B2(net179),
    .C1(_03657_),
    .X(_03659_));
 sky130_fd_sc_hd__a211o_1 _10577_ (.A1(net210),
    .A2(_03647_),
    .B1(_03659_),
    .C1(_03639_),
    .X(_03660_));
 sky130_fd_sc_hd__a31o_1 _10578_ (.A1(_02323_),
    .A2(_03634_),
    .A3(_03635_),
    .B1(_03660_),
    .X(_03661_));
 sky130_fd_sc_hd__a31o_1 _10579_ (.A1(net200),
    .A2(_03632_),
    .A3(_03633_),
    .B1(_03661_),
    .X(_03662_));
 sky130_fd_sc_hd__o21a_4 _10580_ (.A1(net243),
    .A2(_03535_),
    .B1(_03662_),
    .X(dest_val[9]));
 sky130_fd_sc_hd__or4b_4 _10581_ (.A(_03368_),
    .B(_03408_),
    .C(_03631_),
    .D_N(_03500_),
    .X(_03663_));
 sky130_fd_sc_hd__o21ai_1 _10582_ (.A1(_03611_),
    .A2(_03612_),
    .B1(_03614_),
    .Y(_03664_));
 sky130_fd_sc_hd__o22a_1 _10583_ (.A1(net77),
    .A2(net24),
    .B1(net16),
    .B2(net73),
    .X(_03665_));
 sky130_fd_sc_hd__xnor2_1 _10584_ (.A(net70),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__a22o_1 _10585_ (.A1(net102),
    .A2(net40),
    .B1(net37),
    .B2(_00189_),
    .X(_03667_));
 sky130_fd_sc_hd__xor2_1 _10586_ (.A(_00245_),
    .B(_03667_),
    .X(_03668_));
 sky130_fd_sc_hd__inv_2 _10587_ (.A(_03668_),
    .Y(_03669_));
 sky130_fd_sc_hd__xnor2_1 _10588_ (.A(_03666_),
    .B(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__a22o_1 _10589_ (.A1(net44),
    .A2(_00348_),
    .B1(_00354_),
    .B2(net41),
    .X(_03671_));
 sky130_fd_sc_hd__xor2_1 _10590_ (.A(net93),
    .B(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__nand2b_1 _10591_ (.A_N(_03670_),
    .B(_03672_),
    .Y(_03673_));
 sky130_fd_sc_hd__nand2b_1 _10592_ (.A_N(_03672_),
    .B(_03670_),
    .Y(_03674_));
 sky130_fd_sc_hd__nand2_1 _10593_ (.A(_03673_),
    .B(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__a21boi_2 _10594_ (.A1(_03557_),
    .A2(_03563_),
    .B1_N(_03562_),
    .Y(_03676_));
 sky130_fd_sc_hd__o22a_1 _10595_ (.A1(net119),
    .A2(net11),
    .B1(net6),
    .B2(_00290_),
    .X(_03677_));
 sky130_fd_sc_hd__xnor2_2 _10596_ (.A(net19),
    .B(_03677_),
    .Y(_03678_));
 sky130_fd_sc_hd__xnor2_2 _10597_ (.A(_03676_),
    .B(_03678_),
    .Y(_03679_));
 sky130_fd_sc_hd__nor2_1 _10598_ (.A(net112),
    .B(net19),
    .Y(_03680_));
 sky130_fd_sc_hd__or3_1 _10599_ (.A(net112),
    .B(net19),
    .C(_03679_),
    .X(_03681_));
 sky130_fd_sc_hd__xnor2_2 _10600_ (.A(_03679_),
    .B(_03680_),
    .Y(_03682_));
 sky130_fd_sc_hd__o22a_1 _10601_ (.A1(net54),
    .A2(net47),
    .B1(net45),
    .B2(net52),
    .X(_03683_));
 sky130_fd_sc_hd__xnor2_1 _10602_ (.A(net96),
    .B(_03683_),
    .Y(_03684_));
 sky130_fd_sc_hd__o22a_1 _10603_ (.A1(net60),
    .A2(net28),
    .B1(net26),
    .B2(net58),
    .X(_03685_));
 sky130_fd_sc_hd__xnor2_1 _10604_ (.A(_00301_),
    .B(_03685_),
    .Y(_03686_));
 sky130_fd_sc_hd__and2_1 _10605_ (.A(_03684_),
    .B(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__xor2_1 _10606_ (.A(_03684_),
    .B(_03686_),
    .X(_03688_));
 sky130_fd_sc_hd__a22o_1 _10607_ (.A1(_06540_),
    .A2(net32),
    .B1(net30),
    .B2(_06547_),
    .X(_03689_));
 sky130_fd_sc_hd__xnor2_1 _10608_ (.A(net50),
    .B(_03689_),
    .Y(_03690_));
 sky130_fd_sc_hd__xor2_1 _10609_ (.A(_03688_),
    .B(_03690_),
    .X(_03691_));
 sky130_fd_sc_hd__nand2_1 _10610_ (.A(_03682_),
    .B(_03691_),
    .Y(_03692_));
 sky130_fd_sc_hd__xnor2_1 _10611_ (.A(_03682_),
    .B(_03691_),
    .Y(_03693_));
 sky130_fd_sc_hd__xor2_1 _10612_ (.A(_03675_),
    .B(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__a21o_1 _10613_ (.A1(_03594_),
    .A2(_03596_),
    .B1(_03592_),
    .X(_03695_));
 sky130_fd_sc_hd__o21ai_1 _10614_ (.A1(net104),
    .A2(net7),
    .B1(_00342_),
    .Y(_03696_));
 sky130_fd_sc_hd__o31a_2 _10615_ (.A1(_00342_),
    .A2(_00389_),
    .A3(_02067_),
    .B1(_03696_),
    .X(_03697_));
 sky130_fd_sc_hd__xnor2_1 _10616_ (.A(_03695_),
    .B(_03697_),
    .Y(_03698_));
 sky130_fd_sc_hd__a21oi_1 _10617_ (.A1(_03543_),
    .A2(_03547_),
    .B1(_03698_),
    .Y(_03699_));
 sky130_fd_sc_hd__and3_1 _10618_ (.A(_03543_),
    .B(_03547_),
    .C(_03698_),
    .X(_03700_));
 sky130_fd_sc_hd__nor2_1 _10619_ (.A(_03699_),
    .B(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__xnor2_1 _10620_ (.A(_03694_),
    .B(_03701_),
    .Y(_03702_));
 sky130_fd_sc_hd__o21ba_1 _10621_ (.A1(_03436_),
    .A2(_03585_),
    .B1_N(_03584_),
    .X(_03703_));
 sky130_fd_sc_hd__o22a_1 _10622_ (.A1(net83),
    .A2(net14),
    .B1(net12),
    .B2(net87),
    .X(_03704_));
 sky130_fd_sc_hd__xnor2_2 _10623_ (.A(net137),
    .B(_03704_),
    .Y(_03705_));
 sky130_fd_sc_hd__o22a_1 _10624_ (.A1(net67),
    .A2(net36),
    .B1(net34),
    .B2(net66),
    .X(_03706_));
 sky130_fd_sc_hd__xnor2_1 _10625_ (.A(net124),
    .B(_03706_),
    .Y(_03707_));
 sky130_fd_sc_hd__nor2_1 _10626_ (.A(_03705_),
    .B(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__xnor2_1 _10627_ (.A(_03705_),
    .B(_03707_),
    .Y(_03709_));
 sky130_fd_sc_hd__o22a_1 _10628_ (.A1(net55),
    .A2(net75),
    .B1(net17),
    .B2(net79),
    .X(_03710_));
 sky130_fd_sc_hd__xnor2_1 _10629_ (.A(net122),
    .B(_03710_),
    .Y(_03711_));
 sky130_fd_sc_hd__nor2_1 _10630_ (.A(_03709_),
    .B(_03711_),
    .Y(_03712_));
 sky130_fd_sc_hd__and2_1 _10631_ (.A(_03709_),
    .B(_03711_),
    .X(_03713_));
 sky130_fd_sc_hd__or2_1 _10632_ (.A(_03712_),
    .B(_03713_),
    .X(_03714_));
 sky130_fd_sc_hd__a21oi_1 _10633_ (.A1(_03577_),
    .A2(_03580_),
    .B1(_03714_),
    .Y(_03715_));
 sky130_fd_sc_hd__and3_1 _10634_ (.A(_03577_),
    .B(_03580_),
    .C(_03714_),
    .X(_03716_));
 sky130_fd_sc_hd__nor2_1 _10635_ (.A(_03715_),
    .B(_03716_),
    .Y(_03717_));
 sky130_fd_sc_hd__xnor2_1 _10636_ (.A(_03703_),
    .B(_03717_),
    .Y(_03718_));
 sky130_fd_sc_hd__and2b_1 _10637_ (.A_N(_03702_),
    .B(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__xnor2_1 _10638_ (.A(_03702_),
    .B(_03718_),
    .Y(_03720_));
 sky130_fd_sc_hd__a21bo_1 _10639_ (.A1(_03554_),
    .A2(_03601_),
    .B1_N(_03600_),
    .X(_03721_));
 sky130_fd_sc_hd__a21o_1 _10640_ (.A1(_03606_),
    .A2(_03610_),
    .B1(_03609_),
    .X(_03722_));
 sky130_fd_sc_hd__o21ai_1 _10641_ (.A1(_03555_),
    .A2(_03568_),
    .B1(_03567_),
    .Y(_03723_));
 sky130_fd_sc_hd__a32o_1 _10642_ (.A1(_03580_),
    .A2(_03581_),
    .A3(_03598_),
    .B1(_03597_),
    .B2(_03587_),
    .X(_03724_));
 sky130_fd_sc_hd__xor2_1 _10643_ (.A(_03723_),
    .B(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__o21ai_1 _10644_ (.A1(_03550_),
    .A2(_03553_),
    .B1(_03725_),
    .Y(_03726_));
 sky130_fd_sc_hd__or3_1 _10645_ (.A(_03550_),
    .B(_03553_),
    .C(_03725_),
    .X(_03727_));
 sky130_fd_sc_hd__and2_1 _10646_ (.A(_03726_),
    .B(_03727_),
    .X(_03728_));
 sky130_fd_sc_hd__xnor2_1 _10647_ (.A(_03722_),
    .B(_03728_),
    .Y(_03729_));
 sky130_fd_sc_hd__nand2b_1 _10648_ (.A_N(_03729_),
    .B(_03721_),
    .Y(_03730_));
 sky130_fd_sc_hd__xnor2_1 _10649_ (.A(_03721_),
    .B(_03729_),
    .Y(_03731_));
 sky130_fd_sc_hd__nand2_1 _10650_ (.A(_03720_),
    .B(_03731_),
    .Y(_03732_));
 sky130_fd_sc_hd__xnor2_1 _10651_ (.A(_03720_),
    .B(_03731_),
    .Y(_03733_));
 sky130_fd_sc_hd__nand2b_1 _10652_ (.A_N(_03733_),
    .B(_03664_),
    .Y(_03734_));
 sky130_fd_sc_hd__xor2_1 _10653_ (.A(_03664_),
    .B(_03733_),
    .X(_03735_));
 sky130_fd_sc_hd__a21o_2 _10654_ (.A1(_03616_),
    .A2(_03618_),
    .B1(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__nand3_2 _10655_ (.A(_03616_),
    .B(_03618_),
    .C(_03735_),
    .Y(_03737_));
 sky130_fd_sc_hd__nand2_4 _10656_ (.A(_03736_),
    .B(_03737_),
    .Y(_03738_));
 sky130_fd_sc_hd__o21ai_1 _10657_ (.A1(_03418_),
    .A2(_03498_),
    .B1(_03620_),
    .Y(_03739_));
 sky130_fd_sc_hd__and2_1 _10658_ (.A(_03621_),
    .B(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__nor2_1 _10659_ (.A(_03499_),
    .B(_03622_),
    .Y(_03741_));
 sky130_fd_sc_hd__a21oi_1 _10660_ (.A1(_03412_),
    .A2(_03741_),
    .B1(_03740_),
    .Y(_03742_));
 sky130_fd_sc_hd__or4_2 _10661_ (.A(_03222_),
    .B(_03361_),
    .C(_03499_),
    .D(_03622_),
    .X(_03743_));
 sky130_fd_sc_hd__o21bai_2 _10662_ (.A1(_03227_),
    .A2(_03228_),
    .B1_N(_03743_),
    .Y(_03744_));
 sky130_fd_sc_hd__o311ai_4 _10663_ (.A1(_02643_),
    .A2(_03223_),
    .A3(_03743_),
    .B1(_03744_),
    .C1(_03742_),
    .Y(_03745_));
 sky130_fd_sc_hd__xnor2_4 _10664_ (.A(_03738_),
    .B(_03745_),
    .Y(_03746_));
 sky130_fd_sc_hd__a21oi_1 _10665_ (.A1(net161),
    .A2(_03663_),
    .B1(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__a31o_1 _10666_ (.A1(net162),
    .A2(_03663_),
    .A3(_03746_),
    .B1(_02242_),
    .X(_03748_));
 sky130_fd_sc_hd__a22o_1 _10667_ (.A1(net161),
    .A2(_01823_),
    .B1(_01825_),
    .B2(_01826_),
    .X(_03749_));
 sky130_fd_sc_hd__nand4_1 _10668_ (.A(net161),
    .B(_01823_),
    .C(_01825_),
    .D(_01826_),
    .Y(_03750_));
 sky130_fd_sc_hd__nand2_1 _10669_ (.A(_03749_),
    .B(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__o21ai_1 _10670_ (.A1(_06300_),
    .A2(_03636_),
    .B1(_06307_),
    .Y(_03752_));
 sky130_fd_sc_hd__mux2_1 _10671_ (.A0(_06384_),
    .A1(_03752_),
    .S(net285),
    .X(_03753_));
 sky130_fd_sc_hd__nor2_1 _10672_ (.A(_06265_),
    .B(_03753_),
    .Y(_03754_));
 sky130_fd_sc_hd__a21o_1 _10673_ (.A1(_06265_),
    .A2(_03753_),
    .B1(net236),
    .X(_03755_));
 sky130_fd_sc_hd__and2_1 _10674_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .X(_03756_));
 sky130_fd_sc_hd__nand2_1 _10675_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .Y(_03757_));
 sky130_fd_sc_hd__or2_1 _10676_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .X(_03758_));
 sky130_fd_sc_hd__o21ai_1 _10677_ (.A1(_03640_),
    .A2(_03641_),
    .B1(_03642_),
    .Y(_03759_));
 sky130_fd_sc_hd__a21oi_1 _10678_ (.A1(_03757_),
    .A2(_03758_),
    .B1(_03759_),
    .Y(_03760_));
 sky130_fd_sc_hd__and3_1 _10679_ (.A(_03757_),
    .B(_03758_),
    .C(_03759_),
    .X(_03761_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(_02658_),
    .A1(_02664_),
    .S(net222),
    .X(_03762_));
 sky130_fd_sc_hd__inv_2 _10681_ (.A(_03762_),
    .Y(_03763_));
 sky130_fd_sc_hd__mux2_1 _10682_ (.A0(_03102_),
    .A1(_03763_),
    .S(net225),
    .X(_03764_));
 sky130_fd_sc_hd__o21a_1 _10683_ (.A1(_03760_),
    .A2(_03761_),
    .B1(net249),
    .X(_03765_));
 sky130_fd_sc_hd__a211o_1 _10684_ (.A1(net229),
    .A2(_03764_),
    .B1(_03765_),
    .C1(_06476_),
    .X(_03766_));
 sky130_fd_sc_hd__or2_1 _10685_ (.A(\div_res[9] ),
    .B(_03648_),
    .X(_03767_));
 sky130_fd_sc_hd__a21oi_1 _10686_ (.A1(net165),
    .A2(_03767_),
    .B1(\div_res[10] ),
    .Y(_03768_));
 sky130_fd_sc_hd__a31o_1 _10687_ (.A1(\div_res[10] ),
    .A2(net165),
    .A3(_03767_),
    .B1(net195),
    .X(_03769_));
 sky130_fd_sc_hd__mux2_1 _10688_ (.A0(_02320_),
    .A1(_02326_),
    .S(_06256_),
    .X(_03770_));
 sky130_fd_sc_hd__a21oi_1 _10689_ (.A1(net198),
    .A2(_03770_),
    .B1(_06247_),
    .Y(_03771_));
 sky130_fd_sc_hd__or2_1 _10690_ (.A(\div_shifter[41] ),
    .B(_03652_),
    .X(_03772_));
 sky130_fd_sc_hd__a21oi_1 _10691_ (.A1(net234),
    .A2(_03772_),
    .B1(\div_shifter[42] ),
    .Y(_03773_));
 sky130_fd_sc_hd__a311o_1 _10692_ (.A1(\div_shifter[42] ),
    .A2(net234),
    .A3(_03772_),
    .B1(_03773_),
    .C1(net192),
    .X(_03774_));
 sky130_fd_sc_hd__a21oi_1 _10693_ (.A1(_06238_),
    .A2(net241),
    .B1(_03771_),
    .Y(_03775_));
 sky130_fd_sc_hd__o211a_1 _10694_ (.A1(_03768_),
    .A2(_03769_),
    .B1(_03774_),
    .C1(_03775_),
    .X(_03776_));
 sky130_fd_sc_hd__o21ai_2 _10695_ (.A1(net227),
    .A2(_03112_),
    .B1(_02335_),
    .Y(_03777_));
 sky130_fd_sc_hd__o221a_1 _10696_ (.A1(_02314_),
    .A2(_03764_),
    .B1(_03777_),
    .B2(net177),
    .C1(_03776_),
    .X(_03778_));
 sky130_fd_sc_hd__o211a_1 _10697_ (.A1(_03754_),
    .A2(_03755_),
    .B1(_03766_),
    .C1(_03778_),
    .X(_03779_));
 sky130_fd_sc_hd__o221a_1 _10698_ (.A1(_03747_),
    .A2(_03748_),
    .B1(_03751_),
    .B2(_02324_),
    .C1(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__and3_1 _10699_ (.A(curr_PC[9]),
    .B(curr_PC[10]),
    .C(_03532_),
    .X(_03781_));
 sky130_fd_sc_hd__a21oi_1 _10700_ (.A1(curr_PC[9]),
    .A2(_03532_),
    .B1(curr_PC[10]),
    .Y(_03782_));
 sky130_fd_sc_hd__or3_2 _10701_ (.A(net242),
    .B(_03781_),
    .C(_03782_),
    .X(_03783_));
 sky130_fd_sc_hd__o21ai_4 _10702_ (.A1(net248),
    .A2(_03780_),
    .B1(_03783_),
    .Y(dest_val[10]));
 sky130_fd_sc_hd__o21a_1 _10703_ (.A1(_03663_),
    .A2(_03746_),
    .B1(net162),
    .X(_03784_));
 sky130_fd_sc_hd__a21bo_1 _10704_ (.A1(_03722_),
    .A2(_03728_),
    .B1_N(_03730_),
    .X(_03785_));
 sky130_fd_sc_hd__a21oi_1 _10705_ (.A1(_03688_),
    .A2(_03690_),
    .B1(_03687_),
    .Y(_03786_));
 sky130_fd_sc_hd__or2_1 _10706_ (.A(_03697_),
    .B(_03786_),
    .X(_03787_));
 sky130_fd_sc_hd__xor2_1 _10707_ (.A(_03697_),
    .B(_03786_),
    .X(_03788_));
 sky130_fd_sc_hd__o21ai_1 _10708_ (.A1(_03708_),
    .A2(_03712_),
    .B1(_03788_),
    .Y(_03789_));
 sky130_fd_sc_hd__or3_1 _10709_ (.A(_03708_),
    .B(_03712_),
    .C(_03788_),
    .X(_03790_));
 sky130_fd_sc_hd__nand2_1 _10710_ (.A(_03789_),
    .B(_03790_),
    .Y(_03791_));
 sky130_fd_sc_hd__o22a_1 _10711_ (.A1(net62),
    .A2(net47),
    .B1(net45),
    .B2(net54),
    .X(_03792_));
 sky130_fd_sc_hd__xnor2_1 _10712_ (.A(net95),
    .B(_03792_),
    .Y(_03793_));
 sky130_fd_sc_hd__a22o_1 _10713_ (.A1(_00189_),
    .A2(net44),
    .B1(net42),
    .B2(_00348_),
    .X(_03794_));
 sky130_fd_sc_hd__xor2_1 _10714_ (.A(net93),
    .B(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__xor2_1 _10715_ (.A(_03793_),
    .B(_03795_),
    .X(_03796_));
 sky130_fd_sc_hd__a22o_1 _10716_ (.A1(_00172_),
    .A2(net40),
    .B1(net38),
    .B2(net102),
    .X(_03797_));
 sky130_fd_sc_hd__xor2_1 _10717_ (.A(net90),
    .B(_03797_),
    .X(_03798_));
 sky130_fd_sc_hd__and2_1 _10718_ (.A(_03796_),
    .B(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__nor2_1 _10719_ (.A(_03796_),
    .B(_03798_),
    .Y(_03800_));
 sky130_fd_sc_hd__or2_1 _10720_ (.A(_03799_),
    .B(_03800_),
    .X(_03801_));
 sky130_fd_sc_hd__o22a_1 _10721_ (.A1(net73),
    .A2(net11),
    .B1(net6),
    .B2(net120),
    .X(_03802_));
 sky130_fd_sc_hd__xnor2_1 _10722_ (.A(net19),
    .B(_03802_),
    .Y(_03803_));
 sky130_fd_sc_hd__a32o_1 _10723_ (.A1(_00361_),
    .A2(_00686_),
    .A3(_00687_),
    .B1(_00452_),
    .B2(_00354_),
    .X(_03804_));
 sky130_fd_sc_hd__xnor2_1 _10724_ (.A(_00678_),
    .B(_03804_),
    .Y(_03805_));
 sky130_fd_sc_hd__nand2_1 _10725_ (.A(net116),
    .B(_02078_),
    .Y(_03806_));
 sky130_fd_sc_hd__xor2_1 _10726_ (.A(_03805_),
    .B(_03806_),
    .X(_03807_));
 sky130_fd_sc_hd__nand2b_1 _10727_ (.A_N(_03803_),
    .B(_03807_),
    .Y(_03808_));
 sky130_fd_sc_hd__xnor2_1 _10728_ (.A(_03803_),
    .B(_03807_),
    .Y(_03809_));
 sky130_fd_sc_hd__o22a_1 _10729_ (.A1(net55),
    .A2(net36),
    .B1(net34),
    .B2(net67),
    .X(_03810_));
 sky130_fd_sc_hd__xnor2_1 _10730_ (.A(net126),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__a22o_1 _10731_ (.A1(_06563_),
    .A2(net32),
    .B1(net30),
    .B2(_06540_),
    .X(_03812_));
 sky130_fd_sc_hd__xnor2_1 _10732_ (.A(net50),
    .B(_03812_),
    .Y(_03813_));
 sky130_fd_sc_hd__and2_1 _10733_ (.A(_03811_),
    .B(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__xor2_1 _10734_ (.A(_03811_),
    .B(_03813_),
    .X(_03815_));
 sky130_fd_sc_hd__o22a_1 _10735_ (.A1(net66),
    .A2(net28),
    .B1(net26),
    .B2(net60),
    .X(_03816_));
 sky130_fd_sc_hd__xnor2_1 _10736_ (.A(net89),
    .B(_03816_),
    .Y(_03817_));
 sky130_fd_sc_hd__xor2_1 _10737_ (.A(_03815_),
    .B(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__nand2_1 _10738_ (.A(_03809_),
    .B(_03818_),
    .Y(_03819_));
 sky130_fd_sc_hd__or2_1 _10739_ (.A(_03809_),
    .B(_03818_),
    .X(_03820_));
 sky130_fd_sc_hd__nand2_1 _10740_ (.A(_03819_),
    .B(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__xnor2_1 _10741_ (.A(_03801_),
    .B(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__xnor2_1 _10742_ (.A(_03791_),
    .B(_03822_),
    .Y(_03823_));
 sky130_fd_sc_hd__o21ai_2 _10743_ (.A1(_03676_),
    .A2(_03678_),
    .B1(_03681_),
    .Y(_03824_));
 sky130_fd_sc_hd__o22a_1 _10744_ (.A1(net83),
    .A2(net12),
    .B1(net7),
    .B2(net87),
    .X(_03825_));
 sky130_fd_sc_hd__xnor2_1 _10745_ (.A(_00339_),
    .B(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__o22a_1 _10746_ (.A1(net75),
    .A2(net17),
    .B1(net14),
    .B2(net79),
    .X(_03827_));
 sky130_fd_sc_hd__xnor2_1 _10747_ (.A(net122),
    .B(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__nor2_1 _10748_ (.A(_00342_),
    .B(_03828_),
    .Y(_03829_));
 sky130_fd_sc_hd__xnor2_1 _10749_ (.A(net135),
    .B(_03828_),
    .Y(_03830_));
 sky130_fd_sc_hd__and2_1 _10750_ (.A(_03826_),
    .B(_03830_),
    .X(_03831_));
 sky130_fd_sc_hd__nor2_1 _10751_ (.A(_03826_),
    .B(_03830_),
    .Y(_03832_));
 sky130_fd_sc_hd__nor2_1 _10752_ (.A(_03831_),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__o21ai_1 _10753_ (.A1(_03666_),
    .A2(_03669_),
    .B1(_03673_),
    .Y(_03834_));
 sky130_fd_sc_hd__and2_1 _10754_ (.A(_03833_),
    .B(_03834_),
    .X(_03835_));
 sky130_fd_sc_hd__xor2_1 _10755_ (.A(_03833_),
    .B(_03834_),
    .X(_03836_));
 sky130_fd_sc_hd__xnor2_1 _10756_ (.A(_03824_),
    .B(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__or2_1 _10757_ (.A(_03823_),
    .B(_03837_),
    .X(_03838_));
 sky130_fd_sc_hd__nand2_1 _10758_ (.A(_03823_),
    .B(_03837_),
    .Y(_03839_));
 sky130_fd_sc_hd__and2_1 _10759_ (.A(_03838_),
    .B(_03839_),
    .X(_03840_));
 sky130_fd_sc_hd__a21o_1 _10760_ (.A1(_03694_),
    .A2(_03701_),
    .B1(_03719_),
    .X(_03841_));
 sky130_fd_sc_hd__o21bai_2 _10761_ (.A1(_03703_),
    .A2(_03716_),
    .B1_N(_03715_),
    .Y(_03842_));
 sky130_fd_sc_hd__o21a_1 _10762_ (.A1(_03675_),
    .A2(_03693_),
    .B1(_03692_),
    .X(_03843_));
 sky130_fd_sc_hd__a21o_1 _10763_ (.A1(_03695_),
    .A2(_03697_),
    .B1(_03699_),
    .X(_03844_));
 sky130_fd_sc_hd__nand2b_1 _10764_ (.A_N(_03843_),
    .B(_03844_),
    .Y(_03845_));
 sky130_fd_sc_hd__xnor2_1 _10765_ (.A(_03843_),
    .B(_03844_),
    .Y(_03846_));
 sky130_fd_sc_hd__xnor2_1 _10766_ (.A(_03842_),
    .B(_03846_),
    .Y(_03847_));
 sky130_fd_sc_hd__a21boi_1 _10767_ (.A1(_03723_),
    .A2(_03724_),
    .B1_N(_03726_),
    .Y(_03848_));
 sky130_fd_sc_hd__xnor2_1 _10768_ (.A(_03847_),
    .B(_03848_),
    .Y(_03849_));
 sky130_fd_sc_hd__nand2b_1 _10769_ (.A_N(_03849_),
    .B(_03841_),
    .Y(_03850_));
 sky130_fd_sc_hd__xnor2_1 _10770_ (.A(_03841_),
    .B(_03849_),
    .Y(_03851_));
 sky130_fd_sc_hd__nand2_1 _10771_ (.A(_03840_),
    .B(_03851_),
    .Y(_03852_));
 sky130_fd_sc_hd__xnor2_1 _10772_ (.A(_03840_),
    .B(_03851_),
    .Y(_03853_));
 sky130_fd_sc_hd__nand2b_1 _10773_ (.A_N(_03853_),
    .B(_03785_),
    .Y(_03854_));
 sky130_fd_sc_hd__xor2_1 _10774_ (.A(_03785_),
    .B(_03853_),
    .X(_03855_));
 sky130_fd_sc_hd__a21oi_1 _10775_ (.A1(_03732_),
    .A2(_03734_),
    .B1(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__a21o_1 _10776_ (.A1(_03732_),
    .A2(_03734_),
    .B1(_03855_),
    .X(_03857_));
 sky130_fd_sc_hd__and3_1 _10777_ (.A(_03732_),
    .B(_03734_),
    .C(_03855_),
    .X(_03858_));
 sky130_fd_sc_hd__or2_4 _10778_ (.A(_03856_),
    .B(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__nor2_1 _10779_ (.A(_03622_),
    .B(_03738_),
    .Y(_03860_));
 sky130_fd_sc_hd__and2_1 _10780_ (.A(_03623_),
    .B(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__a21boi_1 _10781_ (.A1(_03620_),
    .A2(_03736_),
    .B1_N(_03737_),
    .Y(_03862_));
 sky130_fd_sc_hd__a21o_1 _10782_ (.A1(_03628_),
    .A2(_03860_),
    .B1(_03862_),
    .X(_03863_));
 sky130_fd_sc_hd__a21o_2 _10783_ (.A1(_03367_),
    .A2(_03861_),
    .B1(_03863_),
    .X(_03864_));
 sky130_fd_sc_hd__xnor2_4 _10784_ (.A(_03859_),
    .B(_03864_),
    .Y(_03865_));
 sky130_fd_sc_hd__o21ai_1 _10785_ (.A1(_03784_),
    .A2(_03865_),
    .B1(net200),
    .Y(_03866_));
 sky130_fd_sc_hd__a21oi_1 _10786_ (.A1(_03784_),
    .A2(_03865_),
    .B1(_03866_),
    .Y(_03867_));
 sky130_fd_sc_hd__o21a_1 _10787_ (.A1(net157),
    .A2(_01827_),
    .B1(_01829_),
    .X(_03868_));
 sky130_fd_sc_hd__nor2_1 _10788_ (.A(_02324_),
    .B(_03868_),
    .Y(_03869_));
 sky130_fd_sc_hd__o31a_1 _10789_ (.A1(net157),
    .A2(_01827_),
    .A3(_01829_),
    .B1(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__a21o_1 _10790_ (.A1(_06265_),
    .A2(_03752_),
    .B1(_06256_),
    .X(_03871_));
 sky130_fd_sc_hd__nand2_1 _10791_ (.A(net284),
    .B(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__o21ai_1 _10792_ (.A1(net285),
    .A2(_06386_),
    .B1(_03872_),
    .Y(_03873_));
 sky130_fd_sc_hd__o21ai_1 _10793_ (.A1(_06211_),
    .A2(_03873_),
    .B1(_02317_),
    .Y(_03874_));
 sky130_fd_sc_hd__a21oi_1 _10794_ (.A1(_06211_),
    .A2(_03873_),
    .B1(_03874_),
    .Y(_03875_));
 sky130_fd_sc_hd__and2_1 _10795_ (.A(reg1_val[11]),
    .B(curr_PC[11]),
    .X(_03876_));
 sky130_fd_sc_hd__nand2_1 _10796_ (.A(reg1_val[11]),
    .B(curr_PC[11]),
    .Y(_03877_));
 sky130_fd_sc_hd__or2_1 _10797_ (.A(reg1_val[11]),
    .B(curr_PC[11]),
    .X(_03878_));
 sky130_fd_sc_hd__a211o_1 _10798_ (.A1(_03877_),
    .A2(_03878_),
    .B1(_03756_),
    .C1(_03761_),
    .X(_03879_));
 sky130_fd_sc_hd__o211a_1 _10799_ (.A1(_03756_),
    .A2(_03761_),
    .B1(_03877_),
    .C1(_03878_),
    .X(_03880_));
 sky130_fd_sc_hd__or3b_1 _10800_ (.A(_03880_),
    .B(net229),
    .C_N(_03879_),
    .X(_03881_));
 sky130_fd_sc_hd__mux2_1 _10801_ (.A0(_02812_),
    .A1(_02818_),
    .S(net222),
    .X(_03882_));
 sky130_fd_sc_hd__inv_2 _10802_ (.A(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__mux2_1 _10803_ (.A0(_02967_),
    .A1(_03883_),
    .S(net225),
    .X(_03884_));
 sky130_fd_sc_hd__o21a_1 _10804_ (.A1(net249),
    .A2(_03884_),
    .B1(_03881_),
    .X(_03885_));
 sky130_fd_sc_hd__or2_1 _10805_ (.A(\div_res[10] ),
    .B(_03767_),
    .X(_03886_));
 sky130_fd_sc_hd__a21oi_1 _10806_ (.A1(net165),
    .A2(_03886_),
    .B1(\div_res[11] ),
    .Y(_03887_));
 sky130_fd_sc_hd__a31o_1 _10807_ (.A1(\div_res[11] ),
    .A2(net165),
    .A3(_03886_),
    .B1(net195),
    .X(_03888_));
 sky130_fd_sc_hd__mux2_1 _10808_ (.A0(net197),
    .A1(net196),
    .S(_06193_),
    .X(_03889_));
 sky130_fd_sc_hd__a21o_1 _10809_ (.A1(net198),
    .A2(_03889_),
    .B1(_06202_),
    .X(_03890_));
 sky130_fd_sc_hd__or2_1 _10810_ (.A(\div_shifter[42] ),
    .B(_03772_),
    .X(_03891_));
 sky130_fd_sc_hd__a21oi_1 _10811_ (.A1(net234),
    .A2(_03891_),
    .B1(\div_shifter[43] ),
    .Y(_03892_));
 sky130_fd_sc_hd__a31o_1 _10812_ (.A1(\div_shifter[43] ),
    .A2(net234),
    .A3(_03891_),
    .B1(net193),
    .X(_03893_));
 sky130_fd_sc_hd__nand2_1 _10813_ (.A(_06185_),
    .B(net241),
    .Y(_03894_));
 sky130_fd_sc_hd__o211a_1 _10814_ (.A1(_03892_),
    .A2(_03893_),
    .B1(_03894_),
    .C1(_03890_),
    .X(_03895_));
 sky130_fd_sc_hd__o21ai_2 _10815_ (.A1(net226),
    .A2(_02973_),
    .B1(_02335_),
    .Y(_03896_));
 sky130_fd_sc_hd__o221a_1 _10816_ (.A1(_03887_),
    .A2(_03888_),
    .B1(_03896_),
    .B2(net177),
    .C1(_03895_),
    .X(_03897_));
 sky130_fd_sc_hd__o221a_1 _10817_ (.A1(_02314_),
    .A2(_03884_),
    .B1(_03885_),
    .B2(_06476_),
    .C1(_03897_),
    .X(_03898_));
 sky130_fd_sc_hd__or4b_1 _10818_ (.A(_03867_),
    .B(_03870_),
    .C(_03875_),
    .D_N(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__or2_1 _10819_ (.A(curr_PC[11]),
    .B(_03781_),
    .X(_03900_));
 sky130_fd_sc_hd__and2_1 _10820_ (.A(curr_PC[11]),
    .B(_03781_),
    .X(_03901_));
 sky130_fd_sc_hd__nor2_1 _10821_ (.A(net242),
    .B(_03901_),
    .Y(_03902_));
 sky130_fd_sc_hd__a22o_4 _10822_ (.A1(net242),
    .A2(_03899_),
    .B1(_03900_),
    .B2(_03902_),
    .X(dest_val[11]));
 sky130_fd_sc_hd__or3_1 _10823_ (.A(_03663_),
    .B(_03746_),
    .C(_03865_),
    .X(_03903_));
 sky130_fd_sc_hd__and2_1 _10824_ (.A(net162),
    .B(_03903_),
    .X(_03904_));
 sky130_fd_sc_hd__o21ai_1 _10825_ (.A1(_03847_),
    .A2(_03848_),
    .B1(_03850_),
    .Y(_03905_));
 sky130_fd_sc_hd__o21ai_1 _10826_ (.A1(_03805_),
    .A2(_03806_),
    .B1(_03808_),
    .Y(_03906_));
 sky130_fd_sc_hd__a21o_1 _10827_ (.A1(_03793_),
    .A2(_03795_),
    .B1(_03799_),
    .X(_03907_));
 sky130_fd_sc_hd__o22a_1 _10828_ (.A1(net75),
    .A2(net14),
    .B1(net12),
    .B2(net78),
    .X(_03908_));
 sky130_fd_sc_hd__xnor2_2 _10829_ (.A(net122),
    .B(_03908_),
    .Y(_03909_));
 sky130_fd_sc_hd__inv_2 _10830_ (.A(_03909_),
    .Y(_03910_));
 sky130_fd_sc_hd__o21ai_1 _10831_ (.A1(_00345_),
    .A2(net7),
    .B1(_00339_),
    .Y(_03911_));
 sky130_fd_sc_hd__o31ai_2 _10832_ (.A1(_00339_),
    .A2(_00346_),
    .A3(_02067_),
    .B1(_03911_),
    .Y(_03912_));
 sky130_fd_sc_hd__nor2_1 _10833_ (.A(_03910_),
    .B(_03912_),
    .Y(_03913_));
 sky130_fd_sc_hd__xnor2_1 _10834_ (.A(_03909_),
    .B(_03912_),
    .Y(_03914_));
 sky130_fd_sc_hd__inv_2 _10835_ (.A(_03914_),
    .Y(_03915_));
 sky130_fd_sc_hd__xnor2_1 _10836_ (.A(_03907_),
    .B(_03915_),
    .Y(_03916_));
 sky130_fd_sc_hd__nand2b_1 _10837_ (.A_N(_03916_),
    .B(_03906_),
    .Y(_03917_));
 sky130_fd_sc_hd__xnor2_1 _10838_ (.A(_03906_),
    .B(_03916_),
    .Y(_03918_));
 sky130_fd_sc_hd__a22o_1 _10839_ (.A1(net102),
    .A2(net43),
    .B1(net42),
    .B2(_00189_),
    .X(_03919_));
 sky130_fd_sc_hd__xor2_1 _10840_ (.A(net93),
    .B(_03919_),
    .X(_03920_));
 sky130_fd_sc_hd__o22a_1 _10841_ (.A1(net64),
    .A2(net47),
    .B1(net45),
    .B2(net62),
    .X(_03921_));
 sky130_fd_sc_hd__xnor2_1 _10842_ (.A(net95),
    .B(_03921_),
    .Y(_03922_));
 sky130_fd_sc_hd__and2_1 _10843_ (.A(_03920_),
    .B(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__nor2_1 _10844_ (.A(_03920_),
    .B(_03922_),
    .Y(_03924_));
 sky130_fd_sc_hd__nor2_1 _10845_ (.A(_03923_),
    .B(_03924_),
    .Y(_03925_));
 sky130_fd_sc_hd__a22o_1 _10846_ (.A1(_00163_),
    .A2(net40),
    .B1(net38),
    .B2(_00172_),
    .X(_03926_));
 sky130_fd_sc_hd__xor2_1 _10847_ (.A(net90),
    .B(_03926_),
    .X(_03927_));
 sky130_fd_sc_hd__xnor2_1 _10848_ (.A(_03925_),
    .B(_03927_),
    .Y(_03928_));
 sky130_fd_sc_hd__o32a_1 _10849_ (.A1(net36),
    .A2(_00405_),
    .A3(_00407_),
    .B1(net34),
    .B2(net55),
    .X(_03929_));
 sky130_fd_sc_hd__xnor2_1 _10850_ (.A(net126),
    .B(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__a22o_1 _10851_ (.A1(_06559_),
    .A2(net32),
    .B1(net30),
    .B2(_06563_),
    .X(_03931_));
 sky130_fd_sc_hd__xnor2_1 _10852_ (.A(net50),
    .B(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__nand2_1 _10853_ (.A(_03930_),
    .B(_03932_),
    .Y(_03933_));
 sky130_fd_sc_hd__xor2_1 _10854_ (.A(_03930_),
    .B(_03932_),
    .X(_03934_));
 sky130_fd_sc_hd__o22a_1 _10855_ (.A1(net67),
    .A2(net28),
    .B1(net26),
    .B2(net66),
    .X(_03935_));
 sky130_fd_sc_hd__xnor2_1 _10856_ (.A(net89),
    .B(_03935_),
    .Y(_03936_));
 sky130_fd_sc_hd__nand2_1 _10857_ (.A(_03934_),
    .B(_03936_),
    .Y(_03937_));
 sky130_fd_sc_hd__xor2_1 _10858_ (.A(_03934_),
    .B(_03936_),
    .X(_03938_));
 sky130_fd_sc_hd__o22a_1 _10859_ (.A1(net85),
    .A2(net24),
    .B1(net16),
    .B2(net81),
    .X(_03939_));
 sky130_fd_sc_hd__xnor2_1 _10860_ (.A(net70),
    .B(_03939_),
    .Y(_03940_));
 sky130_fd_sc_hd__o22a_1 _10861_ (.A1(net77),
    .A2(net10),
    .B1(net5),
    .B2(net73),
    .X(_03941_));
 sky130_fd_sc_hd__xnor2_1 _10862_ (.A(net20),
    .B(_03941_),
    .Y(_03942_));
 sky130_fd_sc_hd__or2_1 _10863_ (.A(_03940_),
    .B(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__xor2_1 _10864_ (.A(_03940_),
    .B(_03942_),
    .X(_03944_));
 sky130_fd_sc_hd__nand2_1 _10865_ (.A(_03938_),
    .B(_03944_),
    .Y(_03945_));
 sky130_fd_sc_hd__xnor2_1 _10866_ (.A(_03938_),
    .B(_03944_),
    .Y(_03946_));
 sky130_fd_sc_hd__or2_1 _10867_ (.A(_03928_),
    .B(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__nand2_1 _10868_ (.A(_03928_),
    .B(_03946_),
    .Y(_03948_));
 sky130_fd_sc_hd__nand2_1 _10869_ (.A(_03947_),
    .B(_03948_),
    .Y(_03949_));
 sky130_fd_sc_hd__a21oi_1 _10870_ (.A1(_03815_),
    .A2(_03817_),
    .B1(_03814_),
    .Y(_03950_));
 sky130_fd_sc_hd__nor2_1 _10871_ (.A(net120),
    .B(net19),
    .Y(_03951_));
 sky130_fd_sc_hd__xnor2_1 _10872_ (.A(_03950_),
    .B(_03951_),
    .Y(_03952_));
 sky130_fd_sc_hd__o21ai_1 _10873_ (.A1(_03829_),
    .A2(_03831_),
    .B1(_03952_),
    .Y(_03953_));
 sky130_fd_sc_hd__or3_1 _10874_ (.A(_03829_),
    .B(_03831_),
    .C(_03952_),
    .X(_03954_));
 sky130_fd_sc_hd__nand2_1 _10875_ (.A(_03953_),
    .B(_03954_),
    .Y(_03955_));
 sky130_fd_sc_hd__nor2_1 _10876_ (.A(_03949_),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__and2_1 _10877_ (.A(_03949_),
    .B(_03955_),
    .X(_03957_));
 sky130_fd_sc_hd__nor2_1 _10878_ (.A(_03956_),
    .B(_03957_),
    .Y(_03958_));
 sky130_fd_sc_hd__xor2_1 _10879_ (.A(_03918_),
    .B(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__o21a_1 _10880_ (.A1(_03791_),
    .A2(_03822_),
    .B1(_03838_),
    .X(_03960_));
 sky130_fd_sc_hd__a21o_1 _10881_ (.A1(_03824_),
    .A2(_03836_),
    .B1(_03835_),
    .X(_03961_));
 sky130_fd_sc_hd__nand2_1 _10882_ (.A(_03787_),
    .B(_03789_),
    .Y(_03962_));
 sky130_fd_sc_hd__o21a_1 _10883_ (.A1(_03801_),
    .A2(_03821_),
    .B1(_03819_),
    .X(_03963_));
 sky130_fd_sc_hd__a21oi_1 _10884_ (.A1(_03787_),
    .A2(_03789_),
    .B1(_03963_),
    .Y(_03964_));
 sky130_fd_sc_hd__xnor2_1 _10885_ (.A(_03962_),
    .B(_03963_),
    .Y(_03965_));
 sky130_fd_sc_hd__xnor2_1 _10886_ (.A(_03961_),
    .B(_03965_),
    .Y(_03966_));
 sky130_fd_sc_hd__a21boi_1 _10887_ (.A1(_03842_),
    .A2(_03846_),
    .B1_N(_03845_),
    .Y(_03967_));
 sky130_fd_sc_hd__xor2_1 _10888_ (.A(_03966_),
    .B(_03967_),
    .X(_03968_));
 sky130_fd_sc_hd__nand2b_1 _10889_ (.A_N(_03960_),
    .B(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hd__xnor2_1 _10890_ (.A(_03960_),
    .B(_03968_),
    .Y(_03970_));
 sky130_fd_sc_hd__nand2_1 _10891_ (.A(_03959_),
    .B(_03970_),
    .Y(_03971_));
 sky130_fd_sc_hd__xor2_1 _10892_ (.A(_03959_),
    .B(_03970_),
    .X(_03972_));
 sky130_fd_sc_hd__nand2_1 _10893_ (.A(_03905_),
    .B(_03972_),
    .Y(_03973_));
 sky130_fd_sc_hd__xnor2_1 _10894_ (.A(_03905_),
    .B(_03972_),
    .Y(_03974_));
 sky130_fd_sc_hd__a21oi_1 _10895_ (.A1(_03852_),
    .A2(_03854_),
    .B1(_03974_),
    .Y(_03975_));
 sky130_fd_sc_hd__a21o_1 _10896_ (.A1(_03852_),
    .A2(_03854_),
    .B1(_03974_),
    .X(_03976_));
 sky130_fd_sc_hd__and3_1 _10897_ (.A(_03852_),
    .B(_03854_),
    .C(_03974_),
    .X(_03977_));
 sky130_fd_sc_hd__or2_4 _10898_ (.A(_03975_),
    .B(_03977_),
    .X(_03978_));
 sky130_fd_sc_hd__a21oi_2 _10899_ (.A1(_03736_),
    .A2(_03857_),
    .B1(_03858_),
    .Y(_03979_));
 sky130_fd_sc_hd__nor2_1 _10900_ (.A(_03738_),
    .B(_03859_),
    .Y(_03980_));
 sky130_fd_sc_hd__a21o_1 _10901_ (.A1(_03740_),
    .A2(_03980_),
    .B1(_03979_),
    .X(_03981_));
 sky130_fd_sc_hd__and2_1 _10902_ (.A(_03741_),
    .B(_03980_),
    .X(_03982_));
 sky130_fd_sc_hd__a21o_2 _10903_ (.A1(_03417_),
    .A2(_03982_),
    .B1(_03981_),
    .X(_03983_));
 sky130_fd_sc_hd__xnor2_4 _10904_ (.A(_03978_),
    .B(_03983_),
    .Y(_03984_));
 sky130_fd_sc_hd__a21oi_1 _10905_ (.A1(_03904_),
    .A2(_03984_),
    .B1(_02242_),
    .Y(_03985_));
 sky130_fd_sc_hd__o21a_1 _10906_ (.A1(_03904_),
    .A2(_03984_),
    .B1(_03985_),
    .X(_03986_));
 sky130_fd_sc_hd__a21oi_1 _10907_ (.A1(net161),
    .A2(_01830_),
    .B1(_01835_),
    .Y(_03987_));
 sky130_fd_sc_hd__a311oi_1 _10908_ (.A1(net161),
    .A2(_01830_),
    .A3(_01835_),
    .B1(_02324_),
    .C1(_03987_),
    .Y(_03988_));
 sky130_fd_sc_hd__a21oi_1 _10909_ (.A1(_06211_),
    .A2(_03871_),
    .B1(_06193_),
    .Y(_03989_));
 sky130_fd_sc_hd__mux2_1 _10910_ (.A0(_06388_),
    .A1(_03989_),
    .S(net284),
    .X(_03990_));
 sky130_fd_sc_hd__a21oi_1 _10911_ (.A1(_06169_),
    .A2(_03990_),
    .B1(net236),
    .Y(_03991_));
 sky130_fd_sc_hd__o21a_1 _10912_ (.A1(_06169_),
    .A2(_03990_),
    .B1(_03991_),
    .X(_03992_));
 sky130_fd_sc_hd__mux2_1 _10913_ (.A0(_02970_),
    .A1(_02972_),
    .S(net222),
    .X(_03993_));
 sky130_fd_sc_hd__mux2_1 _10914_ (.A0(_02829_),
    .A1(_03993_),
    .S(net225),
    .X(_03994_));
 sky130_fd_sc_hd__nand2_1 _10915_ (.A(reg1_val[12]),
    .B(curr_PC[12]),
    .Y(_03995_));
 sky130_fd_sc_hd__or2_1 _10916_ (.A(reg1_val[12]),
    .B(curr_PC[12]),
    .X(_03996_));
 sky130_fd_sc_hd__o211a_1 _10917_ (.A1(_03876_),
    .A2(_03880_),
    .B1(_03995_),
    .C1(_03996_),
    .X(_03997_));
 sky130_fd_sc_hd__a211o_1 _10918_ (.A1(_03995_),
    .A2(_03996_),
    .B1(_03876_),
    .C1(_03880_),
    .X(_03998_));
 sky130_fd_sc_hd__nand2_1 _10919_ (.A(net249),
    .B(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hd__a2bb2o_1 _10920_ (.A1_N(_03997_),
    .A2_N(_03999_),
    .B1(net229),
    .B2(_03994_),
    .X(_04000_));
 sky130_fd_sc_hd__or2_1 _10921_ (.A(\div_res[11] ),
    .B(_03886_),
    .X(_04001_));
 sky130_fd_sc_hd__a21o_1 _10922_ (.A1(net165),
    .A2(_04001_),
    .B1(\div_res[12] ),
    .X(_04002_));
 sky130_fd_sc_hd__a31oi_1 _10923_ (.A1(\div_res[12] ),
    .A2(net165),
    .A3(_04001_),
    .B1(net194),
    .Y(_04003_));
 sky130_fd_sc_hd__or2_1 _10924_ (.A(\div_shifter[43] ),
    .B(_03891_),
    .X(_04004_));
 sky130_fd_sc_hd__a21o_1 _10925_ (.A1(net233),
    .A2(_04004_),
    .B1(\div_shifter[44] ),
    .X(_04005_));
 sky130_fd_sc_hd__a31oi_1 _10926_ (.A1(\div_shifter[44] ),
    .A2(net233),
    .A3(_04004_),
    .B1(net192),
    .Y(_04006_));
 sky130_fd_sc_hd__mux2_1 _10927_ (.A0(net197),
    .A1(net196),
    .S(_06157_),
    .X(_04007_));
 sky130_fd_sc_hd__a21oi_1 _10928_ (.A1(net199),
    .A2(_04007_),
    .B1(_06163_),
    .Y(_04008_));
 sky130_fd_sc_hd__a221o_1 _10929_ (.A1(_06151_),
    .A2(net241),
    .B1(_04005_),
    .B2(_04006_),
    .C1(_04008_),
    .X(_04009_));
 sky130_fd_sc_hd__o21a_1 _10930_ (.A1(net226),
    .A2(_02819_),
    .B1(_02335_),
    .X(_04010_));
 sky130_fd_sc_hd__a221o_1 _10931_ (.A1(_04002_),
    .A2(_04003_),
    .B1(_04010_),
    .B2(net179),
    .C1(_04009_),
    .X(_04011_));
 sky130_fd_sc_hd__a221o_1 _10932_ (.A1(_02313_),
    .A2(_03994_),
    .B1(_04000_),
    .B2(net210),
    .C1(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__or4_1 _10933_ (.A(_03986_),
    .B(_03988_),
    .C(_03992_),
    .D(_04012_),
    .X(_04013_));
 sky130_fd_sc_hd__and3_1 _10934_ (.A(curr_PC[11]),
    .B(curr_PC[12]),
    .C(_03781_),
    .X(_04014_));
 sky130_fd_sc_hd__o21ai_1 _10935_ (.A1(curr_PC[12]),
    .A2(_03901_),
    .B1(net248),
    .Y(_04015_));
 sky130_fd_sc_hd__a2bb2o_4 _10936_ (.A1_N(_04014_),
    .A2_N(_04015_),
    .B1(net242),
    .B2(_04013_),
    .X(dest_val[12]));
 sky130_fd_sc_hd__o21a_1 _10937_ (.A1(_03903_),
    .A2(_03984_),
    .B1(net162),
    .X(_04016_));
 sky130_fd_sc_hd__o22a_1 _10938_ (.A1(net99),
    .A2(net24),
    .B1(net16),
    .B2(net85),
    .X(_04017_));
 sky130_fd_sc_hd__xnor2_1 _10939_ (.A(net69),
    .B(_04017_),
    .Y(_04018_));
 sky130_fd_sc_hd__a22o_1 _10940_ (.A1(_06547_),
    .A2(net40),
    .B1(net38),
    .B2(_00163_),
    .X(_04019_));
 sky130_fd_sc_hd__xor2_1 _10941_ (.A(net90),
    .B(_04019_),
    .X(_04020_));
 sky130_fd_sc_hd__nand2b_1 _10942_ (.A_N(_04018_),
    .B(_04020_),
    .Y(_04021_));
 sky130_fd_sc_hd__xor2_1 _10943_ (.A(_04018_),
    .B(_04020_),
    .X(_04022_));
 sky130_fd_sc_hd__a22o_1 _10944_ (.A1(_00172_),
    .A2(net43),
    .B1(net41),
    .B2(net102),
    .X(_04023_));
 sky130_fd_sc_hd__xor2_1 _10945_ (.A(net92),
    .B(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__nand2b_1 _10946_ (.A_N(_04022_),
    .B(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__xnor2_1 _10947_ (.A(_04022_),
    .B(_04024_),
    .Y(_04026_));
 sky130_fd_sc_hd__o22a_1 _10948_ (.A1(net34),
    .A2(net17),
    .B1(net14),
    .B2(net36),
    .X(_04027_));
 sky130_fd_sc_hd__xnor2_2 _10949_ (.A(net126),
    .B(_04027_),
    .Y(_04028_));
 sky130_fd_sc_hd__xnor2_2 _10950_ (.A(_00339_),
    .B(_04028_),
    .Y(_04029_));
 sky130_fd_sc_hd__o22a_1 _10951_ (.A1(net75),
    .A2(net12),
    .B1(_02067_),
    .B2(net78),
    .X(_04030_));
 sky130_fd_sc_hd__xor2_2 _10952_ (.A(net122),
    .B(_04030_),
    .X(_04031_));
 sky130_fd_sc_hd__and2_1 _10953_ (.A(_04029_),
    .B(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__xor2_2 _10954_ (.A(_04029_),
    .B(_04031_),
    .X(_04033_));
 sky130_fd_sc_hd__nand2_1 _10955_ (.A(_04026_),
    .B(_04033_),
    .Y(_04034_));
 sky130_fd_sc_hd__or2_1 _10956_ (.A(_04026_),
    .B(_04033_),
    .X(_04035_));
 sky130_fd_sc_hd__o22a_1 _10957_ (.A1(net58),
    .A2(net47),
    .B1(net45),
    .B2(net64),
    .X(_04036_));
 sky130_fd_sc_hd__xnor2_1 _10958_ (.A(net95),
    .B(_04036_),
    .Y(_04037_));
 sky130_fd_sc_hd__o22a_1 _10959_ (.A1(net55),
    .A2(net28),
    .B1(net26),
    .B2(net67),
    .X(_04038_));
 sky130_fd_sc_hd__xnor2_1 _10960_ (.A(net89),
    .B(_04038_),
    .Y(_04039_));
 sky130_fd_sc_hd__and2_1 _10961_ (.A(_04037_),
    .B(_04039_),
    .X(_04040_));
 sky130_fd_sc_hd__nor2_1 _10962_ (.A(_04037_),
    .B(_04039_),
    .Y(_04041_));
 sky130_fd_sc_hd__nor2_1 _10963_ (.A(_04040_),
    .B(_04041_),
    .Y(_04042_));
 sky130_fd_sc_hd__a22o_1 _10964_ (.A1(_06525_),
    .A2(net32),
    .B1(net30),
    .B2(_06559_),
    .X(_04043_));
 sky130_fd_sc_hd__xnor2_1 _10965_ (.A(net50),
    .B(_04043_),
    .Y(_04044_));
 sky130_fd_sc_hd__xor2_1 _10966_ (.A(_04042_),
    .B(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__and3_1 _10967_ (.A(_04034_),
    .B(_04035_),
    .C(_04045_),
    .X(_04046_));
 sky130_fd_sc_hd__a21oi_1 _10968_ (.A1(_04034_),
    .A2(_04035_),
    .B1(_04045_),
    .Y(_04047_));
 sky130_fd_sc_hd__o22a_1 _10969_ (.A1(net81),
    .A2(net10),
    .B1(net5),
    .B2(net77),
    .X(_04048_));
 sky130_fd_sc_hd__xnor2_1 _10970_ (.A(net19),
    .B(_04048_),
    .Y(_04049_));
 sky130_fd_sc_hd__nor2_1 _10971_ (.A(_03913_),
    .B(_04049_),
    .Y(_04050_));
 sky130_fd_sc_hd__and2_1 _10972_ (.A(_03913_),
    .B(_04049_),
    .X(_04051_));
 sky130_fd_sc_hd__nor2_1 _10973_ (.A(_04050_),
    .B(_04051_),
    .Y(_04052_));
 sky130_fd_sc_hd__nor2_1 _10974_ (.A(net73),
    .B(net20),
    .Y(_04053_));
 sky130_fd_sc_hd__xnor2_1 _10975_ (.A(_04052_),
    .B(_04053_),
    .Y(_04054_));
 sky130_fd_sc_hd__or3_1 _10976_ (.A(_04046_),
    .B(_04047_),
    .C(_04054_),
    .X(_04055_));
 sky130_fd_sc_hd__o21ai_1 _10977_ (.A1(_04046_),
    .A2(_04047_),
    .B1(_04054_),
    .Y(_04056_));
 sky130_fd_sc_hd__a21o_1 _10978_ (.A1(_03925_),
    .A2(_03927_),
    .B1(_03923_),
    .X(_04057_));
 sky130_fd_sc_hd__a21oi_1 _10979_ (.A1(_03933_),
    .A2(_03937_),
    .B1(_03943_),
    .Y(_04058_));
 sky130_fd_sc_hd__and3_1 _10980_ (.A(_03933_),
    .B(_03937_),
    .C(_03943_),
    .X(_04059_));
 sky130_fd_sc_hd__or2_1 _10981_ (.A(_04058_),
    .B(_04059_),
    .X(_04060_));
 sky130_fd_sc_hd__and2b_1 _10982_ (.A_N(_04060_),
    .B(_04057_),
    .X(_04061_));
 sky130_fd_sc_hd__xnor2_1 _10983_ (.A(_04057_),
    .B(_04060_),
    .Y(_04062_));
 sky130_fd_sc_hd__and3_1 _10984_ (.A(_04055_),
    .B(_04056_),
    .C(_04062_),
    .X(_04063_));
 sky130_fd_sc_hd__a21oi_1 _10985_ (.A1(_04055_),
    .A2(_04056_),
    .B1(_04062_),
    .Y(_04064_));
 sky130_fd_sc_hd__nor2_1 _10986_ (.A(_04063_),
    .B(_04064_),
    .Y(_04065_));
 sky130_fd_sc_hd__a21o_1 _10987_ (.A1(_03918_),
    .A2(_03958_),
    .B1(_03956_),
    .X(_04066_));
 sky130_fd_sc_hd__a21o_1 _10988_ (.A1(_03961_),
    .A2(_03965_),
    .B1(_03964_),
    .X(_04067_));
 sky130_fd_sc_hd__a21bo_1 _10989_ (.A1(_03907_),
    .A2(_03915_),
    .B1_N(_03917_),
    .X(_04068_));
 sky130_fd_sc_hd__nand2_1 _10990_ (.A(_03945_),
    .B(_03947_),
    .Y(_04069_));
 sky130_fd_sc_hd__o31a_1 _10991_ (.A1(net120),
    .A2(net19),
    .A3(_03950_),
    .B1(_03953_),
    .X(_04070_));
 sky130_fd_sc_hd__a21o_1 _10992_ (.A1(_03945_),
    .A2(_03947_),
    .B1(_04070_),
    .X(_04071_));
 sky130_fd_sc_hd__xor2_1 _10993_ (.A(_04069_),
    .B(_04070_),
    .X(_04072_));
 sky130_fd_sc_hd__nand2b_1 _10994_ (.A_N(_04072_),
    .B(_04068_),
    .Y(_04073_));
 sky130_fd_sc_hd__xnor2_1 _10995_ (.A(_04068_),
    .B(_04072_),
    .Y(_04074_));
 sky130_fd_sc_hd__nand2_1 _10996_ (.A(_04067_),
    .B(_04074_),
    .Y(_04075_));
 sky130_fd_sc_hd__xor2_1 _10997_ (.A(_04067_),
    .B(_04074_),
    .X(_04076_));
 sky130_fd_sc_hd__xor2_1 _10998_ (.A(_04066_),
    .B(_04076_),
    .X(_04077_));
 sky130_fd_sc_hd__nand2_1 _10999_ (.A(_04065_),
    .B(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__or2_1 _11000_ (.A(_04065_),
    .B(_04077_),
    .X(_04079_));
 sky130_fd_sc_hd__nand2_1 _11001_ (.A(_04078_),
    .B(_04079_),
    .Y(_04080_));
 sky130_fd_sc_hd__o21a_1 _11002_ (.A1(_03966_),
    .A2(_03967_),
    .B1(_03969_),
    .X(_04081_));
 sky130_fd_sc_hd__or2_1 _11003_ (.A(_04080_),
    .B(_04081_),
    .X(_04082_));
 sky130_fd_sc_hd__xnor2_1 _11004_ (.A(_04080_),
    .B(_04081_),
    .Y(_04083_));
 sky130_fd_sc_hd__a21oi_1 _11005_ (.A1(_03971_),
    .A2(_03973_),
    .B1(_04083_),
    .Y(_04084_));
 sky130_fd_sc_hd__and3_1 _11006_ (.A(_03971_),
    .B(_03973_),
    .C(_04083_),
    .X(_04085_));
 sky130_fd_sc_hd__or2_4 _11007_ (.A(_04084_),
    .B(_04085_),
    .X(_04086_));
 sky130_fd_sc_hd__nor2_1 _11008_ (.A(_03859_),
    .B(_03978_),
    .Y(_04087_));
 sky130_fd_sc_hd__nand2_1 _11009_ (.A(_03860_),
    .B(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__a21oi_2 _11010_ (.A1(_03857_),
    .A2(_03976_),
    .B1(_03977_),
    .Y(_04089_));
 sky130_fd_sc_hd__a21o_1 _11011_ (.A1(_03862_),
    .A2(_04087_),
    .B1(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__a31oi_1 _11012_ (.A1(_03629_),
    .A2(_03860_),
    .A3(_04087_),
    .B1(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__o31a_2 _11013_ (.A1(_03092_),
    .A2(_03625_),
    .A3(_04088_),
    .B1(_04091_),
    .X(_04092_));
 sky130_fd_sc_hd__xor2_4 _11014_ (.A(_04086_),
    .B(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__o21ai_1 _11015_ (.A1(_04016_),
    .A2(_04093_),
    .B1(net200),
    .Y(_04094_));
 sky130_fd_sc_hd__a21oi_1 _11016_ (.A1(_04016_),
    .A2(_04093_),
    .B1(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__a21o_1 _11017_ (.A1(net161),
    .A2(_01836_),
    .B1(_01837_),
    .X(_04096_));
 sky130_fd_sc_hd__a31oi_1 _11018_ (.A1(net161),
    .A2(_01836_),
    .A3(_01837_),
    .B1(_02324_),
    .Y(_04097_));
 sky130_fd_sc_hd__o21ba_1 _11019_ (.A1(_06169_),
    .A2(_03989_),
    .B1_N(_06157_),
    .X(_04098_));
 sky130_fd_sc_hd__mux2_1 _11020_ (.A0(_06390_),
    .A1(_04098_),
    .S(net284),
    .X(_04099_));
 sky130_fd_sc_hd__or2_1 _11021_ (.A(_06139_),
    .B(_04099_),
    .X(_04100_));
 sky130_fd_sc_hd__nand2_1 _11022_ (.A(_06139_),
    .B(_04099_),
    .Y(_04101_));
 sky130_fd_sc_hd__nand2_1 _11023_ (.A(reg1_val[13]),
    .B(curr_PC[13]),
    .Y(_04102_));
 sky130_fd_sc_hd__or2_1 _11024_ (.A(reg1_val[13]),
    .B(curr_PC[13]),
    .X(_04103_));
 sky130_fd_sc_hd__nand2_1 _11025_ (.A(_04102_),
    .B(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__a21oi_1 _11026_ (.A1(reg1_val[12]),
    .A2(curr_PC[12]),
    .B1(_03997_),
    .Y(_04105_));
 sky130_fd_sc_hd__xor2_1 _11027_ (.A(_04104_),
    .B(_04105_),
    .X(_04106_));
 sky130_fd_sc_hd__mux2_1 _11028_ (.A0(_03106_),
    .A1(_03110_),
    .S(net223),
    .X(_04107_));
 sky130_fd_sc_hd__mux2_1 _11029_ (.A0(_02650_),
    .A1(_04107_),
    .S(net225),
    .X(_04108_));
 sky130_fd_sc_hd__nand2_1 _11030_ (.A(_06331_),
    .B(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__o211a_1 _11031_ (.A1(_06331_),
    .A2(_04106_),
    .B1(_04109_),
    .C1(net210),
    .X(_04110_));
 sky130_fd_sc_hd__or2_1 _11032_ (.A(\div_res[12] ),
    .B(_04001_),
    .X(_04111_));
 sky130_fd_sc_hd__a21oi_1 _11033_ (.A1(net164),
    .A2(_04111_),
    .B1(\div_res[13] ),
    .Y(_04112_));
 sky130_fd_sc_hd__a31o_1 _11034_ (.A1(\div_res[13] ),
    .A2(net164),
    .A3(_04111_),
    .B1(net194),
    .X(_04113_));
 sky130_fd_sc_hd__or2_1 _11035_ (.A(\div_shifter[44] ),
    .B(_04004_),
    .X(_04114_));
 sky130_fd_sc_hd__a21oi_1 _11036_ (.A1(net232),
    .A2(_04114_),
    .B1(\div_shifter[45] ),
    .Y(_04115_));
 sky130_fd_sc_hd__a31o_1 _11037_ (.A1(\div_shifter[45] ),
    .A2(net232),
    .A3(_04114_),
    .B1(net192),
    .X(_04116_));
 sky130_fd_sc_hd__nand2_1 _11038_ (.A(_06121_),
    .B(net241),
    .Y(_04117_));
 sky130_fd_sc_hd__mux2_1 _11039_ (.A0(net197),
    .A1(net196),
    .S(_06127_),
    .X(_04118_));
 sky130_fd_sc_hd__a21o_1 _11040_ (.A1(net198),
    .A2(_04118_),
    .B1(_06133_),
    .X(_04119_));
 sky130_fd_sc_hd__o211a_1 _11041_ (.A1(_04115_),
    .A2(_04116_),
    .B1(_04117_),
    .C1(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__o21ai_2 _11042_ (.A1(net226),
    .A2(_02665_),
    .B1(_02335_),
    .Y(_04121_));
 sky130_fd_sc_hd__o221a_1 _11043_ (.A1(_04112_),
    .A2(_04113_),
    .B1(_04121_),
    .B2(net177),
    .C1(_04120_),
    .X(_04122_));
 sky130_fd_sc_hd__o21ai_1 _11044_ (.A1(_02314_),
    .A2(_04108_),
    .B1(_04122_),
    .Y(_04123_));
 sky130_fd_sc_hd__a311o_1 _11045_ (.A1(_02317_),
    .A2(_04100_),
    .A3(_04101_),
    .B1(_04110_),
    .C1(_04123_),
    .X(_04124_));
 sky130_fd_sc_hd__a211o_1 _11046_ (.A1(_04096_),
    .A2(_04097_),
    .B1(_04124_),
    .C1(_04095_),
    .X(_04125_));
 sky130_fd_sc_hd__or2_1 _11047_ (.A(curr_PC[13]),
    .B(_04014_),
    .X(_04126_));
 sky130_fd_sc_hd__a21oi_1 _11048_ (.A1(curr_PC[13]),
    .A2(_04014_),
    .B1(net242),
    .Y(_04127_));
 sky130_fd_sc_hd__a22o_4 _11049_ (.A1(net242),
    .A2(_04125_),
    .B1(_04126_),
    .B2(_04127_),
    .X(dest_val[13]));
 sky130_fd_sc_hd__or4_2 _11050_ (.A(_03746_),
    .B(_03865_),
    .C(_03984_),
    .D(_04093_),
    .X(_04128_));
 sky130_fd_sc_hd__nor2_1 _11051_ (.A(_03663_),
    .B(_04128_),
    .Y(_04129_));
 sky130_fd_sc_hd__or2_1 _11052_ (.A(net158),
    .B(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__a21bo_1 _11053_ (.A1(_04066_),
    .A2(_04076_),
    .B1_N(_04075_),
    .X(_04131_));
 sky130_fd_sc_hd__a21o_1 _11054_ (.A1(_04042_),
    .A2(_04044_),
    .B1(_04040_),
    .X(_04132_));
 sky130_fd_sc_hd__nand2_1 _11055_ (.A(_04021_),
    .B(_04025_),
    .Y(_04133_));
 sky130_fd_sc_hd__a21oi_4 _11056_ (.A1(net137),
    .A2(_04028_),
    .B1(_04032_),
    .Y(_04134_));
 sky130_fd_sc_hd__a21o_1 _11057_ (.A1(_04021_),
    .A2(_04025_),
    .B1(_04134_),
    .X(_04135_));
 sky130_fd_sc_hd__xor2_2 _11058_ (.A(_04133_),
    .B(_04134_),
    .X(_04136_));
 sky130_fd_sc_hd__nand2b_1 _11059_ (.A_N(_04136_),
    .B(_04132_),
    .Y(_04137_));
 sky130_fd_sc_hd__xnor2_2 _11060_ (.A(_04132_),
    .B(_04136_),
    .Y(_04138_));
 sky130_fd_sc_hd__o22a_1 _11061_ (.A1(net60),
    .A2(net47),
    .B1(net45),
    .B2(net58),
    .X(_04139_));
 sky130_fd_sc_hd__xnor2_1 _11062_ (.A(net96),
    .B(_04139_),
    .Y(_04140_));
 sky130_fd_sc_hd__o22a_1 _11063_ (.A1(net55),
    .A2(net26),
    .B1(net17),
    .B2(net28),
    .X(_04141_));
 sky130_fd_sc_hd__xnor2_1 _11064_ (.A(net89),
    .B(_04141_),
    .Y(_04142_));
 sky130_fd_sc_hd__nand2_1 _11065_ (.A(_04140_),
    .B(_04142_),
    .Y(_04143_));
 sky130_fd_sc_hd__or2_1 _11066_ (.A(_04140_),
    .B(_04142_),
    .X(_04144_));
 sky130_fd_sc_hd__and2_1 _11067_ (.A(_04143_),
    .B(_04144_),
    .X(_04145_));
 sky130_fd_sc_hd__a22o_1 _11068_ (.A1(_06517_),
    .A2(net32),
    .B1(net30),
    .B2(_06525_),
    .X(_04146_));
 sky130_fd_sc_hd__xnor2_2 _11069_ (.A(net50),
    .B(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__xor2_2 _11070_ (.A(_04145_),
    .B(_04147_),
    .X(_04148_));
 sky130_fd_sc_hd__a22o_1 _11071_ (.A1(_06540_),
    .A2(net40),
    .B1(net38),
    .B2(_06547_),
    .X(_04149_));
 sky130_fd_sc_hd__xor2_1 _11072_ (.A(net90),
    .B(_04149_),
    .X(_04150_));
 sky130_fd_sc_hd__a22o_1 _11073_ (.A1(_00163_),
    .A2(net44),
    .B1(net41),
    .B2(_00172_),
    .X(_04151_));
 sky130_fd_sc_hd__xor2_2 _11074_ (.A(net93),
    .B(_04151_),
    .X(_04152_));
 sky130_fd_sc_hd__nand2_1 _11075_ (.A(_04150_),
    .B(_04152_),
    .Y(_04153_));
 sky130_fd_sc_hd__or2_1 _11076_ (.A(_04150_),
    .B(_04152_),
    .X(_04154_));
 sky130_fd_sc_hd__and2_1 _11077_ (.A(_04153_),
    .B(_04154_),
    .X(_04155_));
 sky130_fd_sc_hd__o22a_1 _11078_ (.A1(net34),
    .A2(net14),
    .B1(net12),
    .B2(net36),
    .X(_04156_));
 sky130_fd_sc_hd__xnor2_1 _11079_ (.A(net126),
    .B(_04156_),
    .Y(_04157_));
 sky130_fd_sc_hd__or2_1 _11080_ (.A(_00359_),
    .B(net7),
    .X(_04158_));
 sky130_fd_sc_hd__nor2_1 _11081_ (.A(_00358_),
    .B(net7),
    .Y(_04159_));
 sky130_fd_sc_hd__mux2_1 _11082_ (.A0(_04158_),
    .A1(_04159_),
    .S(net122),
    .X(_04160_));
 sky130_fd_sc_hd__nor2_1 _11083_ (.A(_04157_),
    .B(_04160_),
    .Y(_04161_));
 sky130_fd_sc_hd__and2_1 _11084_ (.A(_04157_),
    .B(_04160_),
    .X(_04162_));
 sky130_fd_sc_hd__nor2_1 _11085_ (.A(_04161_),
    .B(_04162_),
    .Y(_04163_));
 sky130_fd_sc_hd__and2b_1 _11086_ (.A_N(_04163_),
    .B(_04155_),
    .X(_04164_));
 sky130_fd_sc_hd__xnor2_1 _11087_ (.A(_04155_),
    .B(_04163_),
    .Y(_04165_));
 sky130_fd_sc_hd__xnor2_1 _11088_ (.A(_04148_),
    .B(_04165_),
    .Y(_04166_));
 sky130_fd_sc_hd__o22a_1 _11089_ (.A1(net85),
    .A2(net10),
    .B1(net5),
    .B2(net81),
    .X(_04167_));
 sky130_fd_sc_hd__xnor2_1 _11090_ (.A(net20),
    .B(_04167_),
    .Y(_04168_));
 sky130_fd_sc_hd__o22a_1 _11091_ (.A1(net101),
    .A2(net24),
    .B1(net16),
    .B2(net99),
    .X(_04169_));
 sky130_fd_sc_hd__xnor2_1 _11092_ (.A(net69),
    .B(_04169_),
    .Y(_04170_));
 sky130_fd_sc_hd__nor2_1 _11093_ (.A(net77),
    .B(net19),
    .Y(_04171_));
 sky130_fd_sc_hd__xnor2_1 _11094_ (.A(_04170_),
    .B(_04171_),
    .Y(_04172_));
 sky130_fd_sc_hd__nand2b_1 _11095_ (.A_N(_04168_),
    .B(_04172_),
    .Y(_04173_));
 sky130_fd_sc_hd__xor2_1 _11096_ (.A(_04168_),
    .B(_04172_),
    .X(_04174_));
 sky130_fd_sc_hd__nor2_1 _11097_ (.A(_04166_),
    .B(_04174_),
    .Y(_04175_));
 sky130_fd_sc_hd__nand2_1 _11098_ (.A(_04166_),
    .B(_04174_),
    .Y(_04176_));
 sky130_fd_sc_hd__and2b_1 _11099_ (.A_N(_04175_),
    .B(_04176_),
    .X(_04177_));
 sky130_fd_sc_hd__xor2_2 _11100_ (.A(_04138_),
    .B(_04177_),
    .X(_04178_));
 sky130_fd_sc_hd__a21bo_1 _11101_ (.A1(_04056_),
    .A2(_04062_),
    .B1_N(_04055_),
    .X(_04179_));
 sky130_fd_sc_hd__or2_1 _11102_ (.A(_04058_),
    .B(_04061_),
    .X(_04180_));
 sky130_fd_sc_hd__a21o_1 _11103_ (.A1(_04026_),
    .A2(_04033_),
    .B1(_04046_),
    .X(_04181_));
 sky130_fd_sc_hd__a21o_1 _11104_ (.A1(_04052_),
    .A2(_04053_),
    .B1(_04050_),
    .X(_04182_));
 sky130_fd_sc_hd__nand2_1 _11105_ (.A(_04181_),
    .B(_04182_),
    .Y(_04183_));
 sky130_fd_sc_hd__xor2_2 _11106_ (.A(_04181_),
    .B(_04182_),
    .X(_04184_));
 sky130_fd_sc_hd__xnor2_2 _11107_ (.A(_04180_),
    .B(_04184_),
    .Y(_04185_));
 sky130_fd_sc_hd__and2_1 _11108_ (.A(_04071_),
    .B(_04073_),
    .X(_04186_));
 sky130_fd_sc_hd__xnor2_1 _11109_ (.A(_04185_),
    .B(_04186_),
    .Y(_04187_));
 sky130_fd_sc_hd__nand2b_1 _11110_ (.A_N(_04187_),
    .B(_04179_),
    .Y(_04188_));
 sky130_fd_sc_hd__xnor2_1 _11111_ (.A(_04179_),
    .B(_04187_),
    .Y(_04189_));
 sky130_fd_sc_hd__nand2_1 _11112_ (.A(_04178_),
    .B(_04189_),
    .Y(_04190_));
 sky130_fd_sc_hd__xnor2_1 _11113_ (.A(_04178_),
    .B(_04189_),
    .Y(_04191_));
 sky130_fd_sc_hd__nand2b_1 _11114_ (.A_N(_04191_),
    .B(_04131_),
    .Y(_04192_));
 sky130_fd_sc_hd__xor2_1 _11115_ (.A(_04131_),
    .B(_04191_),
    .X(_04193_));
 sky130_fd_sc_hd__a21oi_1 _11116_ (.A1(_04078_),
    .A2(_04082_),
    .B1(_04193_),
    .Y(_04194_));
 sky130_fd_sc_hd__and3_1 _11117_ (.A(_04078_),
    .B(_04082_),
    .C(_04193_),
    .X(_04195_));
 sky130_fd_sc_hd__or2_2 _11118_ (.A(_04194_),
    .B(_04195_),
    .X(_04196_));
 sky130_fd_sc_hd__o21ba_1 _11119_ (.A1(_03975_),
    .A2(_04084_),
    .B1_N(_04085_),
    .X(_04197_));
 sky130_fd_sc_hd__nor2_1 _11120_ (.A(_03978_),
    .B(_04086_),
    .Y(_04198_));
 sky130_fd_sc_hd__a21o_1 _11121_ (.A1(_03979_),
    .A2(_04198_),
    .B1(_04197_),
    .X(_04199_));
 sky130_fd_sc_hd__and2_1 _11122_ (.A(_03980_),
    .B(_04198_),
    .X(_04200_));
 sky130_fd_sc_hd__a21oi_4 _11123_ (.A1(net3),
    .A2(_04200_),
    .B1(_04199_),
    .Y(_04201_));
 sky130_fd_sc_hd__xnor2_4 _11124_ (.A(_04196_),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__a21oi_1 _11125_ (.A1(_04130_),
    .A2(_04202_),
    .B1(_02242_),
    .Y(_04203_));
 sky130_fd_sc_hd__o21a_1 _11126_ (.A1(_04130_),
    .A2(_04202_),
    .B1(_04203_),
    .X(_04204_));
 sky130_fd_sc_hd__a211o_1 _11127_ (.A1(net161),
    .A2(_01838_),
    .B1(_01840_),
    .C1(_01841_),
    .X(_04205_));
 sky130_fd_sc_hd__or3b_1 _11128_ (.A(net157),
    .B(_01842_),
    .C_N(_01838_),
    .X(_04206_));
 sky130_fd_sc_hd__o21bai_1 _11129_ (.A1(_06139_),
    .A2(_04098_),
    .B1_N(_06127_),
    .Y(_04207_));
 sky130_fd_sc_hd__mux2_1 _11130_ (.A0(_06392_),
    .A1(_04207_),
    .S(net284),
    .X(_04208_));
 sky130_fd_sc_hd__nand2_1 _11131_ (.A(_06109_),
    .B(_04208_),
    .Y(_04209_));
 sky130_fd_sc_hd__o211a_1 _11132_ (.A1(_06109_),
    .A2(_04208_),
    .B1(_04209_),
    .C1(_02317_),
    .X(_04210_));
 sky130_fd_sc_hd__nand2_1 _11133_ (.A(net291),
    .B(curr_PC[14]),
    .Y(_04211_));
 sky130_fd_sc_hd__or2_1 _11134_ (.A(net291),
    .B(curr_PC[14]),
    .X(_04212_));
 sky130_fd_sc_hd__nand2_1 _11135_ (.A(_04211_),
    .B(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__o21a_1 _11136_ (.A1(_04104_),
    .A2(_04105_),
    .B1(_04102_),
    .X(_04214_));
 sky130_fd_sc_hd__xor2_1 _11137_ (.A(_04213_),
    .B(_04214_),
    .X(_04215_));
 sky130_fd_sc_hd__or2_1 _11138_ (.A(net224),
    .B(_03249_),
    .X(_04216_));
 sky130_fd_sc_hd__o211a_1 _11139_ (.A1(net222),
    .A2(_03247_),
    .B1(_04216_),
    .C1(net225),
    .X(_04217_));
 sky130_fd_sc_hd__a21oi_2 _11140_ (.A1(net227),
    .A2(_02528_),
    .B1(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__nand2_1 _11141_ (.A(net229),
    .B(_04218_),
    .Y(_04219_));
 sky130_fd_sc_hd__o211a_1 _11142_ (.A1(net229),
    .A2(_04215_),
    .B1(_04219_),
    .C1(net210),
    .X(_04220_));
 sky130_fd_sc_hd__or2_1 _11143_ (.A(\div_shifter[45] ),
    .B(_04114_),
    .X(_04221_));
 sky130_fd_sc_hd__a21oi_1 _11144_ (.A1(net234),
    .A2(_04221_),
    .B1(\div_shifter[46] ),
    .Y(_04222_));
 sky130_fd_sc_hd__a31o_1 _11145_ (.A1(\div_shifter[46] ),
    .A2(net234),
    .A3(_04221_),
    .B1(net192),
    .X(_04223_));
 sky130_fd_sc_hd__or2_1 _11146_ (.A(_04222_),
    .B(_04223_),
    .X(_04224_));
 sky130_fd_sc_hd__or2_1 _11147_ (.A(\div_res[13] ),
    .B(_04111_),
    .X(_04225_));
 sky130_fd_sc_hd__a21oi_1 _11148_ (.A1(net164),
    .A2(_04225_),
    .B1(\div_res[14] ),
    .Y(_04226_));
 sky130_fd_sc_hd__a31o_1 _11149_ (.A1(\div_res[14] ),
    .A2(net164),
    .A3(_04225_),
    .B1(net194),
    .X(_04227_));
 sky130_fd_sc_hd__mux2_1 _11150_ (.A0(net197),
    .A1(net196),
    .S(_06103_),
    .X(_04228_));
 sky130_fd_sc_hd__a21oi_1 _11151_ (.A1(net198),
    .A2(_04228_),
    .B1(_06097_),
    .Y(_04229_));
 sky130_fd_sc_hd__a21oi_1 _11152_ (.A1(_06086_),
    .A2(net241),
    .B1(_04229_),
    .Y(_04230_));
 sky130_fd_sc_hd__o211a_1 _11153_ (.A1(_04226_),
    .A2(_04227_),
    .B1(_04230_),
    .C1(_04224_),
    .X(_04231_));
 sky130_fd_sc_hd__o21a_1 _11154_ (.A1(net226),
    .A2(_02498_),
    .B1(_02335_),
    .X(_04232_));
 sky130_fd_sc_hd__inv_2 _11155_ (.A(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__o221a_1 _11156_ (.A1(_02314_),
    .A2(_04218_),
    .B1(_04233_),
    .B2(net177),
    .C1(_04231_),
    .X(_04234_));
 sky130_fd_sc_hd__or3b_1 _11157_ (.A(_04210_),
    .B(_04220_),
    .C_N(_04234_),
    .X(_04235_));
 sky130_fd_sc_hd__a311o_1 _11158_ (.A1(_02323_),
    .A2(_04205_),
    .A3(_04206_),
    .B1(_04235_),
    .C1(_04204_),
    .X(_04236_));
 sky130_fd_sc_hd__and3_1 _11159_ (.A(curr_PC[13]),
    .B(curr_PC[14]),
    .C(_04014_),
    .X(_04237_));
 sky130_fd_sc_hd__a21oi_1 _11160_ (.A1(curr_PC[13]),
    .A2(_04014_),
    .B1(curr_PC[14]),
    .Y(_04238_));
 sky130_fd_sc_hd__nor2_1 _11161_ (.A(_04237_),
    .B(_04238_),
    .Y(_04239_));
 sky130_fd_sc_hd__mux2_8 _11162_ (.A0(_04236_),
    .A1(_04239_),
    .S(net248),
    .X(dest_val[14]));
 sky130_fd_sc_hd__a21oi_1 _11163_ (.A1(_04129_),
    .A2(_04202_),
    .B1(net158),
    .Y(_04240_));
 sky130_fd_sc_hd__o22a_1 _11164_ (.A1(net99),
    .A2(net10),
    .B1(net5),
    .B2(net85),
    .X(_04241_));
 sky130_fd_sc_hd__xnor2_1 _11165_ (.A(net19),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__a22o_1 _11166_ (.A1(_06547_),
    .A2(net43),
    .B1(net41),
    .B2(_00163_),
    .X(_04243_));
 sky130_fd_sc_hd__xor2_1 _11167_ (.A(net93),
    .B(_04243_),
    .X(_04244_));
 sky130_fd_sc_hd__nand2b_1 _11168_ (.A_N(_04242_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__nand2b_1 _11169_ (.A_N(_04244_),
    .B(_04242_),
    .Y(_04246_));
 sky130_fd_sc_hd__nand2_1 _11170_ (.A(_04245_),
    .B(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__o22a_1 _11171_ (.A1(net52),
    .A2(net23),
    .B1(net16),
    .B2(net101),
    .X(_04248_));
 sky130_fd_sc_hd__xnor2_1 _11172_ (.A(net69),
    .B(_04248_),
    .Y(_04249_));
 sky130_fd_sc_hd__or2_1 _11173_ (.A(_04247_),
    .B(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__nand2_1 _11174_ (.A(_04247_),
    .B(_04249_),
    .Y(_04251_));
 sky130_fd_sc_hd__nand2_1 _11175_ (.A(_04250_),
    .B(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__o22a_1 _11176_ (.A1(net26),
    .A2(net17),
    .B1(net14),
    .B2(net28),
    .X(_04253_));
 sky130_fd_sc_hd__xnor2_1 _11177_ (.A(net89),
    .B(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__and2_1 _11178_ (.A(net122),
    .B(_04254_),
    .X(_04255_));
 sky130_fd_sc_hd__nor2_1 _11179_ (.A(net122),
    .B(_04254_),
    .Y(_04256_));
 sky130_fd_sc_hd__nor2_1 _11180_ (.A(_04255_),
    .B(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__o22a_1 _11181_ (.A1(net34),
    .A2(net12),
    .B1(net7),
    .B2(net36),
    .X(_04258_));
 sky130_fd_sc_hd__xnor2_2 _11182_ (.A(net126),
    .B(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__xor2_2 _11183_ (.A(_04257_),
    .B(_04259_),
    .X(_04260_));
 sky130_fd_sc_hd__a22o_1 _11184_ (.A1(_06563_),
    .A2(net40),
    .B1(net38),
    .B2(_06540_),
    .X(_04261_));
 sky130_fd_sc_hd__xor2_1 _11185_ (.A(net90),
    .B(_04261_),
    .X(_04262_));
 sky130_fd_sc_hd__a22o_1 _11186_ (.A1(_00143_),
    .A2(net32),
    .B1(net30),
    .B2(_06517_),
    .X(_04263_));
 sky130_fd_sc_hd__xnor2_1 _11187_ (.A(net50),
    .B(_04263_),
    .Y(_04264_));
 sky130_fd_sc_hd__and2_1 _11188_ (.A(_04262_),
    .B(_04264_),
    .X(_04265_));
 sky130_fd_sc_hd__nor2_1 _11189_ (.A(_04262_),
    .B(_04264_),
    .Y(_04266_));
 sky130_fd_sc_hd__nor2_1 _11190_ (.A(_04265_),
    .B(_04266_),
    .Y(_04267_));
 sky130_fd_sc_hd__o22a_1 _11191_ (.A1(net66),
    .A2(net47),
    .B1(net45),
    .B2(net60),
    .X(_04268_));
 sky130_fd_sc_hd__xnor2_2 _11192_ (.A(net96),
    .B(_04268_),
    .Y(_04269_));
 sky130_fd_sc_hd__xor2_2 _11193_ (.A(_04267_),
    .B(_04269_),
    .X(_04270_));
 sky130_fd_sc_hd__xnor2_2 _11194_ (.A(_04153_),
    .B(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__xnor2_2 _11195_ (.A(_04260_),
    .B(_04271_),
    .Y(_04272_));
 sky130_fd_sc_hd__xnor2_2 _11196_ (.A(_04252_),
    .B(_04272_),
    .Y(_04273_));
 sky130_fd_sc_hd__a21bo_1 _11197_ (.A1(_04145_),
    .A2(_04147_),
    .B1_N(_04143_),
    .X(_04274_));
 sky130_fd_sc_hd__nor2_1 _11198_ (.A(net81),
    .B(net19),
    .Y(_04275_));
 sky130_fd_sc_hd__xnor2_1 _11199_ (.A(_04274_),
    .B(_04275_),
    .Y(_04276_));
 sky130_fd_sc_hd__or2_1 _11200_ (.A(_04161_),
    .B(_04276_),
    .X(_04277_));
 sky130_fd_sc_hd__nand2_1 _11201_ (.A(_04161_),
    .B(_04276_),
    .Y(_04278_));
 sky130_fd_sc_hd__and2_1 _11202_ (.A(_04277_),
    .B(_04278_),
    .X(_04279_));
 sky130_fd_sc_hd__nand2b_1 _11203_ (.A_N(_04273_),
    .B(_04279_),
    .Y(_04280_));
 sky130_fd_sc_hd__xnor2_2 _11204_ (.A(_04273_),
    .B(_04279_),
    .Y(_04281_));
 sky130_fd_sc_hd__a21o_1 _11205_ (.A1(_04138_),
    .A2(_04176_),
    .B1(_04175_),
    .X(_04282_));
 sky130_fd_sc_hd__a21bo_1 _11206_ (.A1(_04180_),
    .A2(_04184_),
    .B1_N(_04183_),
    .X(_04283_));
 sky130_fd_sc_hd__nand2_2 _11207_ (.A(_04135_),
    .B(_04137_),
    .Y(_04284_));
 sky130_fd_sc_hd__a21o_1 _11208_ (.A1(_04148_),
    .A2(_04165_),
    .B1(_04164_),
    .X(_04285_));
 sky130_fd_sc_hd__o31a_1 _11209_ (.A1(net77),
    .A2(net19),
    .A3(_04170_),
    .B1(_04173_),
    .X(_04286_));
 sky130_fd_sc_hd__inv_2 _11210_ (.A(_04286_),
    .Y(_04287_));
 sky130_fd_sc_hd__and2_1 _11211_ (.A(_04285_),
    .B(_04287_),
    .X(_04288_));
 sky130_fd_sc_hd__xnor2_2 _11212_ (.A(_04285_),
    .B(_04287_),
    .Y(_04289_));
 sky130_fd_sc_hd__inv_2 _11213_ (.A(_04289_),
    .Y(_04290_));
 sky130_fd_sc_hd__xnor2_2 _11214_ (.A(_04284_),
    .B(_04289_),
    .Y(_04291_));
 sky130_fd_sc_hd__xnor2_2 _11215_ (.A(_04283_),
    .B(_04291_),
    .Y(_04292_));
 sky130_fd_sc_hd__nand2b_1 _11216_ (.A_N(_04292_),
    .B(_04282_),
    .Y(_04293_));
 sky130_fd_sc_hd__xnor2_2 _11217_ (.A(_04282_),
    .B(_04292_),
    .Y(_04294_));
 sky130_fd_sc_hd__nand2_1 _11218_ (.A(_04281_),
    .B(_04294_),
    .Y(_04295_));
 sky130_fd_sc_hd__xnor2_2 _11219_ (.A(_04281_),
    .B(_04294_),
    .Y(_04296_));
 sky130_fd_sc_hd__o21ai_2 _11220_ (.A1(_04185_),
    .A2(_04186_),
    .B1(_04188_),
    .Y(_04297_));
 sky130_fd_sc_hd__nand2b_1 _11221_ (.A_N(_04296_),
    .B(_04297_),
    .Y(_04298_));
 sky130_fd_sc_hd__xor2_2 _11222_ (.A(_04296_),
    .B(_04297_),
    .X(_04299_));
 sky130_fd_sc_hd__a21oi_1 _11223_ (.A1(_04190_),
    .A2(_04192_),
    .B1(_04299_),
    .Y(_04300_));
 sky130_fd_sc_hd__nand3_2 _11224_ (.A(_04190_),
    .B(_04192_),
    .C(_04299_),
    .Y(_04301_));
 sky130_fd_sc_hd__nand2b_4 _11225_ (.A_N(_04300_),
    .B(_04301_),
    .Y(_04302_));
 sky130_fd_sc_hd__o21ba_1 _11226_ (.A1(_04084_),
    .A2(_04194_),
    .B1_N(_04195_),
    .X(_04303_));
 sky130_fd_sc_hd__nor2_1 _11227_ (.A(_04086_),
    .B(_04196_),
    .Y(_04304_));
 sky130_fd_sc_hd__a21o_1 _11228_ (.A1(_04089_),
    .A2(_04304_),
    .B1(_04303_),
    .X(_04305_));
 sky130_fd_sc_hd__and2_1 _11229_ (.A(_04087_),
    .B(_04304_),
    .X(_04306_));
 sky130_fd_sc_hd__a21o_1 _11230_ (.A1(_03863_),
    .A2(_04306_),
    .B1(_04305_),
    .X(_04307_));
 sky130_fd_sc_hd__a31o_2 _11231_ (.A1(_03367_),
    .A2(_03861_),
    .A3(_04306_),
    .B1(_04307_),
    .X(_04308_));
 sky130_fd_sc_hd__xnor2_4 _11232_ (.A(_04302_),
    .B(_04308_),
    .Y(_04309_));
 sky130_fd_sc_hd__or2_1 _11233_ (.A(_04240_),
    .B(_04309_),
    .X(_04310_));
 sky130_fd_sc_hd__nand2_1 _11234_ (.A(_04240_),
    .B(_04309_),
    .Y(_04311_));
 sky130_fd_sc_hd__a21oi_1 _11235_ (.A1(net161),
    .A2(_01843_),
    .B1(_01845_),
    .Y(_04312_));
 sky130_fd_sc_hd__a311oi_1 _11236_ (.A1(net161),
    .A2(_01843_),
    .A3(_01845_),
    .B1(_02324_),
    .C1(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__a21o_1 _11237_ (.A1(_06109_),
    .A2(_04207_),
    .B1(_06103_),
    .X(_04314_));
 sky130_fd_sc_hd__mux2_1 _11238_ (.A0(_06394_),
    .A1(_04314_),
    .S(net284),
    .X(_04315_));
 sky130_fd_sc_hd__nand2_1 _11239_ (.A(_06064_),
    .B(_04315_),
    .Y(_04316_));
 sky130_fd_sc_hd__o211a_1 _11240_ (.A1(_06064_),
    .A2(_04315_),
    .B1(_04316_),
    .C1(_02317_),
    .X(_04317_));
 sky130_fd_sc_hd__and2_1 _11241_ (.A(net290),
    .B(curr_PC[15]),
    .X(_04318_));
 sky130_fd_sc_hd__nor2_1 _11242_ (.A(net290),
    .B(curr_PC[15]),
    .Y(_04319_));
 sky130_fd_sc_hd__nor2_1 _11243_ (.A(_04318_),
    .B(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__o21a_1 _11244_ (.A1(_04213_),
    .A2(_04214_),
    .B1(_04211_),
    .X(_04321_));
 sky130_fd_sc_hd__xnor2_1 _11245_ (.A(_04320_),
    .B(_04321_),
    .Y(_04322_));
 sky130_fd_sc_hd__mux2_1 _11246_ (.A0(_03380_),
    .A1(_03382_),
    .S(net222),
    .X(_04323_));
 sky130_fd_sc_hd__and3_1 _11247_ (.A(net226),
    .B(_02340_),
    .C(_02342_),
    .X(_04324_));
 sky130_fd_sc_hd__a21oi_2 _11248_ (.A1(net225),
    .A2(_04323_),
    .B1(_04324_),
    .Y(_04325_));
 sky130_fd_sc_hd__nand2_1 _11249_ (.A(net229),
    .B(_04325_),
    .Y(_04326_));
 sky130_fd_sc_hd__o211a_1 _11250_ (.A1(net229),
    .A2(_04322_),
    .B1(_04326_),
    .C1(_06475_),
    .X(_04327_));
 sky130_fd_sc_hd__or2_1 _11251_ (.A(\div_res[14] ),
    .B(_04225_),
    .X(_04328_));
 sky130_fd_sc_hd__and3_1 _11252_ (.A(\div_res[15] ),
    .B(net164),
    .C(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__a21oi_1 _11253_ (.A1(net164),
    .A2(_04328_),
    .B1(\div_res[15] ),
    .Y(_04330_));
 sky130_fd_sc_hd__or3_1 _11254_ (.A(net194),
    .B(_04329_),
    .C(_04330_),
    .X(_04331_));
 sky130_fd_sc_hd__or2_1 _11255_ (.A(\div_shifter[46] ),
    .B(_04221_),
    .X(_04332_));
 sky130_fd_sc_hd__a21oi_1 _11256_ (.A1(net232),
    .A2(_04332_),
    .B1(\div_shifter[47] ),
    .Y(_04333_));
 sky130_fd_sc_hd__a31o_1 _11257_ (.A1(\div_shifter[47] ),
    .A2(net232),
    .A3(_04332_),
    .B1(net192),
    .X(_04334_));
 sky130_fd_sc_hd__nor2_1 _11258_ (.A(_04333_),
    .B(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__mux2_1 _11259_ (.A0(net197),
    .A1(net196),
    .S(_06042_),
    .X(_04336_));
 sky130_fd_sc_hd__a21oi_1 _11260_ (.A1(net198),
    .A2(_04336_),
    .B1(_06053_),
    .Y(_04337_));
 sky130_fd_sc_hd__a211o_1 _11261_ (.A1(_06031_),
    .A2(net241),
    .B1(_04335_),
    .C1(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__o21a_1 _11262_ (.A1(net226),
    .A2(_02307_),
    .B1(_02335_),
    .X(_04339_));
 sky130_fd_sc_hd__a2bb2o_1 _11263_ (.A1_N(_02314_),
    .A2_N(_04325_),
    .B1(_04339_),
    .B2(net179),
    .X(_04340_));
 sky130_fd_sc_hd__or3b_1 _11264_ (.A(_04338_),
    .B(_04340_),
    .C_N(_04331_),
    .X(_04341_));
 sky130_fd_sc_hd__or3_1 _11265_ (.A(_04317_),
    .B(_04327_),
    .C(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__a311o_1 _11266_ (.A1(net200),
    .A2(_04310_),
    .A3(_04311_),
    .B1(_04313_),
    .C1(_04342_),
    .X(_04343_));
 sky130_fd_sc_hd__or2_1 _11267_ (.A(curr_PC[15]),
    .B(_04237_),
    .X(_04344_));
 sky130_fd_sc_hd__and2_1 _11268_ (.A(curr_PC[15]),
    .B(_04237_),
    .X(_04345_));
 sky130_fd_sc_hd__nor2_1 _11269_ (.A(net243),
    .B(_04345_),
    .Y(_04346_));
 sky130_fd_sc_hd__a22o_4 _11270_ (.A1(net243),
    .A2(_04343_),
    .B1(_04344_),
    .B2(_04346_),
    .X(dest_val[15]));
 sky130_fd_sc_hd__nor4b_4 _11271_ (.A(_03663_),
    .B(_04309_),
    .C(_04128_),
    .D_N(_04202_),
    .Y(_04347_));
 sky130_fd_sc_hd__or2_1 _11272_ (.A(net158),
    .B(_04347_),
    .X(_04348_));
 sky130_fd_sc_hd__a21oi_1 _11273_ (.A1(_04267_),
    .A2(_04269_),
    .B1(_04265_),
    .Y(_04349_));
 sky130_fd_sc_hd__o22a_1 _11274_ (.A1(net67),
    .A2(net47),
    .B1(net45),
    .B2(net66),
    .X(_04350_));
 sky130_fd_sc_hd__xnor2_1 _11275_ (.A(net95),
    .B(_04350_),
    .Y(_04351_));
 sky130_fd_sc_hd__a22oi_1 _11276_ (.A1(_00143_),
    .A2(net30),
    .B1(_00408_),
    .B2(net32),
    .Y(_04352_));
 sky130_fd_sc_hd__xnor2_1 _11277_ (.A(_00216_),
    .B(_04352_),
    .Y(_04353_));
 sky130_fd_sc_hd__nand2_1 _11278_ (.A(_04351_),
    .B(_04353_),
    .Y(_04354_));
 sky130_fd_sc_hd__or2_1 _11279_ (.A(_04351_),
    .B(_04353_),
    .X(_04355_));
 sky130_fd_sc_hd__nand2_1 _11280_ (.A(_04354_),
    .B(_04355_),
    .Y(_04356_));
 sky130_fd_sc_hd__nor2_1 _11281_ (.A(_04349_),
    .B(_04356_),
    .Y(_04357_));
 sky130_fd_sc_hd__xnor2_1 _11282_ (.A(_04349_),
    .B(_04356_),
    .Y(_04358_));
 sky130_fd_sc_hd__o22a_1 _11283_ (.A1(net26),
    .A2(net14),
    .B1(net12),
    .B2(net28),
    .X(_04359_));
 sky130_fd_sc_hd__xnor2_1 _11284_ (.A(_00301_),
    .B(_04359_),
    .Y(_04360_));
 sky130_fd_sc_hd__o21ai_1 _11285_ (.A1(_00282_),
    .A2(net8),
    .B1(net125),
    .Y(_04361_));
 sky130_fd_sc_hd__o21ai_2 _11286_ (.A1(_00292_),
    .A2(net8),
    .B1(_04361_),
    .Y(_04362_));
 sky130_fd_sc_hd__nor2_1 _11287_ (.A(_04360_),
    .B(_04362_),
    .Y(_04363_));
 sky130_fd_sc_hd__and2_1 _11288_ (.A(_04360_),
    .B(_04362_),
    .X(_04364_));
 sky130_fd_sc_hd__nor2_1 _11289_ (.A(_04363_),
    .B(_04364_),
    .Y(_04365_));
 sky130_fd_sc_hd__nor2_1 _11290_ (.A(_04358_),
    .B(_04365_),
    .Y(_04366_));
 sky130_fd_sc_hd__and2_1 _11291_ (.A(_04358_),
    .B(_04365_),
    .X(_04367_));
 sky130_fd_sc_hd__or2_1 _11292_ (.A(_04366_),
    .B(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__o22a_1 _11293_ (.A1(net54),
    .A2(net23),
    .B1(net15),
    .B2(net52),
    .X(_04369_));
 sky130_fd_sc_hd__xnor2_1 _11294_ (.A(net69),
    .B(_04369_),
    .Y(_04370_));
 sky130_fd_sc_hd__inv_2 _11295_ (.A(_04370_),
    .Y(_04371_));
 sky130_fd_sc_hd__a22o_1 _11296_ (.A1(_06559_),
    .A2(net40),
    .B1(net38),
    .B2(_06563_),
    .X(_04372_));
 sky130_fd_sc_hd__xor2_1 _11297_ (.A(_00245_),
    .B(_04372_),
    .X(_04373_));
 sky130_fd_sc_hd__xor2_1 _11298_ (.A(_04370_),
    .B(_04373_),
    .X(_04374_));
 sky130_fd_sc_hd__a22o_1 _11299_ (.A1(_06540_),
    .A2(net43),
    .B1(net42),
    .B2(_06547_),
    .X(_04375_));
 sky130_fd_sc_hd__xor2_1 _11300_ (.A(net93),
    .B(_04375_),
    .X(_04376_));
 sky130_fd_sc_hd__and2b_1 _11301_ (.A_N(_04374_),
    .B(_04376_),
    .X(_04377_));
 sky130_fd_sc_hd__and2b_1 _11302_ (.A_N(_04376_),
    .B(_04374_),
    .X(_04378_));
 sky130_fd_sc_hd__or2_1 _11303_ (.A(_04377_),
    .B(_04378_),
    .X(_04379_));
 sky130_fd_sc_hd__xnor2_2 _11304_ (.A(_04368_),
    .B(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__a21oi_2 _11305_ (.A1(_04257_),
    .A2(_04259_),
    .B1(_04255_),
    .Y(_04381_));
 sky130_fd_sc_hd__o22a_1 _11306_ (.A1(net101),
    .A2(net10),
    .B1(net5),
    .B2(net99),
    .X(_04382_));
 sky130_fd_sc_hd__xnor2_1 _11307_ (.A(net20),
    .B(_04382_),
    .Y(_04383_));
 sky130_fd_sc_hd__xnor2_1 _11308_ (.A(_04381_),
    .B(_04383_),
    .Y(_04384_));
 sky130_fd_sc_hd__or3_1 _11309_ (.A(net85),
    .B(net20),
    .C(_04384_),
    .X(_04385_));
 sky130_fd_sc_hd__o21ai_1 _11310_ (.A1(net85),
    .A2(net20),
    .B1(_04384_),
    .Y(_04386_));
 sky130_fd_sc_hd__and2_1 _11311_ (.A(_04385_),
    .B(_04386_),
    .X(_04387_));
 sky130_fd_sc_hd__and2b_1 _11312_ (.A_N(_04380_),
    .B(_04387_),
    .X(_04388_));
 sky130_fd_sc_hd__xnor2_2 _11313_ (.A(_04380_),
    .B(_04387_),
    .Y(_04389_));
 sky130_fd_sc_hd__o21ai_2 _11314_ (.A1(_04252_),
    .A2(_04272_),
    .B1(_04280_),
    .Y(_04390_));
 sky130_fd_sc_hd__a21bo_1 _11315_ (.A1(_04274_),
    .A2(_04275_),
    .B1_N(_04277_),
    .X(_04391_));
 sky130_fd_sc_hd__a32oi_2 _11316_ (.A1(_04150_),
    .A2(_04152_),
    .A3(_04270_),
    .B1(_04271_),
    .B2(_04260_),
    .Y(_04392_));
 sky130_fd_sc_hd__a21oi_1 _11317_ (.A1(_04245_),
    .A2(_04250_),
    .B1(_04392_),
    .Y(_04393_));
 sky130_fd_sc_hd__and3_1 _11318_ (.A(_04245_),
    .B(_04250_),
    .C(_04392_),
    .X(_04394_));
 sky130_fd_sc_hd__nor2_1 _11319_ (.A(_04393_),
    .B(_04394_),
    .Y(_04395_));
 sky130_fd_sc_hd__xnor2_2 _11320_ (.A(_04391_),
    .B(_04395_),
    .Y(_04396_));
 sky130_fd_sc_hd__a21oi_2 _11321_ (.A1(_04284_),
    .A2(_04290_),
    .B1(_04288_),
    .Y(_04397_));
 sky130_fd_sc_hd__xnor2_1 _11322_ (.A(_04396_),
    .B(_04397_),
    .Y(_04398_));
 sky130_fd_sc_hd__nand2b_1 _11323_ (.A_N(_04398_),
    .B(_04390_),
    .Y(_04399_));
 sky130_fd_sc_hd__xnor2_2 _11324_ (.A(_04390_),
    .B(_04398_),
    .Y(_04401_));
 sky130_fd_sc_hd__nand2_1 _11325_ (.A(_04389_),
    .B(_04401_),
    .Y(_04402_));
 sky130_fd_sc_hd__xnor2_2 _11326_ (.A(_04389_),
    .B(_04401_),
    .Y(_04403_));
 sky130_fd_sc_hd__a21boi_2 _11327_ (.A1(_04283_),
    .A2(_04291_),
    .B1_N(_04293_),
    .Y(_04404_));
 sky130_fd_sc_hd__or2_1 _11328_ (.A(_04403_),
    .B(_04404_),
    .X(_04405_));
 sky130_fd_sc_hd__xnor2_2 _11329_ (.A(_04403_),
    .B(_04404_),
    .Y(_04406_));
 sky130_fd_sc_hd__a21oi_2 _11330_ (.A1(_04295_),
    .A2(_04298_),
    .B1(_04406_),
    .Y(_04407_));
 sky130_fd_sc_hd__nand3_2 _11331_ (.A(_04295_),
    .B(_04298_),
    .C(_04406_),
    .Y(_04408_));
 sky130_fd_sc_hd__nand2b_2 _11332_ (.A_N(_04407_),
    .B(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__nor2_1 _11333_ (.A(_04196_),
    .B(_04302_),
    .Y(_04410_));
 sky130_fd_sc_hd__and2_1 _11334_ (.A(_04198_),
    .B(_04410_),
    .X(_04412_));
 sky130_fd_sc_hd__o21a_1 _11335_ (.A1(_04194_),
    .A2(_04300_),
    .B1(_04301_),
    .X(_04413_));
 sky130_fd_sc_hd__a21oi_1 _11336_ (.A1(_04197_),
    .A2(_04410_),
    .B1(_04413_),
    .Y(_04414_));
 sky130_fd_sc_hd__a21bo_1 _11337_ (.A1(_03981_),
    .A2(_04412_),
    .B1_N(_04414_),
    .X(_04415_));
 sky130_fd_sc_hd__a31o_1 _11338_ (.A1(_03417_),
    .A2(_03982_),
    .A3(_04412_),
    .B1(_04415_),
    .X(_04416_));
 sky130_fd_sc_hd__nor2_1 _11339_ (.A(_04409_),
    .B(_04416_),
    .Y(_04417_));
 sky130_fd_sc_hd__and2_1 _11340_ (.A(_04409_),
    .B(_04416_),
    .X(_04418_));
 sky130_fd_sc_hd__nor2_2 _11341_ (.A(_04417_),
    .B(_04418_),
    .Y(_04419_));
 sky130_fd_sc_hd__o21ai_1 _11342_ (.A1(_04348_),
    .A2(_04419_),
    .B1(net200),
    .Y(_04420_));
 sky130_fd_sc_hd__a21oi_1 _11343_ (.A1(_04348_),
    .A2(_04419_),
    .B1(_04420_),
    .Y(_04421_));
 sky130_fd_sc_hd__a22o_1 _11344_ (.A1(net161),
    .A2(_01846_),
    .B1(_01850_),
    .B2(_01851_),
    .X(_04423_));
 sky130_fd_sc_hd__nand4_1 _11345_ (.A(net161),
    .B(_01846_),
    .C(_01850_),
    .D(_01851_),
    .Y(_04424_));
 sky130_fd_sc_hd__a21o_1 _11346_ (.A1(_06064_),
    .A2(_04314_),
    .B1(_06042_),
    .X(_04425_));
 sky130_fd_sc_hd__mux2_1 _11347_ (.A0(_06396_),
    .A1(_04425_),
    .S(net284),
    .X(_04426_));
 sky130_fd_sc_hd__nand2_1 _11348_ (.A(_06009_),
    .B(_04426_),
    .Y(_04427_));
 sky130_fd_sc_hd__or2_1 _11349_ (.A(_06009_),
    .B(_04426_),
    .X(_04428_));
 sky130_fd_sc_hd__o21ba_1 _11350_ (.A1(_04319_),
    .A2(_04321_),
    .B1_N(_04318_),
    .X(_04429_));
 sky130_fd_sc_hd__nor2_1 _11351_ (.A(reg1_val[16]),
    .B(curr_PC[16]),
    .Y(_04430_));
 sky130_fd_sc_hd__nand2_1 _11352_ (.A(reg1_val[16]),
    .B(curr_PC[16]),
    .Y(_04431_));
 sky130_fd_sc_hd__and2b_1 _11353_ (.A_N(_04430_),
    .B(_04431_),
    .X(_04432_));
 sky130_fd_sc_hd__xnor2_1 _11354_ (.A(_04429_),
    .B(_04432_),
    .Y(_04434_));
 sky130_fd_sc_hd__mux2_1 _11355_ (.A0(_04339_),
    .A1(_04434_),
    .S(net249),
    .X(_04435_));
 sky130_fd_sc_hd__or2_1 _11356_ (.A(\div_shifter[47] ),
    .B(_04332_),
    .X(_04436_));
 sky130_fd_sc_hd__a21oi_1 _11357_ (.A1(net232),
    .A2(_04436_),
    .B1(\div_shifter[48] ),
    .Y(_04437_));
 sky130_fd_sc_hd__a31o_1 _11358_ (.A1(\div_shifter[48] ),
    .A2(net232),
    .A3(_04436_),
    .B1(net192),
    .X(_04438_));
 sky130_fd_sc_hd__nor2_1 _11359_ (.A(_04437_),
    .B(_04438_),
    .Y(_04439_));
 sky130_fd_sc_hd__o21ai_1 _11360_ (.A1(_05987_),
    .A2(net197),
    .B1(net198),
    .Y(_04440_));
 sky130_fd_sc_hd__a22o_1 _11361_ (.A1(_05980_),
    .A2(net241),
    .B1(_02325_),
    .B2(_05987_),
    .X(_04441_));
 sky130_fd_sc_hd__a211o_1 _11362_ (.A1(_05998_),
    .A2(_04440_),
    .B1(_04441_),
    .C1(_04439_),
    .X(_04442_));
 sky130_fd_sc_hd__or2_1 _11363_ (.A(\div_res[15] ),
    .B(_04328_),
    .X(_04443_));
 sky130_fd_sc_hd__a21oi_1 _11364_ (.A1(net164),
    .A2(_04443_),
    .B1(\div_res[16] ),
    .Y(_04445_));
 sky130_fd_sc_hd__a31o_1 _11365_ (.A1(\div_res[16] ),
    .A2(net164),
    .A3(_04443_),
    .B1(net194),
    .X(_04446_));
 sky130_fd_sc_hd__o2bb2a_1 _11366_ (.A1_N(_02313_),
    .A2_N(_04339_),
    .B1(_04445_),
    .B2(_04446_),
    .X(_04447_));
 sky130_fd_sc_hd__o21ai_1 _11367_ (.A1(net177),
    .A2(_04325_),
    .B1(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__a211o_1 _11368_ (.A1(_06475_),
    .A2(_04435_),
    .B1(_04442_),
    .C1(_04448_),
    .X(_04449_));
 sky130_fd_sc_hd__a31o_1 _11369_ (.A1(_02317_),
    .A2(_04427_),
    .A3(_04428_),
    .B1(_04449_),
    .X(_04450_));
 sky130_fd_sc_hd__a311o_1 _11370_ (.A1(_02323_),
    .A2(_04423_),
    .A3(_04424_),
    .B1(_04450_),
    .C1(_04421_),
    .X(_04451_));
 sky130_fd_sc_hd__nand2_1 _11371_ (.A(curr_PC[16]),
    .B(_04345_),
    .Y(_04452_));
 sky130_fd_sc_hd__o21a_1 _11372_ (.A1(curr_PC[16]),
    .A2(_04345_),
    .B1(net248),
    .X(_04453_));
 sky130_fd_sc_hd__a22o_4 _11373_ (.A1(net243),
    .A2(_04451_),
    .B1(_04452_),
    .B2(_04453_),
    .X(dest_val[16]));
 sky130_fd_sc_hd__a21oi_1 _11374_ (.A1(curr_PC[16]),
    .A2(_04345_),
    .B1(curr_PC[17]),
    .Y(_04455_));
 sky130_fd_sc_hd__and3_1 _11375_ (.A(curr_PC[16]),
    .B(curr_PC[17]),
    .C(_04345_),
    .X(_04456_));
 sky130_fd_sc_hd__o21a_2 _11376_ (.A1(_04455_),
    .A2(_04456_),
    .B1(net248),
    .X(_04457_));
 sky130_fd_sc_hd__a21oi_1 _11377_ (.A1(_04347_),
    .A2(_04419_),
    .B1(net158),
    .Y(_04458_));
 sky130_fd_sc_hd__a22o_1 _11378_ (.A1(net30),
    .A2(_00408_),
    .B1(_00700_),
    .B2(net32),
    .X(_04459_));
 sky130_fd_sc_hd__xnor2_1 _11379_ (.A(net50),
    .B(_04459_),
    .Y(_04460_));
 sky130_fd_sc_hd__and2_1 _11380_ (.A(net124),
    .B(_04460_),
    .X(_04461_));
 sky130_fd_sc_hd__xnor2_1 _11381_ (.A(net124),
    .B(_04460_),
    .Y(_04462_));
 sky130_fd_sc_hd__o22a_1 _11382_ (.A1(net26),
    .A2(net12),
    .B1(net8),
    .B2(_00323_),
    .X(_04463_));
 sky130_fd_sc_hd__xnor2_1 _11383_ (.A(net89),
    .B(_04463_),
    .Y(_04464_));
 sky130_fd_sc_hd__and2b_1 _11384_ (.A_N(_04462_),
    .B(_04464_),
    .X(_04466_));
 sky130_fd_sc_hd__xor2_1 _11385_ (.A(_04462_),
    .B(_04464_),
    .X(_04467_));
 sky130_fd_sc_hd__or2_1 _11386_ (.A(_04363_),
    .B(_04467_),
    .X(_04468_));
 sky130_fd_sc_hd__xor2_1 _11387_ (.A(_04363_),
    .B(_04467_),
    .X(_04469_));
 sky130_fd_sc_hd__nand2b_1 _11388_ (.A_N(_04354_),
    .B(_04469_),
    .Y(_04470_));
 sky130_fd_sc_hd__xnor2_1 _11389_ (.A(_04354_),
    .B(_04469_),
    .Y(_04471_));
 sky130_fd_sc_hd__a22o_1 _11390_ (.A1(_06563_),
    .A2(_00249_),
    .B1(net42),
    .B2(_06540_),
    .X(_04472_));
 sky130_fd_sc_hd__xor2_1 _11391_ (.A(net93),
    .B(_04472_),
    .X(_04473_));
 sky130_fd_sc_hd__o22a_1 _11392_ (.A1(net55),
    .A2(_00223_),
    .B1(net46),
    .B2(net67),
    .X(_04474_));
 sky130_fd_sc_hd__xnor2_1 _11393_ (.A(net96),
    .B(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__and2_1 _11394_ (.A(_04473_),
    .B(_04475_),
    .X(_04477_));
 sky130_fd_sc_hd__nor2_1 _11395_ (.A(_04473_),
    .B(_04475_),
    .Y(_04478_));
 sky130_fd_sc_hd__nor2_1 _11396_ (.A(_04477_),
    .B(_04478_),
    .Y(_04479_));
 sky130_fd_sc_hd__a22o_1 _11397_ (.A1(_06525_),
    .A2(net40),
    .B1(net38),
    .B2(_06559_),
    .X(_04480_));
 sky130_fd_sc_hd__xor2_1 _11398_ (.A(_00245_),
    .B(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__xor2_1 _11399_ (.A(_04479_),
    .B(_04481_),
    .X(_04482_));
 sky130_fd_sc_hd__nand2_1 _11400_ (.A(_04471_),
    .B(_04482_),
    .Y(_04483_));
 sky130_fd_sc_hd__or2_1 _11401_ (.A(_04471_),
    .B(_04482_),
    .X(_04484_));
 sky130_fd_sc_hd__o22a_1 _11402_ (.A1(net52),
    .A2(net10),
    .B1(net5),
    .B2(net101),
    .X(_04485_));
 sky130_fd_sc_hd__xnor2_1 _11403_ (.A(net20),
    .B(_04485_),
    .Y(_04486_));
 sky130_fd_sc_hd__o22a_1 _11404_ (.A1(net62),
    .A2(net23),
    .B1(net15),
    .B2(net54),
    .X(_04488_));
 sky130_fd_sc_hd__xnor2_1 _11405_ (.A(net69),
    .B(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__nor2_1 _11406_ (.A(net99),
    .B(net20),
    .Y(_04490_));
 sky130_fd_sc_hd__xnor2_1 _11407_ (.A(_04489_),
    .B(_04490_),
    .Y(_04491_));
 sky130_fd_sc_hd__nand2b_1 _11408_ (.A_N(_04486_),
    .B(_04491_),
    .Y(_04492_));
 sky130_fd_sc_hd__xnor2_1 _11409_ (.A(_04486_),
    .B(_04491_),
    .Y(_04493_));
 sky130_fd_sc_hd__and3_1 _11410_ (.A(_04483_),
    .B(_04484_),
    .C(_04493_),
    .X(_04494_));
 sky130_fd_sc_hd__a21oi_1 _11411_ (.A1(_04483_),
    .A2(_04484_),
    .B1(_04493_),
    .Y(_04495_));
 sky130_fd_sc_hd__nor2_1 _11412_ (.A(_04494_),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__o21ba_1 _11413_ (.A1(_04368_),
    .A2(_04379_),
    .B1_N(_04388_),
    .X(_04497_));
 sky130_fd_sc_hd__o21ai_2 _11414_ (.A1(_04381_),
    .A2(_04383_),
    .B1(_04385_),
    .Y(_04499_));
 sky130_fd_sc_hd__a21oi_1 _11415_ (.A1(_04371_),
    .A2(_04373_),
    .B1(_04377_),
    .Y(_04500_));
 sky130_fd_sc_hd__o21ba_1 _11416_ (.A1(_04357_),
    .A2(_04366_),
    .B1_N(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__or3b_1 _11417_ (.A(_04357_),
    .B(_04366_),
    .C_N(_04500_),
    .X(_04502_));
 sky130_fd_sc_hd__and2b_1 _11418_ (.A_N(_04501_),
    .B(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__xnor2_2 _11419_ (.A(_04499_),
    .B(_04503_),
    .Y(_04504_));
 sky130_fd_sc_hd__a21o_1 _11420_ (.A1(_04391_),
    .A2(_04395_),
    .B1(_04393_),
    .X(_04505_));
 sky130_fd_sc_hd__nand2b_1 _11421_ (.A_N(_04504_),
    .B(_04505_),
    .Y(_04506_));
 sky130_fd_sc_hd__xnor2_2 _11422_ (.A(_04504_),
    .B(_04505_),
    .Y(_04507_));
 sky130_fd_sc_hd__nand2b_1 _11423_ (.A_N(_04497_),
    .B(_04507_),
    .Y(_04508_));
 sky130_fd_sc_hd__xnor2_2 _11424_ (.A(_04497_),
    .B(_04507_),
    .Y(_04510_));
 sky130_fd_sc_hd__nand2_1 _11425_ (.A(_04496_),
    .B(_04510_),
    .Y(_04511_));
 sky130_fd_sc_hd__xnor2_2 _11426_ (.A(_04496_),
    .B(_04510_),
    .Y(_04512_));
 sky130_fd_sc_hd__o21ai_2 _11427_ (.A1(_04396_),
    .A2(_04397_),
    .B1(_04399_),
    .Y(_04513_));
 sky130_fd_sc_hd__nand2b_1 _11428_ (.A_N(_04512_),
    .B(_04513_),
    .Y(_04514_));
 sky130_fd_sc_hd__xor2_2 _11429_ (.A(_04512_),
    .B(_04513_),
    .X(_04515_));
 sky130_fd_sc_hd__a21oi_2 _11430_ (.A1(_04402_),
    .A2(_04405_),
    .B1(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__nand3_2 _11431_ (.A(_04402_),
    .B(_04405_),
    .C(_04515_),
    .Y(_04517_));
 sky130_fd_sc_hd__nand2b_2 _11432_ (.A_N(_04516_),
    .B(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__nor2_1 _11433_ (.A(_04302_),
    .B(_04409_),
    .Y(_04519_));
 sky130_fd_sc_hd__and2_1 _11434_ (.A(_04304_),
    .B(_04519_),
    .X(_04521_));
 sky130_fd_sc_hd__inv_2 _11435_ (.A(_04521_),
    .Y(_04522_));
 sky130_fd_sc_hd__o21a_1 _11436_ (.A1(_04300_),
    .A2(_04407_),
    .B1(_04408_),
    .X(_04523_));
 sky130_fd_sc_hd__a21o_1 _11437_ (.A1(_04303_),
    .A2(_04519_),
    .B1(_04523_),
    .X(_04524_));
 sky130_fd_sc_hd__a21oi_1 _11438_ (.A1(_04090_),
    .A2(_04521_),
    .B1(_04524_),
    .Y(_04525_));
 sky130_fd_sc_hd__o31ai_4 _11439_ (.A1(_03630_),
    .A2(_04088_),
    .A3(_04522_),
    .B1(_04525_),
    .Y(_04526_));
 sky130_fd_sc_hd__xnor2_4 _11440_ (.A(_04518_),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__inv_2 _11441_ (.A(_04527_),
    .Y(_04528_));
 sky130_fd_sc_hd__o21ai_1 _11442_ (.A1(_04458_),
    .A2(_04527_),
    .B1(net200),
    .Y(_04529_));
 sky130_fd_sc_hd__a21o_1 _11443_ (.A1(_04458_),
    .A2(_04527_),
    .B1(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__nor3_1 _11444_ (.A(net157),
    .B(_01852_),
    .C(_01853_),
    .Y(_04532_));
 sky130_fd_sc_hd__o21a_1 _11445_ (.A1(net157),
    .A2(_01852_),
    .B1(_01853_),
    .X(_04533_));
 sky130_fd_sc_hd__a21o_1 _11446_ (.A1(_05998_),
    .A2(_04425_),
    .B1(_05987_),
    .X(_04534_));
 sky130_fd_sc_hd__nand2_1 _11447_ (.A(net284),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__o21ai_1 _11448_ (.A1(net284),
    .A2(_06398_),
    .B1(_04535_),
    .Y(_04536_));
 sky130_fd_sc_hd__xor2_1 _11449_ (.A(_05956_),
    .B(_04536_),
    .X(_04537_));
 sky130_fd_sc_hd__o21a_1 _11450_ (.A1(_04429_),
    .A2(_04430_),
    .B1(_04431_),
    .X(_04538_));
 sky130_fd_sc_hd__nor2_1 _11451_ (.A(reg1_val[17]),
    .B(curr_PC[17]),
    .Y(_04539_));
 sky130_fd_sc_hd__nand2_1 _11452_ (.A(reg1_val[17]),
    .B(curr_PC[17]),
    .Y(_04540_));
 sky130_fd_sc_hd__nand2b_1 _11453_ (.A_N(_04539_),
    .B(_04540_),
    .Y(_04541_));
 sky130_fd_sc_hd__xnor2_1 _11454_ (.A(_04538_),
    .B(_04541_),
    .Y(_04543_));
 sky130_fd_sc_hd__nor2_1 _11455_ (.A(net249),
    .B(_04232_),
    .Y(_04544_));
 sky130_fd_sc_hd__a211o_1 _11456_ (.A1(net250),
    .A2(_04543_),
    .B1(_04544_),
    .C1(_06476_),
    .X(_04545_));
 sky130_fd_sc_hd__o21ai_1 _11457_ (.A1(_05943_),
    .A2(net197),
    .B1(net198),
    .Y(_04546_));
 sky130_fd_sc_hd__o21ai_1 _11458_ (.A1(_05934_),
    .A2(net209),
    .B1(net245),
    .Y(_04547_));
 sky130_fd_sc_hd__a221o_1 _11459_ (.A1(_05943_),
    .A2(_02325_),
    .B1(_04546_),
    .B2(_05950_),
    .C1(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__a21oi_1 _11460_ (.A1(_02313_),
    .A2(_04232_),
    .B1(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__or2_1 _11461_ (.A(\div_res[16] ),
    .B(_04443_),
    .X(_04550_));
 sky130_fd_sc_hd__and3_1 _11462_ (.A(\div_res[17] ),
    .B(net164),
    .C(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__a21oi_1 _11463_ (.A1(net164),
    .A2(_04550_),
    .B1(\div_res[17] ),
    .Y(_04552_));
 sky130_fd_sc_hd__o21a_1 _11464_ (.A1(\div_shifter[48] ),
    .A2(_04436_),
    .B1(net232),
    .X(_04554_));
 sky130_fd_sc_hd__o21ai_1 _11465_ (.A1(\div_shifter[49] ),
    .A2(_04554_),
    .B1(_02330_),
    .Y(_04555_));
 sky130_fd_sc_hd__a21o_1 _11466_ (.A1(\div_shifter[49] ),
    .A2(_04554_),
    .B1(_04555_),
    .X(_04556_));
 sky130_fd_sc_hd__o31a_1 _11467_ (.A1(net194),
    .A2(_04551_),
    .A3(_04552_),
    .B1(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__o211a_1 _11468_ (.A1(net177),
    .A2(_04218_),
    .B1(_04549_),
    .C1(_04557_),
    .X(_04558_));
 sky130_fd_sc_hd__o211a_1 _11469_ (.A1(net236),
    .A2(_04537_),
    .B1(_04545_),
    .C1(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__o311a_2 _11470_ (.A1(_02324_),
    .A2(_04532_),
    .A3(_04533_),
    .B1(_04559_),
    .C1(_04530_),
    .X(_04560_));
 sky130_fd_sc_hd__nor2_8 _11471_ (.A(_04457_),
    .B(_04560_),
    .Y(dest_val[17]));
 sky130_fd_sc_hd__and3_1 _11472_ (.A(_04347_),
    .B(_04419_),
    .C(_04528_),
    .X(_04561_));
 sky130_fd_sc_hd__nand2_1 _11473_ (.A(_00322_),
    .B(net9),
    .Y(_04562_));
 sky130_fd_sc_hd__a22o_4 _11474_ (.A1(_00326_),
    .A2(net9),
    .B1(_04562_),
    .B2(net89),
    .X(_04564_));
 sky130_fd_sc_hd__o21a_1 _11475_ (.A1(net101),
    .A2(net18),
    .B1(_04564_),
    .X(_04565_));
 sky130_fd_sc_hd__nor3_1 _11476_ (.A(net101),
    .B(net18),
    .C(_04564_),
    .Y(_04566_));
 sky130_fd_sc_hd__nor2_1 _11477_ (.A(_04565_),
    .B(_04566_),
    .Y(_04567_));
 sky130_fd_sc_hd__o21a_1 _11478_ (.A1(_04461_),
    .A2(_04466_),
    .B1(_04567_),
    .X(_04568_));
 sky130_fd_sc_hd__nor3_1 _11479_ (.A(_04461_),
    .B(_04466_),
    .C(_04567_),
    .Y(_04569_));
 sky130_fd_sc_hd__nor2_1 _11480_ (.A(_04568_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__a22o_1 _11481_ (.A1(_06517_),
    .A2(net40),
    .B1(net38),
    .B2(_06525_),
    .X(_04571_));
 sky130_fd_sc_hd__xor2_1 _11482_ (.A(net90),
    .B(_04571_),
    .X(_04572_));
 sky130_fd_sc_hd__a22o_1 _11483_ (.A1(net30),
    .A2(_00700_),
    .B1(_01951_),
    .B2(net32),
    .X(_04573_));
 sky130_fd_sc_hd__xnor2_1 _11484_ (.A(_00217_),
    .B(_04573_),
    .Y(_04575_));
 sky130_fd_sc_hd__and2_1 _11485_ (.A(_04572_),
    .B(_04575_),
    .X(_04576_));
 sky130_fd_sc_hd__nor2_1 _11486_ (.A(_04572_),
    .B(_04575_),
    .Y(_04577_));
 sky130_fd_sc_hd__nor2_1 _11487_ (.A(_04576_),
    .B(_04577_),
    .Y(_04578_));
 sky130_fd_sc_hd__o22a_1 _11488_ (.A1(net55),
    .A2(net45),
    .B1(net17),
    .B2(net47),
    .X(_04579_));
 sky130_fd_sc_hd__xnor2_1 _11489_ (.A(net95),
    .B(_04579_),
    .Y(_04580_));
 sky130_fd_sc_hd__xor2_1 _11490_ (.A(_04578_),
    .B(_04580_),
    .X(_04581_));
 sky130_fd_sc_hd__nand2_1 _11491_ (.A(_04570_),
    .B(_04581_),
    .Y(_04582_));
 sky130_fd_sc_hd__or2_1 _11492_ (.A(_04570_),
    .B(_04581_),
    .X(_04583_));
 sky130_fd_sc_hd__nand2_1 _11493_ (.A(_04582_),
    .B(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__o22a_1 _11494_ (.A1(net64),
    .A2(net23),
    .B1(net15),
    .B2(net62),
    .X(_04586_));
 sky130_fd_sc_hd__xnor2_2 _11495_ (.A(net69),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__o22a_1 _11496_ (.A1(net54),
    .A2(net10),
    .B1(net5),
    .B2(net52),
    .X(_04588_));
 sky130_fd_sc_hd__xnor2_1 _11497_ (.A(net21),
    .B(_04588_),
    .Y(_04589_));
 sky130_fd_sc_hd__a22o_1 _11498_ (.A1(_06559_),
    .A2(net43),
    .B1(net41),
    .B2(_06563_),
    .X(_04590_));
 sky130_fd_sc_hd__xor2_1 _11499_ (.A(net93),
    .B(_04590_),
    .X(_04591_));
 sky130_fd_sc_hd__nand2b_1 _11500_ (.A_N(_04589_),
    .B(_04591_),
    .Y(_04592_));
 sky130_fd_sc_hd__nand2b_1 _11501_ (.A_N(_04591_),
    .B(_04589_),
    .Y(_04593_));
 sky130_fd_sc_hd__nand2_1 _11502_ (.A(_04592_),
    .B(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__xnor2_2 _11503_ (.A(_04587_),
    .B(_04594_),
    .Y(_04595_));
 sky130_fd_sc_hd__xor2_1 _11504_ (.A(_04584_),
    .B(_04595_),
    .X(_04597_));
 sky130_fd_sc_hd__a21o_1 _11505_ (.A1(_04471_),
    .A2(_04482_),
    .B1(_04494_),
    .X(_04598_));
 sky130_fd_sc_hd__o31a_1 _11506_ (.A1(net99),
    .A2(net20),
    .A3(_04489_),
    .B1(_04492_),
    .X(_04599_));
 sky130_fd_sc_hd__a21oi_1 _11507_ (.A1(_04479_),
    .A2(_04481_),
    .B1(_04477_),
    .Y(_04600_));
 sky130_fd_sc_hd__a21oi_1 _11508_ (.A1(_04468_),
    .A2(_04470_),
    .B1(_04600_),
    .Y(_04601_));
 sky130_fd_sc_hd__and3_1 _11509_ (.A(_04468_),
    .B(_04470_),
    .C(_04600_),
    .X(_04602_));
 sky130_fd_sc_hd__nor2_1 _11510_ (.A(_04601_),
    .B(_04602_),
    .Y(_04603_));
 sky130_fd_sc_hd__xor2_1 _11511_ (.A(_04599_),
    .B(_04603_),
    .X(_04604_));
 sky130_fd_sc_hd__a21oi_1 _11512_ (.A1(_04499_),
    .A2(_04502_),
    .B1(_04501_),
    .Y(_04605_));
 sky130_fd_sc_hd__or2_1 _11513_ (.A(_04604_),
    .B(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__xnor2_1 _11514_ (.A(_04604_),
    .B(_04605_),
    .Y(_04608_));
 sky130_fd_sc_hd__nand2b_1 _11515_ (.A_N(_04608_),
    .B(_04598_),
    .Y(_04609_));
 sky130_fd_sc_hd__xnor2_1 _11516_ (.A(_04598_),
    .B(_04608_),
    .Y(_04610_));
 sky130_fd_sc_hd__nand2_1 _11517_ (.A(_04597_),
    .B(_04610_),
    .Y(_04611_));
 sky130_fd_sc_hd__or2_1 _11518_ (.A(_04597_),
    .B(_04610_),
    .X(_04612_));
 sky130_fd_sc_hd__nand2_1 _11519_ (.A(_04611_),
    .B(_04612_),
    .Y(_04613_));
 sky130_fd_sc_hd__nand2_1 _11520_ (.A(_04506_),
    .B(_04508_),
    .Y(_04614_));
 sky130_fd_sc_hd__nand2b_1 _11521_ (.A_N(_04613_),
    .B(_04614_),
    .Y(_04615_));
 sky130_fd_sc_hd__xor2_2 _11522_ (.A(_04613_),
    .B(_04614_),
    .X(_04616_));
 sky130_fd_sc_hd__a21oi_2 _11523_ (.A1(_04511_),
    .A2(_04514_),
    .B1(_04616_),
    .Y(_04617_));
 sky130_fd_sc_hd__nand3_2 _11524_ (.A(_04511_),
    .B(_04514_),
    .C(_04616_),
    .Y(_04619_));
 sky130_fd_sc_hd__nand2b_4 _11525_ (.A_N(_04617_),
    .B(_04619_),
    .Y(_04620_));
 sky130_fd_sc_hd__nor2_1 _11526_ (.A(_04409_),
    .B(_04518_),
    .Y(_04621_));
 sky130_fd_sc_hd__and2_1 _11527_ (.A(_04410_),
    .B(_04621_),
    .X(_04622_));
 sky130_fd_sc_hd__nand2_1 _11528_ (.A(_04410_),
    .B(_04621_),
    .Y(_04623_));
 sky130_fd_sc_hd__o21a_1 _11529_ (.A1(_04407_),
    .A2(_04516_),
    .B1(_04517_),
    .X(_04624_));
 sky130_fd_sc_hd__a21o_1 _11530_ (.A1(_04413_),
    .A2(_04621_),
    .B1(_04624_),
    .X(_04625_));
 sky130_fd_sc_hd__a21o_1 _11531_ (.A1(_04199_),
    .A2(_04622_),
    .B1(_04625_),
    .X(_04626_));
 sky130_fd_sc_hd__a31o_1 _11532_ (.A1(net3),
    .A2(_04200_),
    .A3(_04622_),
    .B1(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__xor2_4 _11533_ (.A(_04620_),
    .B(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__o21ai_1 _11534_ (.A1(net158),
    .A2(_04561_),
    .B1(_04628_),
    .Y(_04629_));
 sky130_fd_sc_hd__o31a_1 _11535_ (.A1(net158),
    .A2(_04561_),
    .A3(_04628_),
    .B1(net200),
    .X(_04630_));
 sky130_fd_sc_hd__nand2_1 _11536_ (.A(_04629_),
    .B(_04630_),
    .Y(_04631_));
 sky130_fd_sc_hd__a21oi_1 _11537_ (.A1(net162),
    .A2(_01854_),
    .B1(_01858_),
    .Y(_04632_));
 sky130_fd_sc_hd__and3_1 _11538_ (.A(net162),
    .B(_01854_),
    .C(_01858_),
    .X(_04633_));
 sky130_fd_sc_hd__a21oi_1 _11539_ (.A1(_05950_),
    .A2(_04534_),
    .B1(_05943_),
    .Y(_04634_));
 sky130_fd_sc_hd__mux2_1 _11540_ (.A0(_06400_),
    .A1(_04634_),
    .S(net284),
    .X(_04635_));
 sky130_fd_sc_hd__nand2_1 _11541_ (.A(_05907_),
    .B(_04635_),
    .Y(_04636_));
 sky130_fd_sc_hd__o21a_1 _11542_ (.A1(_05907_),
    .A2(_04635_),
    .B1(_02317_),
    .X(_04637_));
 sky130_fd_sc_hd__nand2_1 _11543_ (.A(reg1_val[18]),
    .B(curr_PC[18]),
    .Y(_04638_));
 sky130_fd_sc_hd__or2_1 _11544_ (.A(reg1_val[18]),
    .B(curr_PC[18]),
    .X(_04640_));
 sky130_fd_sc_hd__nand2_1 _11545_ (.A(_04638_),
    .B(_04640_),
    .Y(_04641_));
 sky130_fd_sc_hd__o21ai_1 _11546_ (.A1(_04538_),
    .A2(_04539_),
    .B1(_04540_),
    .Y(_04642_));
 sky130_fd_sc_hd__xor2_1 _11547_ (.A(_04641_),
    .B(_04642_),
    .X(_04643_));
 sky130_fd_sc_hd__mux2_1 _11548_ (.A0(_04121_),
    .A1(_04643_),
    .S(net249),
    .X(_04644_));
 sky130_fd_sc_hd__or3_1 _11549_ (.A(\div_shifter[49] ),
    .B(\div_shifter[48] ),
    .C(_04436_),
    .X(_04645_));
 sky130_fd_sc_hd__a21oi_1 _11550_ (.A1(net232),
    .A2(_04645_),
    .B1(\div_shifter[50] ),
    .Y(_04646_));
 sky130_fd_sc_hd__a31o_1 _11551_ (.A1(\div_shifter[50] ),
    .A2(net232),
    .A3(_04645_),
    .B1(net192),
    .X(_04647_));
 sky130_fd_sc_hd__or2_1 _11552_ (.A(_04646_),
    .B(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__mux2_1 _11553_ (.A0(_02319_),
    .A1(_02325_),
    .S(_05889_),
    .X(_04649_));
 sky130_fd_sc_hd__nor2_1 _11554_ (.A(_02315_),
    .B(_04649_),
    .Y(_04650_));
 sky130_fd_sc_hd__o22a_1 _11555_ (.A1(_05872_),
    .A2(net209),
    .B1(_04650_),
    .B2(_05898_),
    .X(_04651_));
 sky130_fd_sc_hd__o221a_1 _11556_ (.A1(net177),
    .A2(_04108_),
    .B1(_04121_),
    .B2(_02314_),
    .C1(_04651_),
    .X(_04652_));
 sky130_fd_sc_hd__or2_1 _11557_ (.A(\div_res[17] ),
    .B(_04550_),
    .X(_04653_));
 sky130_fd_sc_hd__a21oi_1 _11558_ (.A1(net164),
    .A2(_04653_),
    .B1(\div_res[18] ),
    .Y(_04654_));
 sky130_fd_sc_hd__a31o_1 _11559_ (.A1(\div_res[18] ),
    .A2(net164),
    .A3(_04653_),
    .B1(net194),
    .X(_04655_));
 sky130_fd_sc_hd__o211a_1 _11560_ (.A1(_04654_),
    .A2(_04655_),
    .B1(_04648_),
    .C1(_04652_),
    .X(_04656_));
 sky130_fd_sc_hd__o21ai_1 _11561_ (.A1(_06476_),
    .A2(_04644_),
    .B1(_04656_),
    .Y(_04657_));
 sky130_fd_sc_hd__a21oi_2 _11562_ (.A1(_04636_),
    .A2(_04637_),
    .B1(_04657_),
    .Y(_04658_));
 sky130_fd_sc_hd__o311a_1 _11563_ (.A1(_02324_),
    .A2(_04632_),
    .A3(_04633_),
    .B1(_04658_),
    .C1(_04631_),
    .X(_04659_));
 sky130_fd_sc_hd__and2_2 _11564_ (.A(curr_PC[18]),
    .B(_04456_),
    .X(_04661_));
 sky130_fd_sc_hd__o21ai_1 _11565_ (.A1(curr_PC[18]),
    .A2(_04456_),
    .B1(net248),
    .Y(_04662_));
 sky130_fd_sc_hd__o22ai_4 _11566_ (.A1(net248),
    .A2(_04659_),
    .B1(_04661_),
    .B2(_04662_),
    .Y(dest_val[18]));
 sky130_fd_sc_hd__and4_1 _11567_ (.A(_04347_),
    .B(_04419_),
    .C(_04528_),
    .D(_04628_),
    .X(_04663_));
 sky130_fd_sc_hd__o22a_1 _11568_ (.A1(net58),
    .A2(net23),
    .B1(net15),
    .B2(net64),
    .X(_04664_));
 sky130_fd_sc_hd__xnor2_1 _11569_ (.A(net69),
    .B(_04664_),
    .Y(_04665_));
 sky130_fd_sc_hd__a22o_1 _11570_ (.A1(_00143_),
    .A2(net40),
    .B1(net38),
    .B2(_06517_),
    .X(_04666_));
 sky130_fd_sc_hd__xor2_1 _11571_ (.A(net90),
    .B(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__nand2b_1 _11572_ (.A_N(_04665_),
    .B(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__nand2b_1 _11573_ (.A_N(_04667_),
    .B(_04665_),
    .Y(_04669_));
 sky130_fd_sc_hd__nand2_1 _11574_ (.A(_04668_),
    .B(_04669_),
    .Y(_04670_));
 sky130_fd_sc_hd__a22o_1 _11575_ (.A1(_06525_),
    .A2(net43),
    .B1(net41),
    .B2(_06559_),
    .X(_04671_));
 sky130_fd_sc_hd__xor2_2 _11576_ (.A(net93),
    .B(_04671_),
    .X(_04672_));
 sky130_fd_sc_hd__nand2b_1 _11577_ (.A_N(_04670_),
    .B(_04672_),
    .Y(_04673_));
 sky130_fd_sc_hd__xnor2_2 _11578_ (.A(_04670_),
    .B(_04672_),
    .Y(_04674_));
 sky130_fd_sc_hd__o22a_1 _11579_ (.A1(net45),
    .A2(net17),
    .B1(net14),
    .B2(net47),
    .X(_04675_));
 sky130_fd_sc_hd__xor2_1 _11580_ (.A(net95),
    .B(_04675_),
    .X(_04676_));
 sky130_fd_sc_hd__or2_1 _11581_ (.A(net89),
    .B(_04676_),
    .X(_04677_));
 sky130_fd_sc_hd__xnor2_1 _11582_ (.A(net89),
    .B(_04676_),
    .Y(_04678_));
 sky130_fd_sc_hd__a22o_1 _11583_ (.A1(net30),
    .A2(_01951_),
    .B1(_02066_),
    .B2(net32),
    .X(_04679_));
 sky130_fd_sc_hd__xnor2_1 _11584_ (.A(_00216_),
    .B(_04679_),
    .Y(_04681_));
 sky130_fd_sc_hd__or2_2 _11585_ (.A(_04678_),
    .B(_04681_),
    .X(_04682_));
 sky130_fd_sc_hd__nand2_1 _11586_ (.A(_04678_),
    .B(_04681_),
    .Y(_04683_));
 sky130_fd_sc_hd__nand2_1 _11587_ (.A(_04682_),
    .B(_04683_),
    .Y(_04684_));
 sky130_fd_sc_hd__o22a_2 _11588_ (.A1(net62),
    .A2(net10),
    .B1(net5),
    .B2(net54),
    .X(_04685_));
 sky130_fd_sc_hd__xnor2_4 _11589_ (.A(net22),
    .B(_04685_),
    .Y(_04686_));
 sky130_fd_sc_hd__nand2_1 _11590_ (.A(_04564_),
    .B(_04686_),
    .Y(_04687_));
 sky130_fd_sc_hd__xnor2_4 _11591_ (.A(_04564_),
    .B(_04686_),
    .Y(_04688_));
 sky130_fd_sc_hd__nand2_2 _11592_ (.A(_00172_),
    .B(_02078_),
    .Y(_04689_));
 sky130_fd_sc_hd__xor2_4 _11593_ (.A(_04688_),
    .B(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__xnor2_2 _11594_ (.A(_04684_),
    .B(_04690_),
    .Y(_04691_));
 sky130_fd_sc_hd__xor2_1 _11595_ (.A(_04674_),
    .B(_04691_),
    .X(_04692_));
 sky130_fd_sc_hd__o21ai_1 _11596_ (.A1(_04584_),
    .A2(_04595_),
    .B1(_04582_),
    .Y(_04693_));
 sky130_fd_sc_hd__o21ai_2 _11597_ (.A1(_04587_),
    .A2(_04594_),
    .B1(_04592_),
    .Y(_04694_));
 sky130_fd_sc_hd__a21oi_1 _11598_ (.A1(_04578_),
    .A2(_04580_),
    .B1(_04576_),
    .Y(_04695_));
 sky130_fd_sc_hd__o21bai_2 _11599_ (.A1(_04566_),
    .A2(_04568_),
    .B1_N(_04695_),
    .Y(_04696_));
 sky130_fd_sc_hd__or3b_1 _11600_ (.A(_04566_),
    .B(_04568_),
    .C_N(_04695_),
    .X(_04697_));
 sky130_fd_sc_hd__nand2_1 _11601_ (.A(_04696_),
    .B(_04697_),
    .Y(_04698_));
 sky130_fd_sc_hd__nand2b_1 _11602_ (.A_N(_04698_),
    .B(_04694_),
    .Y(_04699_));
 sky130_fd_sc_hd__xor2_1 _11603_ (.A(_04694_),
    .B(_04698_),
    .X(_04700_));
 sky130_fd_sc_hd__o21ba_1 _11604_ (.A1(_04599_),
    .A2(_04602_),
    .B1_N(_04601_),
    .X(_04702_));
 sky130_fd_sc_hd__or2_1 _11605_ (.A(_04700_),
    .B(_04702_),
    .X(_04703_));
 sky130_fd_sc_hd__nand2_1 _11606_ (.A(_04700_),
    .B(_04702_),
    .Y(_04704_));
 sky130_fd_sc_hd__nand2_1 _11607_ (.A(_04703_),
    .B(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__nand2b_1 _11608_ (.A_N(_04705_),
    .B(_04693_),
    .Y(_04706_));
 sky130_fd_sc_hd__xnor2_1 _11609_ (.A(_04693_),
    .B(_04705_),
    .Y(_04707_));
 sky130_fd_sc_hd__xnor2_1 _11610_ (.A(_04692_),
    .B(_04707_),
    .Y(_04708_));
 sky130_fd_sc_hd__a21oi_1 _11611_ (.A1(_04606_),
    .A2(_04609_),
    .B1(_04708_),
    .Y(_04709_));
 sky130_fd_sc_hd__and3_1 _11612_ (.A(_04606_),
    .B(_04609_),
    .C(_04708_),
    .X(_04710_));
 sky130_fd_sc_hd__or2_1 _11613_ (.A(_04709_),
    .B(_04710_),
    .X(_04711_));
 sky130_fd_sc_hd__a21o_1 _11614_ (.A1(_04611_),
    .A2(_04615_),
    .B1(_04711_),
    .X(_04712_));
 sky130_fd_sc_hd__inv_2 _11615_ (.A(_04712_),
    .Y(_04713_));
 sky130_fd_sc_hd__nand3_1 _11616_ (.A(_04611_),
    .B(_04615_),
    .C(_04711_),
    .Y(_04714_));
 sky130_fd_sc_hd__nand2_2 _11617_ (.A(_04712_),
    .B(_04714_),
    .Y(_04715_));
 sky130_fd_sc_hd__nor2_1 _11618_ (.A(_04518_),
    .B(_04620_),
    .Y(_04716_));
 sky130_fd_sc_hd__nand2_1 _11619_ (.A(_04519_),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__inv_2 _11620_ (.A(_04717_),
    .Y(_04718_));
 sky130_fd_sc_hd__o21a_1 _11621_ (.A1(_04516_),
    .A2(_04617_),
    .B1(_04619_),
    .X(_04719_));
 sky130_fd_sc_hd__a21o_1 _11622_ (.A1(_04523_),
    .A2(_04716_),
    .B1(_04719_),
    .X(_04720_));
 sky130_fd_sc_hd__and3_1 _11623_ (.A(_04305_),
    .B(_04519_),
    .C(_04716_),
    .X(_04721_));
 sky130_fd_sc_hd__a311o_2 _11624_ (.A1(_03864_),
    .A2(_04306_),
    .A3(_04718_),
    .B1(_04720_),
    .C1(_04721_),
    .X(_04723_));
 sky130_fd_sc_hd__xnor2_4 _11625_ (.A(_04715_),
    .B(_04723_),
    .Y(_04724_));
 sky130_fd_sc_hd__inv_2 _11626_ (.A(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__o21a_1 _11627_ (.A1(net158),
    .A2(_04663_),
    .B1(_04725_),
    .X(_04726_));
 sky130_fd_sc_hd__o31ai_1 _11628_ (.A1(net158),
    .A2(_04663_),
    .A3(_04725_),
    .B1(net200),
    .Y(_04727_));
 sky130_fd_sc_hd__o21ai_1 _11629_ (.A1(net157),
    .A2(_01859_),
    .B1(_01861_),
    .Y(_04728_));
 sky130_fd_sc_hd__or3_1 _11630_ (.A(net157),
    .B(_01859_),
    .C(_01861_),
    .X(_04729_));
 sky130_fd_sc_hd__nand2_1 _11631_ (.A(_04728_),
    .B(_04729_),
    .Y(_04730_));
 sky130_fd_sc_hd__or2_1 _11632_ (.A(net284),
    .B(_06402_),
    .X(_04731_));
 sky130_fd_sc_hd__o21ba_1 _11633_ (.A1(_05907_),
    .A2(_04634_),
    .B1_N(_05889_),
    .X(_04732_));
 sky130_fd_sc_hd__or2_1 _11634_ (.A(net295),
    .B(_04732_),
    .X(_04733_));
 sky130_fd_sc_hd__a21oi_1 _11635_ (.A1(_04731_),
    .A2(_04733_),
    .B1(_05845_),
    .Y(_04734_));
 sky130_fd_sc_hd__and3_1 _11636_ (.A(_05845_),
    .B(_04731_),
    .C(_04733_),
    .X(_04735_));
 sky130_fd_sc_hd__or3_1 _11637_ (.A(net236),
    .B(_04734_),
    .C(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__nand2_1 _11638_ (.A(reg1_val[19]),
    .B(curr_PC[19]),
    .Y(_04737_));
 sky130_fd_sc_hd__or2_1 _11639_ (.A(reg1_val[19]),
    .B(curr_PC[19]),
    .X(_04738_));
 sky130_fd_sc_hd__nand2_1 _11640_ (.A(_04737_),
    .B(_04738_),
    .Y(_04739_));
 sky130_fd_sc_hd__a21boi_1 _11641_ (.A1(_04640_),
    .A2(_04642_),
    .B1_N(_04638_),
    .Y(_04740_));
 sky130_fd_sc_hd__xnor2_1 _11642_ (.A(_04739_),
    .B(_04740_),
    .Y(_04741_));
 sky130_fd_sc_hd__nor2_1 _11643_ (.A(net250),
    .B(_04010_),
    .Y(_04742_));
 sky130_fd_sc_hd__a211o_1 _11644_ (.A1(net249),
    .A2(_04741_),
    .B1(_04742_),
    .C1(_06476_),
    .X(_04744_));
 sky130_fd_sc_hd__or2_1 _11645_ (.A(\div_res[18] ),
    .B(_04653_),
    .X(_04745_));
 sky130_fd_sc_hd__and3_1 _11646_ (.A(\div_res[19] ),
    .B(net164),
    .C(_04745_),
    .X(_04746_));
 sky130_fd_sc_hd__a21oi_1 _11647_ (.A1(net164),
    .A2(_04745_),
    .B1(\div_res[19] ),
    .Y(_04747_));
 sky130_fd_sc_hd__or3_1 _11648_ (.A(net194),
    .B(_04746_),
    .C(_04747_),
    .X(_04748_));
 sky130_fd_sc_hd__or2_1 _11649_ (.A(\div_shifter[50] ),
    .B(_04645_),
    .X(_04749_));
 sky130_fd_sc_hd__nand3_1 _11650_ (.A(\div_shifter[51] ),
    .B(net232),
    .C(_04749_),
    .Y(_04750_));
 sky130_fd_sc_hd__a21o_1 _11651_ (.A1(net232),
    .A2(_04749_),
    .B1(\div_shifter[51] ),
    .X(_04751_));
 sky130_fd_sc_hd__mux2_1 _11652_ (.A0(_02320_),
    .A1(net196),
    .S(_05817_),
    .X(_04752_));
 sky130_fd_sc_hd__a21o_1 _11653_ (.A1(net198),
    .A2(_04752_),
    .B1(_05826_),
    .X(_04753_));
 sky130_fd_sc_hd__o21ai_1 _11654_ (.A1(_05808_),
    .A2(net209),
    .B1(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__a221o_1 _11655_ (.A1(net179),
    .A2(_03994_),
    .B1(_04010_),
    .B2(_02313_),
    .C1(_04754_),
    .X(_04755_));
 sky130_fd_sc_hd__a31o_1 _11656_ (.A1(_02330_),
    .A2(_04750_),
    .A3(_04751_),
    .B1(_04755_),
    .X(_04756_));
 sky130_fd_sc_hd__and4b_1 _11657_ (.A_N(_04756_),
    .B(_04748_),
    .C(_04744_),
    .D(_04736_),
    .X(_04757_));
 sky130_fd_sc_hd__o221a_1 _11658_ (.A1(_04726_),
    .A2(_04727_),
    .B1(_04730_),
    .B2(_02324_),
    .C1(_04757_),
    .X(_04758_));
 sky130_fd_sc_hd__a21oi_1 _11659_ (.A1(curr_PC[19]),
    .A2(_04661_),
    .B1(net243),
    .Y(_04759_));
 sky130_fd_sc_hd__o21ai_2 _11660_ (.A1(curr_PC[19]),
    .A2(_04661_),
    .B1(_04759_),
    .Y(_04760_));
 sky130_fd_sc_hd__o21ai_4 _11661_ (.A1(net248),
    .A2(_04758_),
    .B1(_04760_),
    .Y(dest_val[19]));
 sky130_fd_sc_hd__a21o_1 _11662_ (.A1(_04663_),
    .A2(_04725_),
    .B1(net158),
    .X(_04761_));
 sky130_fd_sc_hd__o22a_1 _11663_ (.A1(net45),
    .A2(net14),
    .B1(net12),
    .B2(net47),
    .X(_04762_));
 sky130_fd_sc_hd__xnor2_1 _11664_ (.A(net95),
    .B(_04762_),
    .Y(_04763_));
 sky130_fd_sc_hd__a21oi_1 _11665_ (.A1(_00310_),
    .A2(_02066_),
    .B1(_00216_),
    .Y(_04764_));
 sky130_fd_sc_hd__a31o_1 _11666_ (.A1(_00216_),
    .A2(_00303_),
    .A3(_02066_),
    .B1(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__and2b_1 _11667_ (.A_N(_04763_),
    .B(_04765_),
    .X(_04766_));
 sky130_fd_sc_hd__and2b_1 _11668_ (.A_N(_04765_),
    .B(_04763_),
    .X(_04767_));
 sky130_fd_sc_hd__nor2_1 _11669_ (.A(_04766_),
    .B(_04767_),
    .Y(_04768_));
 sky130_fd_sc_hd__o22a_1 _11670_ (.A1(net64),
    .A2(net10),
    .B1(net5),
    .B2(net62),
    .X(_04769_));
 sky130_fd_sc_hd__nand2_1 _11671_ (.A(net54),
    .B(net22),
    .Y(_04770_));
 sky130_fd_sc_hd__xnor2_1 _11672_ (.A(_04769_),
    .B(_04770_),
    .Y(_04771_));
 sky130_fd_sc_hd__or2_1 _11673_ (.A(_04768_),
    .B(_04771_),
    .X(_04772_));
 sky130_fd_sc_hd__nand2_1 _11674_ (.A(_04768_),
    .B(_04771_),
    .Y(_04774_));
 sky130_fd_sc_hd__nand2_1 _11675_ (.A(_04772_),
    .B(_04774_),
    .Y(_04775_));
 sky130_fd_sc_hd__o22a_1 _11676_ (.A1(net60),
    .A2(net23),
    .B1(net15),
    .B2(net58),
    .X(_04776_));
 sky130_fd_sc_hd__xnor2_1 _11677_ (.A(net69),
    .B(_04776_),
    .Y(_04777_));
 sky130_fd_sc_hd__o22a_1 _11678_ (.A1(net55),
    .A2(_00267_),
    .B1(net17),
    .B2(_00263_),
    .X(_04778_));
 sky130_fd_sc_hd__xnor2_1 _11679_ (.A(net90),
    .B(_04778_),
    .Y(_04779_));
 sky130_fd_sc_hd__and2b_1 _11680_ (.A_N(_04777_),
    .B(_04779_),
    .X(_04780_));
 sky130_fd_sc_hd__xor2_1 _11681_ (.A(_04777_),
    .B(_04779_),
    .X(_04781_));
 sky130_fd_sc_hd__a22o_1 _11682_ (.A1(_06517_),
    .A2(net43),
    .B1(net41),
    .B2(_06525_),
    .X(_04782_));
 sky130_fd_sc_hd__xor2_1 _11683_ (.A(net93),
    .B(_04782_),
    .X(_04783_));
 sky130_fd_sc_hd__and2b_1 _11684_ (.A_N(_04781_),
    .B(_04783_),
    .X(_04785_));
 sky130_fd_sc_hd__and2b_1 _11685_ (.A_N(_04783_),
    .B(_04781_),
    .X(_04786_));
 sky130_fd_sc_hd__or2_1 _11686_ (.A(_04785_),
    .B(_04786_),
    .X(_04787_));
 sky130_fd_sc_hd__xor2_2 _11687_ (.A(_04775_),
    .B(_04787_),
    .X(_04788_));
 sky130_fd_sc_hd__a32oi_4 _11688_ (.A1(_04682_),
    .A2(_04683_),
    .A3(_04690_),
    .B1(_04691_),
    .B2(_04674_),
    .Y(_04789_));
 sky130_fd_sc_hd__nand2_1 _11689_ (.A(_04668_),
    .B(_04673_),
    .Y(_04790_));
 sky130_fd_sc_hd__o21a_1 _11690_ (.A1(_04688_),
    .A2(_04689_),
    .B1(_04687_),
    .X(_04791_));
 sky130_fd_sc_hd__a21oi_1 _11691_ (.A1(_04677_),
    .A2(_04682_),
    .B1(_04791_),
    .Y(_04792_));
 sky130_fd_sc_hd__and3_1 _11692_ (.A(_04677_),
    .B(_04682_),
    .C(_04791_),
    .X(_04793_));
 sky130_fd_sc_hd__nor2_1 _11693_ (.A(_04792_),
    .B(_04793_),
    .Y(_04794_));
 sky130_fd_sc_hd__and2_1 _11694_ (.A(_04790_),
    .B(_04794_),
    .X(_04796_));
 sky130_fd_sc_hd__or2_1 _11695_ (.A(_04790_),
    .B(_04794_),
    .X(_04797_));
 sky130_fd_sc_hd__nand2b_1 _11696_ (.A_N(_04796_),
    .B(_04797_),
    .Y(_04798_));
 sky130_fd_sc_hd__a21oi_1 _11697_ (.A1(_04696_),
    .A2(_04699_),
    .B1(_04798_),
    .Y(_04799_));
 sky130_fd_sc_hd__and3_1 _11698_ (.A(_04696_),
    .B(_04699_),
    .C(_04798_),
    .X(_04800_));
 sky130_fd_sc_hd__nor2_1 _11699_ (.A(_04799_),
    .B(_04800_),
    .Y(_04801_));
 sky130_fd_sc_hd__and2b_1 _11700_ (.A_N(_04789_),
    .B(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__xnor2_1 _11701_ (.A(_04789_),
    .B(_04801_),
    .Y(_04803_));
 sky130_fd_sc_hd__nand2_1 _11702_ (.A(_04788_),
    .B(_04803_),
    .Y(_04804_));
 sky130_fd_sc_hd__xnor2_1 _11703_ (.A(_04788_),
    .B(_04803_),
    .Y(_04805_));
 sky130_fd_sc_hd__a21o_1 _11704_ (.A1(_04703_),
    .A2(_04706_),
    .B1(_04805_),
    .X(_04807_));
 sky130_fd_sc_hd__nand3_1 _11705_ (.A(_04703_),
    .B(_04706_),
    .C(_04805_),
    .Y(_04808_));
 sky130_fd_sc_hd__nand2_1 _11706_ (.A(_04807_),
    .B(_04808_),
    .Y(_04809_));
 sky130_fd_sc_hd__a21oi_1 _11707_ (.A1(_04692_),
    .A2(_04707_),
    .B1(_04709_),
    .Y(_04810_));
 sky130_fd_sc_hd__or2_2 _11708_ (.A(_04809_),
    .B(_04810_),
    .X(_04811_));
 sky130_fd_sc_hd__nand2_1 _11709_ (.A(_04809_),
    .B(_04810_),
    .Y(_04812_));
 sky130_fd_sc_hd__nand2_4 _11710_ (.A(_04811_),
    .B(_04812_),
    .Y(_04813_));
 sky130_fd_sc_hd__nor2_1 _11711_ (.A(_04620_),
    .B(_04715_),
    .Y(_04814_));
 sky130_fd_sc_hd__nand2_1 _11712_ (.A(_04621_),
    .B(_04814_),
    .Y(_04815_));
 sky130_fd_sc_hd__inv_2 _11713_ (.A(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__o21a_1 _11714_ (.A1(_04617_),
    .A2(_04713_),
    .B1(_04714_),
    .X(_04818_));
 sky130_fd_sc_hd__a21o_1 _11715_ (.A1(_04624_),
    .A2(_04814_),
    .B1(_04818_),
    .X(_04819_));
 sky130_fd_sc_hd__nor2_1 _11716_ (.A(_04414_),
    .B(_04815_),
    .Y(_04820_));
 sky130_fd_sc_hd__a311oi_4 _11717_ (.A1(_03983_),
    .A2(_04412_),
    .A3(_04816_),
    .B1(_04819_),
    .C1(_04820_),
    .Y(_04821_));
 sky130_fd_sc_hd__xor2_1 _11718_ (.A(_04813_),
    .B(_04821_),
    .X(_04822_));
 sky130_fd_sc_hd__xnor2_4 _11719_ (.A(_04813_),
    .B(_04821_),
    .Y(_04823_));
 sky130_fd_sc_hd__nand2_1 _11720_ (.A(_04761_),
    .B(_04823_),
    .Y(_04824_));
 sky130_fd_sc_hd__o21a_1 _11721_ (.A1(_04761_),
    .A2(_04823_),
    .B1(net200),
    .X(_04825_));
 sky130_fd_sc_hd__a21o_1 _11722_ (.A1(_01859_),
    .A2(_01861_),
    .B1(net157),
    .X(_04826_));
 sky130_fd_sc_hd__xnor2_1 _11723_ (.A(_01866_),
    .B(_04826_),
    .Y(_04827_));
 sky130_fd_sc_hd__o21bai_1 _11724_ (.A1(_05845_),
    .A2(_04732_),
    .B1_N(_05817_),
    .Y(_04829_));
 sky130_fd_sc_hd__mux2_1 _11725_ (.A0(_06404_),
    .A1(_04829_),
    .S(net284),
    .X(_04830_));
 sky130_fd_sc_hd__nand2_1 _11726_ (.A(_05696_),
    .B(_04830_),
    .Y(_04831_));
 sky130_fd_sc_hd__o211a_1 _11727_ (.A1(_05696_),
    .A2(_04830_),
    .B1(_04831_),
    .C1(_02317_),
    .X(_04832_));
 sky130_fd_sc_hd__nand2_1 _11728_ (.A(reg1_val[20]),
    .B(curr_PC[20]),
    .Y(_04833_));
 sky130_fd_sc_hd__or2_1 _11729_ (.A(reg1_val[20]),
    .B(curr_PC[20]),
    .X(_04834_));
 sky130_fd_sc_hd__nand2_1 _11730_ (.A(_04833_),
    .B(_04834_),
    .Y(_04835_));
 sky130_fd_sc_hd__o21a_1 _11731_ (.A1(_04739_),
    .A2(_04740_),
    .B1(_04737_),
    .X(_04836_));
 sky130_fd_sc_hd__xor2_1 _11732_ (.A(_04835_),
    .B(_04836_),
    .X(_04837_));
 sky130_fd_sc_hd__nand2_1 _11733_ (.A(net229),
    .B(_03896_),
    .Y(_04838_));
 sky130_fd_sc_hd__o211a_1 _11734_ (.A1(net229),
    .A2(_04837_),
    .B1(_04838_),
    .C1(_06475_),
    .X(_04840_));
 sky130_fd_sc_hd__or2_1 _11735_ (.A(\div_res[19] ),
    .B(_04745_),
    .X(_04841_));
 sky130_fd_sc_hd__a21oi_1 _11736_ (.A1(net164),
    .A2(_04841_),
    .B1(\div_res[20] ),
    .Y(_04842_));
 sky130_fd_sc_hd__a31o_1 _11737_ (.A1(\div_res[20] ),
    .A2(net164),
    .A3(_04841_),
    .B1(net194),
    .X(_04843_));
 sky130_fd_sc_hd__nor2_1 _11738_ (.A(_04842_),
    .B(_04843_),
    .Y(_04844_));
 sky130_fd_sc_hd__or2_1 _11739_ (.A(\div_shifter[51] ),
    .B(_04749_),
    .X(_04845_));
 sky130_fd_sc_hd__a21oi_1 _11740_ (.A1(net232),
    .A2(_04845_),
    .B1(\div_shifter[52] ),
    .Y(_04846_));
 sky130_fd_sc_hd__a31o_1 _11741_ (.A1(\div_shifter[52] ),
    .A2(net232),
    .A3(_04845_),
    .B1(net192),
    .X(_04847_));
 sky130_fd_sc_hd__nand2_1 _11742_ (.A(_05677_),
    .B(_02319_),
    .Y(_04848_));
 sky130_fd_sc_hd__o211a_1 _11743_ (.A1(_05677_),
    .A2(net196),
    .B1(_04848_),
    .C1(net198),
    .X(_04849_));
 sky130_fd_sc_hd__o22a_1 _11744_ (.A1(_05668_),
    .A2(net209),
    .B1(_04849_),
    .B2(_05687_),
    .X(_04851_));
 sky130_fd_sc_hd__o221a_1 _11745_ (.A1(net177),
    .A2(_03884_),
    .B1(_03896_),
    .B2(_02314_),
    .C1(_04851_),
    .X(_04852_));
 sky130_fd_sc_hd__o21ai_1 _11746_ (.A1(_04846_),
    .A2(_04847_),
    .B1(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__or4_2 _11747_ (.A(_04832_),
    .B(_04840_),
    .C(_04844_),
    .D(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__a221o_1 _11748_ (.A1(_04824_),
    .A2(_04825_),
    .B1(_04827_),
    .B2(_02323_),
    .C1(_04854_),
    .X(_04855_));
 sky130_fd_sc_hd__and3_1 _11749_ (.A(curr_PC[19]),
    .B(curr_PC[20]),
    .C(_04661_),
    .X(_04856_));
 sky130_fd_sc_hd__a21oi_1 _11750_ (.A1(curr_PC[19]),
    .A2(_04661_),
    .B1(curr_PC[20]),
    .Y(_04857_));
 sky130_fd_sc_hd__nor2_1 _11751_ (.A(_04856_),
    .B(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__mux2_8 _11752_ (.A0(_04855_),
    .A1(_04858_),
    .S(net248),
    .X(dest_val[20]));
 sky130_fd_sc_hd__a31o_1 _11753_ (.A1(_04663_),
    .A2(_04725_),
    .A3(_04823_),
    .B1(net158),
    .X(_04859_));
 sky130_fd_sc_hd__o22a_1 _11754_ (.A1(net66),
    .A2(net23),
    .B1(net15),
    .B2(net60),
    .X(_04861_));
 sky130_fd_sc_hd__xnor2_1 _11755_ (.A(net69),
    .B(_04861_),
    .Y(_04862_));
 sky130_fd_sc_hd__o22a_1 _11756_ (.A1(net58),
    .A2(net10),
    .B1(net5),
    .B2(net64),
    .X(_04863_));
 sky130_fd_sc_hd__xnor2_1 _11757_ (.A(net18),
    .B(_04863_),
    .Y(_04864_));
 sky130_fd_sc_hd__a22o_1 _11758_ (.A1(_00143_),
    .A2(net43),
    .B1(net41),
    .B2(_06517_),
    .X(_04865_));
 sky130_fd_sc_hd__xor2_1 _11759_ (.A(net93),
    .B(_04865_),
    .X(_04866_));
 sky130_fd_sc_hd__nand2b_1 _11760_ (.A_N(_04864_),
    .B(_04866_),
    .Y(_04867_));
 sky130_fd_sc_hd__nand2b_1 _11761_ (.A_N(_04866_),
    .B(_04864_),
    .Y(_04868_));
 sky130_fd_sc_hd__nand2_1 _11762_ (.A(_04867_),
    .B(_04868_),
    .Y(_04869_));
 sky130_fd_sc_hd__xor2_1 _11763_ (.A(_04862_),
    .B(_04869_),
    .X(_04870_));
 sky130_fd_sc_hd__and3_1 _11764_ (.A(_00163_),
    .B(net22),
    .C(_04769_),
    .X(_04872_));
 sky130_fd_sc_hd__nand2_1 _11765_ (.A(_04870_),
    .B(_04872_),
    .Y(_04873_));
 sky130_fd_sc_hd__or2_1 _11766_ (.A(_04870_),
    .B(_04872_),
    .X(_04874_));
 sky130_fd_sc_hd__nand2_1 _11767_ (.A(_04873_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__o22a_1 _11768_ (.A1(_00267_),
    .A2(net17),
    .B1(_00699_),
    .B2(_00263_),
    .X(_04876_));
 sky130_fd_sc_hd__xnor2_1 _11769_ (.A(net90),
    .B(_04876_),
    .Y(_04877_));
 sky130_fd_sc_hd__xnor2_1 _11770_ (.A(net50),
    .B(_04877_),
    .Y(_04878_));
 sky130_fd_sc_hd__o22a_1 _11771_ (.A1(net45),
    .A2(net12),
    .B1(net7),
    .B2(net47),
    .X(_04879_));
 sky130_fd_sc_hd__xnor2_1 _11772_ (.A(net95),
    .B(_04879_),
    .Y(_04880_));
 sky130_fd_sc_hd__and2b_1 _11773_ (.A_N(_04878_),
    .B(_04880_),
    .X(_04881_));
 sky130_fd_sc_hd__and2b_1 _11774_ (.A_N(_04880_),
    .B(_04878_),
    .X(_04883_));
 sky130_fd_sc_hd__or2_1 _11775_ (.A(_04881_),
    .B(_04883_),
    .X(_04884_));
 sky130_fd_sc_hd__xor2_1 _11776_ (.A(_04875_),
    .B(_04884_),
    .X(_04885_));
 sky130_fd_sc_hd__o21a_1 _11777_ (.A1(_04775_),
    .A2(_04787_),
    .B1(_04772_),
    .X(_04886_));
 sky130_fd_sc_hd__nor2_1 _11778_ (.A(_04780_),
    .B(_04785_),
    .Y(_04887_));
 sky130_fd_sc_hd__nand2_1 _11779_ (.A(_06547_),
    .B(_02078_),
    .Y(_04888_));
 sky130_fd_sc_hd__nor2_1 _11780_ (.A(_04887_),
    .B(_04888_),
    .Y(_04889_));
 sky130_fd_sc_hd__xnor2_1 _11781_ (.A(_04887_),
    .B(_04888_),
    .Y(_04890_));
 sky130_fd_sc_hd__nor2_1 _11782_ (.A(_04766_),
    .B(_04890_),
    .Y(_04891_));
 sky130_fd_sc_hd__xor2_1 _11783_ (.A(_04766_),
    .B(_04890_),
    .X(_04892_));
 sky130_fd_sc_hd__o21a_1 _11784_ (.A1(_04792_),
    .A2(_04796_),
    .B1(_04892_),
    .X(_04894_));
 sky130_fd_sc_hd__nor3_1 _11785_ (.A(_04792_),
    .B(_04796_),
    .C(_04892_),
    .Y(_04895_));
 sky130_fd_sc_hd__nor2_1 _11786_ (.A(_04894_),
    .B(_04895_),
    .Y(_04896_));
 sky130_fd_sc_hd__and2b_1 _11787_ (.A_N(_04886_),
    .B(_04896_),
    .X(_04897_));
 sky130_fd_sc_hd__xnor2_1 _11788_ (.A(_04886_),
    .B(_04896_),
    .Y(_04898_));
 sky130_fd_sc_hd__nand2_1 _11789_ (.A(_04885_),
    .B(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__or2_1 _11790_ (.A(_04885_),
    .B(_04898_),
    .X(_04900_));
 sky130_fd_sc_hd__and2_1 _11791_ (.A(_04899_),
    .B(_04900_),
    .X(_04901_));
 sky130_fd_sc_hd__o21ai_1 _11792_ (.A1(_04799_),
    .A2(_04802_),
    .B1(_04901_),
    .Y(_04902_));
 sky130_fd_sc_hd__or3_1 _11793_ (.A(_04799_),
    .B(_04802_),
    .C(_04901_),
    .X(_04903_));
 sky130_fd_sc_hd__nand2_1 _11794_ (.A(_04902_),
    .B(_04903_),
    .Y(_04905_));
 sky130_fd_sc_hd__a21oi_1 _11795_ (.A1(_04804_),
    .A2(_04807_),
    .B1(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__a21o_1 _11796_ (.A1(_04804_),
    .A2(_04807_),
    .B1(_04905_),
    .X(_04907_));
 sky130_fd_sc_hd__and3_1 _11797_ (.A(_04804_),
    .B(_04807_),
    .C(_04905_),
    .X(_04908_));
 sky130_fd_sc_hd__or2_4 _11798_ (.A(_04906_),
    .B(_04908_),
    .X(_04909_));
 sky130_fd_sc_hd__nor2_1 _11799_ (.A(_04715_),
    .B(_04813_),
    .Y(_04910_));
 sky130_fd_sc_hd__and2_1 _11800_ (.A(_04716_),
    .B(_04910_),
    .X(_04911_));
 sky130_fd_sc_hd__nand2_1 _11801_ (.A(_04521_),
    .B(_04911_),
    .Y(_04912_));
 sky130_fd_sc_hd__nand2_1 _11802_ (.A(_04524_),
    .B(_04911_),
    .Y(_04913_));
 sky130_fd_sc_hd__a21boi_1 _11803_ (.A1(_04712_),
    .A2(_04811_),
    .B1_N(_04812_),
    .Y(_04914_));
 sky130_fd_sc_hd__a21oi_1 _11804_ (.A1(_04719_),
    .A2(_04910_),
    .B1(_04914_),
    .Y(_04916_));
 sky130_fd_sc_hd__o211a_2 _11805_ (.A1(_04092_),
    .A2(_04912_),
    .B1(_04913_),
    .C1(_04916_),
    .X(_04917_));
 sky130_fd_sc_hd__xnor2_4 _11806_ (.A(_04909_),
    .B(_04917_),
    .Y(_04918_));
 sky130_fd_sc_hd__nor2_1 _11807_ (.A(_04859_),
    .B(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__a21o_1 _11808_ (.A1(_04859_),
    .A2(_04918_),
    .B1(_02242_),
    .X(_04920_));
 sky130_fd_sc_hd__nand2_1 _11809_ (.A(net161),
    .B(_01867_),
    .Y(_04921_));
 sky130_fd_sc_hd__xor2_1 _11810_ (.A(_01868_),
    .B(_04921_),
    .X(_04922_));
 sky130_fd_sc_hd__o21a_1 _11811_ (.A1(_05696_),
    .A2(_06404_),
    .B1(_06406_),
    .X(_04923_));
 sky130_fd_sc_hd__a21bo_1 _11812_ (.A1(_05696_),
    .A2(_04829_),
    .B1_N(_05677_),
    .X(_04924_));
 sky130_fd_sc_hd__mux2_1 _11813_ (.A0(_04923_),
    .A1(_04924_),
    .S(net284),
    .X(_04925_));
 sky130_fd_sc_hd__xnor2_1 _11814_ (.A(_05763_),
    .B(_04925_),
    .Y(_04927_));
 sky130_fd_sc_hd__nand2_1 _11815_ (.A(reg1_val[21]),
    .B(curr_PC[21]),
    .Y(_04928_));
 sky130_fd_sc_hd__or2_1 _11816_ (.A(reg1_val[21]),
    .B(curr_PC[21]),
    .X(_04929_));
 sky130_fd_sc_hd__nand2_1 _11817_ (.A(_04928_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__o21a_1 _11818_ (.A1(_04835_),
    .A2(_04836_),
    .B1(_04833_),
    .X(_04931_));
 sky130_fd_sc_hd__xor2_1 _11819_ (.A(_04930_),
    .B(_04931_),
    .X(_04932_));
 sky130_fd_sc_hd__nor2_1 _11820_ (.A(net229),
    .B(_04932_),
    .Y(_04933_));
 sky130_fd_sc_hd__a211o_1 _11821_ (.A1(net229),
    .A2(_03777_),
    .B1(_04933_),
    .C1(_06476_),
    .X(_04934_));
 sky130_fd_sc_hd__or2_1 _11822_ (.A(\div_shifter[52] ),
    .B(_04845_),
    .X(_04935_));
 sky130_fd_sc_hd__a21oi_1 _11823_ (.A1(net232),
    .A2(_04935_),
    .B1(\div_shifter[53] ),
    .Y(_04936_));
 sky130_fd_sc_hd__a31o_1 _11824_ (.A1(\div_shifter[53] ),
    .A2(net232),
    .A3(_04935_),
    .B1(net192),
    .X(_04938_));
 sky130_fd_sc_hd__or2_1 _11825_ (.A(_04936_),
    .B(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__or2_1 _11826_ (.A(\div_res[20] ),
    .B(_04841_),
    .X(_04940_));
 sky130_fd_sc_hd__a21oi_1 _11827_ (.A1(net165),
    .A2(_04940_),
    .B1(\div_res[21] ),
    .Y(_04941_));
 sky130_fd_sc_hd__a31o_1 _11828_ (.A1(\div_res[21] ),
    .A2(net165),
    .A3(_04940_),
    .B1(net194),
    .X(_04942_));
 sky130_fd_sc_hd__nand2_1 _11829_ (.A(_05744_),
    .B(_02319_),
    .Y(_04943_));
 sky130_fd_sc_hd__o211a_1 _11830_ (.A1(_05744_),
    .A2(net196),
    .B1(_04943_),
    .C1(net198),
    .X(_04944_));
 sky130_fd_sc_hd__o22a_1 _11831_ (.A1(_05725_),
    .A2(net209),
    .B1(_04944_),
    .B2(_05753_),
    .X(_04945_));
 sky130_fd_sc_hd__o221a_1 _11832_ (.A1(net177),
    .A2(_03764_),
    .B1(_03777_),
    .B2(_02314_),
    .C1(_04945_),
    .X(_04946_));
 sky130_fd_sc_hd__o211a_1 _11833_ (.A1(_04941_),
    .A2(_04942_),
    .B1(_04946_),
    .C1(_04939_),
    .X(_04947_));
 sky130_fd_sc_hd__o211a_1 _11834_ (.A1(net236),
    .A2(_04927_),
    .B1(_04934_),
    .C1(_04947_),
    .X(_04949_));
 sky130_fd_sc_hd__o221a_1 _11835_ (.A1(_04919_),
    .A2(_04920_),
    .B1(_04922_),
    .B2(_02324_),
    .C1(_04949_),
    .X(_04950_));
 sky130_fd_sc_hd__nor2_1 _11836_ (.A(curr_PC[21]),
    .B(_04856_),
    .Y(_04951_));
 sky130_fd_sc_hd__and2_1 _11837_ (.A(curr_PC[21]),
    .B(_04856_),
    .X(_04952_));
 sky130_fd_sc_hd__or3_1 _11838_ (.A(net243),
    .B(_04951_),
    .C(_04952_),
    .X(_04953_));
 sky130_fd_sc_hd__o21ai_4 _11839_ (.A1(net248),
    .A2(_04950_),
    .B1(_04953_),
    .Y(dest_val[21]));
 sky130_fd_sc_hd__or4b_1 _11840_ (.A(_04417_),
    .B(_04418_),
    .C(_04527_),
    .D_N(_04628_),
    .X(_04954_));
 sky130_fd_sc_hd__nor4b_2 _11841_ (.A(_04724_),
    .B(_04822_),
    .C(_04954_),
    .D_N(_04918_),
    .Y(_04955_));
 sky130_fd_sc_hd__and2_1 _11842_ (.A(_04347_),
    .B(_04955_),
    .X(_04956_));
 sky130_fd_sc_hd__o22a_1 _11843_ (.A1(net67),
    .A2(net23),
    .B1(net15),
    .B2(net66),
    .X(_04957_));
 sky130_fd_sc_hd__xnor2_1 _11844_ (.A(_00678_),
    .B(_04957_),
    .Y(_04959_));
 sky130_fd_sc_hd__a22oi_1 _11845_ (.A1(_00143_),
    .A2(net41),
    .B1(_00408_),
    .B2(net43),
    .Y(_04960_));
 sky130_fd_sc_hd__xnor2_1 _11846_ (.A(net93),
    .B(_04960_),
    .Y(_04961_));
 sky130_fd_sc_hd__nand2_1 _11847_ (.A(_04959_),
    .B(_04961_),
    .Y(_04962_));
 sky130_fd_sc_hd__or2_1 _11848_ (.A(_04959_),
    .B(_04961_),
    .X(_04963_));
 sky130_fd_sc_hd__nand2_1 _11849_ (.A(_04962_),
    .B(_04963_),
    .Y(_04964_));
 sky130_fd_sc_hd__o21a_1 _11850_ (.A1(_04862_),
    .A2(_04869_),
    .B1(_04867_),
    .X(_04965_));
 sky130_fd_sc_hd__xnor2_1 _11851_ (.A(_04964_),
    .B(_04965_),
    .Y(_04966_));
 sky130_fd_sc_hd__a22o_1 _11852_ (.A1(net38),
    .A2(_00700_),
    .B1(_01951_),
    .B2(net40),
    .X(_04967_));
 sky130_fd_sc_hd__xor2_1 _11853_ (.A(net90),
    .B(_04967_),
    .X(_04968_));
 sky130_fd_sc_hd__or2_1 _11854_ (.A(_00222_),
    .B(net7),
    .X(_04970_));
 sky130_fd_sc_hd__a22o_1 _11855_ (.A1(_00228_),
    .A2(net9),
    .B1(_04970_),
    .B2(net95),
    .X(_04971_));
 sky130_fd_sc_hd__or2_1 _11856_ (.A(_04968_),
    .B(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__nand2_1 _11857_ (.A(_04968_),
    .B(_04971_),
    .Y(_04973_));
 sky130_fd_sc_hd__and2_1 _11858_ (.A(_04972_),
    .B(_04973_),
    .X(_04974_));
 sky130_fd_sc_hd__or2_1 _11859_ (.A(_04966_),
    .B(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__nand2_1 _11860_ (.A(_04966_),
    .B(_04974_),
    .Y(_04976_));
 sky130_fd_sc_hd__nand2_1 _11861_ (.A(_04975_),
    .B(_04976_),
    .Y(_04977_));
 sky130_fd_sc_hd__o21ai_1 _11862_ (.A1(_04875_),
    .A2(_04884_),
    .B1(_04873_),
    .Y(_04978_));
 sky130_fd_sc_hd__a21oi_1 _11863_ (.A1(net50),
    .A2(_04877_),
    .B1(_04881_),
    .Y(_04979_));
 sky130_fd_sc_hd__o22a_1 _11864_ (.A1(net60),
    .A2(net10),
    .B1(net5),
    .B2(net58),
    .X(_04981_));
 sky130_fd_sc_hd__xnor2_1 _11865_ (.A(net18),
    .B(_04981_),
    .Y(_04982_));
 sky130_fd_sc_hd__nor2_1 _11866_ (.A(_04979_),
    .B(_04982_),
    .Y(_04983_));
 sky130_fd_sc_hd__xnor2_1 _11867_ (.A(_04979_),
    .B(_04982_),
    .Y(_04984_));
 sky130_fd_sc_hd__nor2_1 _11868_ (.A(net64),
    .B(net18),
    .Y(_04985_));
 sky130_fd_sc_hd__and2b_1 _11869_ (.A_N(_04984_),
    .B(_04985_),
    .X(_04986_));
 sky130_fd_sc_hd__xnor2_1 _11870_ (.A(_04984_),
    .B(_04985_),
    .Y(_04987_));
 sky130_fd_sc_hd__o21a_1 _11871_ (.A1(_04889_),
    .A2(_04891_),
    .B1(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__nor3_1 _11872_ (.A(_04889_),
    .B(_04891_),
    .C(_04987_),
    .Y(_04989_));
 sky130_fd_sc_hd__nor2_1 _11873_ (.A(_04988_),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__xnor2_1 _11874_ (.A(_04978_),
    .B(_04990_),
    .Y(_04992_));
 sky130_fd_sc_hd__or2_1 _11875_ (.A(_04977_),
    .B(_04992_),
    .X(_04993_));
 sky130_fd_sc_hd__xor2_1 _11876_ (.A(_04977_),
    .B(_04992_),
    .X(_04994_));
 sky130_fd_sc_hd__o21ai_1 _11877_ (.A1(_04894_),
    .A2(_04897_),
    .B1(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hd__or3_1 _11878_ (.A(_04894_),
    .B(_04897_),
    .C(_04994_),
    .X(_04996_));
 sky130_fd_sc_hd__nand2_1 _11879_ (.A(_04995_),
    .B(_04996_),
    .Y(_04997_));
 sky130_fd_sc_hd__a21o_1 _11880_ (.A1(_04899_),
    .A2(_04902_),
    .B1(_04997_),
    .X(_04998_));
 sky130_fd_sc_hd__and3_1 _11881_ (.A(_04899_),
    .B(_04902_),
    .C(_04997_),
    .X(_04999_));
 sky130_fd_sc_hd__inv_2 _11882_ (.A(_04999_),
    .Y(_05000_));
 sky130_fd_sc_hd__nand2_4 _11883_ (.A(_04998_),
    .B(_05000_),
    .Y(_05001_));
 sky130_fd_sc_hd__nor2_2 _11884_ (.A(_04813_),
    .B(_04909_),
    .Y(_05003_));
 sky130_fd_sc_hd__and2_1 _11885_ (.A(_04814_),
    .B(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__inv_2 _11886_ (.A(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__a21oi_2 _11887_ (.A1(_04811_),
    .A2(_04907_),
    .B1(_04908_),
    .Y(_05006_));
 sky130_fd_sc_hd__a221oi_2 _11888_ (.A1(_04818_),
    .A2(_05003_),
    .B1(_05004_),
    .B2(_04625_),
    .C1(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__o31ai_4 _11889_ (.A1(_04201_),
    .A2(_04623_),
    .A3(_05005_),
    .B1(_05007_),
    .Y(_05008_));
 sky130_fd_sc_hd__xor2_4 _11890_ (.A(_05001_),
    .B(_05008_),
    .X(_05009_));
 sky130_fd_sc_hd__o21ai_1 _11891_ (.A1(net160),
    .A2(_04956_),
    .B1(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__or3_1 _11892_ (.A(net160),
    .B(_04956_),
    .C(_05009_),
    .X(_05011_));
 sky130_fd_sc_hd__or2_1 _11893_ (.A(net158),
    .B(_01869_),
    .X(_05012_));
 sky130_fd_sc_hd__a21oi_1 _11894_ (.A1(_01875_),
    .A2(_05012_),
    .B1(_02324_),
    .Y(_05014_));
 sky130_fd_sc_hd__o21a_2 _11895_ (.A1(_01875_),
    .A2(_05012_),
    .B1(_05014_),
    .X(_05015_));
 sky130_fd_sc_hd__a21bo_1 _11896_ (.A1(_05763_),
    .A2(_04924_),
    .B1_N(_05744_),
    .X(_05016_));
 sky130_fd_sc_hd__o21a_1 _11897_ (.A1(_05763_),
    .A2(_04923_),
    .B1(_06405_),
    .X(_05017_));
 sky130_fd_sc_hd__mux2_1 _11898_ (.A0(_05016_),
    .A1(_05017_),
    .S(net295),
    .X(_05018_));
 sky130_fd_sc_hd__o21ai_1 _11899_ (.A1(_05639_),
    .A2(_05018_),
    .B1(_02317_),
    .Y(_05019_));
 sky130_fd_sc_hd__a21oi_1 _11900_ (.A1(_05639_),
    .A2(_05018_),
    .B1(_05019_),
    .Y(_05020_));
 sky130_fd_sc_hd__nand2_1 _11901_ (.A(reg1_val[22]),
    .B(curr_PC[22]),
    .Y(_05021_));
 sky130_fd_sc_hd__or2_1 _11902_ (.A(reg1_val[22]),
    .B(curr_PC[22]),
    .X(_05022_));
 sky130_fd_sc_hd__nand2_1 _11903_ (.A(_05021_),
    .B(_05022_),
    .Y(_05023_));
 sky130_fd_sc_hd__o21a_1 _11904_ (.A1(_04930_),
    .A2(_04931_),
    .B1(_04928_),
    .X(_05025_));
 sky130_fd_sc_hd__xor2_1 _11905_ (.A(_05023_),
    .B(_05025_),
    .X(_05026_));
 sky130_fd_sc_hd__mux2_1 _11906_ (.A0(_03658_),
    .A1(_05026_),
    .S(net250),
    .X(_05027_));
 sky130_fd_sc_hd__or2_1 _11907_ (.A(\div_res[21] ),
    .B(_04940_),
    .X(_05028_));
 sky130_fd_sc_hd__a21oi_1 _11908_ (.A1(net166),
    .A2(_05028_),
    .B1(\div_res[22] ),
    .Y(_05029_));
 sky130_fd_sc_hd__a31o_1 _11909_ (.A1(\div_res[22] ),
    .A2(net166),
    .A3(_05028_),
    .B1(net194),
    .X(_05030_));
 sky130_fd_sc_hd__or2_1 _11910_ (.A(\div_shifter[53] ),
    .B(_04935_),
    .X(_05031_));
 sky130_fd_sc_hd__a21oi_1 _11911_ (.A1(net234),
    .A2(_05031_),
    .B1(\div_shifter[54] ),
    .Y(_05032_));
 sky130_fd_sc_hd__a31o_1 _11912_ (.A1(\div_shifter[54] ),
    .A2(net234),
    .A3(_05031_),
    .B1(net192),
    .X(_05033_));
 sky130_fd_sc_hd__mux2_1 _11913_ (.A0(_02320_),
    .A1(_02326_),
    .S(_05620_),
    .X(_05034_));
 sky130_fd_sc_hd__a21o_1 _11914_ (.A1(net198),
    .A2(_05034_),
    .B1(_05629_),
    .X(_05036_));
 sky130_fd_sc_hd__o21ai_1 _11915_ (.A1(_05609_),
    .A2(net209),
    .B1(_05036_),
    .Y(_05037_));
 sky130_fd_sc_hd__a221o_1 _11916_ (.A1(_02244_),
    .A2(_03646_),
    .B1(_03658_),
    .B2(_02313_),
    .C1(_05037_),
    .X(_05038_));
 sky130_fd_sc_hd__o21ba_1 _11917_ (.A1(_05032_),
    .A2(_05033_),
    .B1_N(_05038_),
    .X(_05039_));
 sky130_fd_sc_hd__o21ai_1 _11918_ (.A1(_05029_),
    .A2(_05030_),
    .B1(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__a211o_1 _11919_ (.A1(net210),
    .A2(_05027_),
    .B1(_05040_),
    .C1(_05020_),
    .X(_05041_));
 sky130_fd_sc_hd__a311o_1 _11920_ (.A1(_02241_),
    .A2(_05010_),
    .A3(_05011_),
    .B1(_05015_),
    .C1(_05041_),
    .X(_05042_));
 sky130_fd_sc_hd__or2_1 _11921_ (.A(curr_PC[22]),
    .B(_04952_),
    .X(_05043_));
 sky130_fd_sc_hd__a21oi_1 _11922_ (.A1(curr_PC[22]),
    .A2(_04952_),
    .B1(net247),
    .Y(_05044_));
 sky130_fd_sc_hd__a22o_4 _11923_ (.A1(net246),
    .A2(_05042_),
    .B1(_05043_),
    .B2(_05044_),
    .X(dest_val[22]));
 sky130_fd_sc_hd__a31o_1 _11924_ (.A1(_04347_),
    .A2(_04955_),
    .A3(_05009_),
    .B1(net160),
    .X(_05046_));
 sky130_fd_sc_hd__a21o_1 _11925_ (.A1(_04978_),
    .A2(_04990_),
    .B1(_04988_),
    .X(_05047_));
 sky130_fd_sc_hd__a22o_1 _11926_ (.A1(net41),
    .A2(_00408_),
    .B1(_00700_),
    .B2(net43),
    .X(_05048_));
 sky130_fd_sc_hd__xor2_1 _11927_ (.A(net93),
    .B(_05048_),
    .X(_05049_));
 sky130_fd_sc_hd__and2b_1 _11928_ (.A_N(net95),
    .B(_05049_),
    .X(_05050_));
 sky130_fd_sc_hd__xor2_1 _11929_ (.A(net95),
    .B(_05049_),
    .X(_05051_));
 sky130_fd_sc_hd__o22a_1 _11930_ (.A1(_00267_),
    .A2(net12),
    .B1(net7),
    .B2(_00263_),
    .X(_05052_));
 sky130_fd_sc_hd__xnor2_1 _11931_ (.A(net90),
    .B(_05052_),
    .Y(_05053_));
 sky130_fd_sc_hd__and2b_1 _11932_ (.A_N(_05051_),
    .B(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__and2b_1 _11933_ (.A_N(_05053_),
    .B(_05051_),
    .X(_05055_));
 sky130_fd_sc_hd__or2_1 _11934_ (.A(_05054_),
    .B(_05055_),
    .X(_05057_));
 sky130_fd_sc_hd__nand2b_1 _11935_ (.A_N(_05057_),
    .B(_04972_),
    .Y(_05058_));
 sky130_fd_sc_hd__nand2b_1 _11936_ (.A_N(_04972_),
    .B(_05057_),
    .Y(_05059_));
 sky130_fd_sc_hd__nand2_1 _11937_ (.A(_05058_),
    .B(_05059_),
    .Y(_05060_));
 sky130_fd_sc_hd__or2_1 _11938_ (.A(_04962_),
    .B(_05060_),
    .X(_05061_));
 sky130_fd_sc_hd__nand2_1 _11939_ (.A(_04962_),
    .B(_05060_),
    .Y(_05062_));
 sky130_fd_sc_hd__and2_1 _11940_ (.A(_05061_),
    .B(_05062_),
    .X(_05063_));
 sky130_fd_sc_hd__o21a_1 _11941_ (.A1(_04964_),
    .A2(_04965_),
    .B1(_04975_),
    .X(_05064_));
 sky130_fd_sc_hd__o22a_1 _11942_ (.A1(net66),
    .A2(net10),
    .B1(net5),
    .B2(net60),
    .X(_05065_));
 sky130_fd_sc_hd__xnor2_1 _11943_ (.A(_02079_),
    .B(_05065_),
    .Y(_05066_));
 sky130_fd_sc_hd__o22a_1 _11944_ (.A1(net55),
    .A2(net23),
    .B1(net15),
    .B2(net67),
    .X(_05068_));
 sky130_fd_sc_hd__xnor2_1 _11945_ (.A(net69),
    .B(_05068_),
    .Y(_05069_));
 sky130_fd_sc_hd__and3b_1 _11946_ (.A_N(_05069_),
    .B(_06563_),
    .C(net22),
    .X(_05070_));
 sky130_fd_sc_hd__o21a_1 _11947_ (.A1(net58),
    .A2(_02079_),
    .B1(_05069_),
    .X(_05071_));
 sky130_fd_sc_hd__nor2_1 _11948_ (.A(_05070_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__and2b_1 _11949_ (.A_N(_05066_),
    .B(_05072_),
    .X(_05073_));
 sky130_fd_sc_hd__xnor2_1 _11950_ (.A(_05066_),
    .B(_05072_),
    .Y(_05074_));
 sky130_fd_sc_hd__o21ai_1 _11951_ (.A1(_04983_),
    .A2(_04986_),
    .B1(_05074_),
    .Y(_05075_));
 sky130_fd_sc_hd__or3_1 _11952_ (.A(_04983_),
    .B(_04986_),
    .C(_05074_),
    .X(_05076_));
 sky130_fd_sc_hd__and2_1 _11953_ (.A(_05075_),
    .B(_05076_),
    .X(_05077_));
 sky130_fd_sc_hd__nand2b_1 _11954_ (.A_N(_05064_),
    .B(_05077_),
    .Y(_05079_));
 sky130_fd_sc_hd__xnor2_1 _11955_ (.A(_05064_),
    .B(_05077_),
    .Y(_05080_));
 sky130_fd_sc_hd__nand2_1 _11956_ (.A(_05063_),
    .B(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__xor2_1 _11957_ (.A(_05063_),
    .B(_05080_),
    .X(_05082_));
 sky130_fd_sc_hd__nand2_1 _11958_ (.A(_05047_),
    .B(_05082_),
    .Y(_05083_));
 sky130_fd_sc_hd__or2_1 _11959_ (.A(_05047_),
    .B(_05082_),
    .X(_05084_));
 sky130_fd_sc_hd__nand2_1 _11960_ (.A(_05083_),
    .B(_05084_),
    .Y(_05085_));
 sky130_fd_sc_hd__a21o_1 _11961_ (.A1(_04993_),
    .A2(_04995_),
    .B1(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__and3_1 _11962_ (.A(_04993_),
    .B(_04995_),
    .C(_05085_),
    .X(_05087_));
 sky130_fd_sc_hd__inv_2 _11963_ (.A(_05087_),
    .Y(_05088_));
 sky130_fd_sc_hd__nand2_2 _11964_ (.A(_05086_),
    .B(_05088_),
    .Y(_05090_));
 sky130_fd_sc_hd__nor2_1 _11965_ (.A(_04909_),
    .B(_05001_),
    .Y(_05091_));
 sky130_fd_sc_hd__nand2_1 _11966_ (.A(_04910_),
    .B(_05091_),
    .Y(_05092_));
 sky130_fd_sc_hd__inv_2 _11967_ (.A(_05092_),
    .Y(_05093_));
 sky130_fd_sc_hd__nor2_1 _11968_ (.A(_04717_),
    .B(_05092_),
    .Y(_05094_));
 sky130_fd_sc_hd__a21oi_2 _11969_ (.A1(_04907_),
    .A2(_04998_),
    .B1(_04999_),
    .Y(_05095_));
 sky130_fd_sc_hd__a21o_1 _11970_ (.A1(_04914_),
    .A2(_05091_),
    .B1(_05095_),
    .X(_05096_));
 sky130_fd_sc_hd__a221o_2 _11971_ (.A1(_04720_),
    .A2(_05093_),
    .B1(_05094_),
    .B2(_04308_),
    .C1(_05096_),
    .X(_05097_));
 sky130_fd_sc_hd__xor2_2 _11972_ (.A(_05090_),
    .B(_05097_),
    .X(_05098_));
 sky130_fd_sc_hd__nor2_1 _11973_ (.A(_05046_),
    .B(_05098_),
    .Y(_05099_));
 sky130_fd_sc_hd__a21o_1 _11974_ (.A1(_05046_),
    .A2(_05098_),
    .B1(_02242_),
    .X(_05101_));
 sky130_fd_sc_hd__a21oi_1 _11975_ (.A1(net161),
    .A2(_01876_),
    .B1(_01878_),
    .Y(_05102_));
 sky130_fd_sc_hd__a31o_1 _11976_ (.A1(net161),
    .A2(_01876_),
    .A3(_01878_),
    .B1(_02324_),
    .X(_05103_));
 sky130_fd_sc_hd__or2_2 _11977_ (.A(_05102_),
    .B(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__o211a_1 _11978_ (.A1(_05639_),
    .A2(_05017_),
    .B1(_06409_),
    .C1(net295),
    .X(_05105_));
 sky130_fd_sc_hd__a21o_1 _11979_ (.A1(_05639_),
    .A2(_05016_),
    .B1(_05620_),
    .X(_05106_));
 sky130_fd_sc_hd__a21o_1 _11980_ (.A1(net284),
    .A2(_05106_),
    .B1(_05105_),
    .X(_05107_));
 sky130_fd_sc_hd__o21ai_1 _11981_ (.A1(_05577_),
    .A2(_05107_),
    .B1(_02317_),
    .Y(_05108_));
 sky130_fd_sc_hd__a21o_1 _11982_ (.A1(_05577_),
    .A2(_05107_),
    .B1(_05108_),
    .X(_05109_));
 sky130_fd_sc_hd__nand2_1 _11983_ (.A(reg1_val[23]),
    .B(curr_PC[23]),
    .Y(_05110_));
 sky130_fd_sc_hd__or2_1 _11984_ (.A(reg1_val[23]),
    .B(curr_PC[23]),
    .X(_05112_));
 sky130_fd_sc_hd__nand2_1 _11985_ (.A(_05110_),
    .B(_05112_),
    .Y(_05113_));
 sky130_fd_sc_hd__o21a_1 _11986_ (.A1(_05023_),
    .A2(_05025_),
    .B1(_05021_),
    .X(_05114_));
 sky130_fd_sc_hd__xnor2_1 _11987_ (.A(_05113_),
    .B(_05114_),
    .Y(_05115_));
 sky130_fd_sc_hd__mux2_1 _11988_ (.A0(_03528_),
    .A1(_05115_),
    .S(net250),
    .X(_05116_));
 sky130_fd_sc_hd__or2_1 _11989_ (.A(\div_res[22] ),
    .B(_05028_),
    .X(_05117_));
 sky130_fd_sc_hd__a21oi_1 _11990_ (.A1(net165),
    .A2(_05117_),
    .B1(\div_res[23] ),
    .Y(_05118_));
 sky130_fd_sc_hd__a31o_1 _11991_ (.A1(\div_res[23] ),
    .A2(net166),
    .A3(_05117_),
    .B1(net195),
    .X(_05119_));
 sky130_fd_sc_hd__or2_1 _11992_ (.A(\div_shifter[54] ),
    .B(_05031_),
    .X(_05120_));
 sky130_fd_sc_hd__a21oi_1 _11993_ (.A1(net232),
    .A2(_05120_),
    .B1(\div_shifter[55] ),
    .Y(_05121_));
 sky130_fd_sc_hd__a311o_1 _11994_ (.A1(\div_shifter[55] ),
    .A2(net234),
    .A3(_05120_),
    .B1(_05121_),
    .C1(net192),
    .X(_05123_));
 sky130_fd_sc_hd__nand2_1 _11995_ (.A(_05555_),
    .B(_02325_),
    .Y(_05124_));
 sky130_fd_sc_hd__o211a_1 _11996_ (.A1(_05555_),
    .A2(_02320_),
    .B1(_05124_),
    .C1(net198),
    .X(_05125_));
 sky130_fd_sc_hd__o22a_1 _11997_ (.A1(_05544_),
    .A2(net209),
    .B1(_05125_),
    .B2(_05566_),
    .X(_05126_));
 sky130_fd_sc_hd__o221a_1 _11998_ (.A1(net177),
    .A2(_03516_),
    .B1(_03528_),
    .B2(_02314_),
    .C1(_05126_),
    .X(_05127_));
 sky130_fd_sc_hd__o211a_1 _11999_ (.A1(_05118_),
    .A2(_05119_),
    .B1(_05123_),
    .C1(_05127_),
    .X(_05128_));
 sky130_fd_sc_hd__o211a_1 _12000_ (.A1(_06476_),
    .A2(_05116_),
    .B1(_05128_),
    .C1(_05109_),
    .X(_05129_));
 sky130_fd_sc_hd__o211a_1 _12001_ (.A1(_05099_),
    .A2(_05101_),
    .B1(_05104_),
    .C1(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__a21oi_1 _12002_ (.A1(curr_PC[22]),
    .A2(_04952_),
    .B1(curr_PC[23]),
    .Y(_05131_));
 sky130_fd_sc_hd__and3_1 _12003_ (.A(curr_PC[22]),
    .B(curr_PC[23]),
    .C(_04952_),
    .X(_05132_));
 sky130_fd_sc_hd__or3_1 _12004_ (.A(net246),
    .B(_05131_),
    .C(_05132_),
    .X(_05134_));
 sky130_fd_sc_hd__o21ai_4 _12005_ (.A1(_06457_),
    .A2(_05130_),
    .B1(_05134_),
    .Y(dest_val[23]));
 sky130_fd_sc_hd__o31a_1 _12006_ (.A1(net95),
    .A2(_00259_),
    .A3(net8),
    .B1(net90),
    .X(_05135_));
 sky130_fd_sc_hd__nor2_1 _12007_ (.A(net90),
    .B(net7),
    .Y(_05136_));
 sky130_fd_sc_hd__a21o_2 _12008_ (.A1(_00260_),
    .A2(_05136_),
    .B1(_05135_),
    .X(_05137_));
 sky130_fd_sc_hd__nor2_1 _12009_ (.A(net60),
    .B(_02079_),
    .Y(_05138_));
 sky130_fd_sc_hd__xnor2_1 _12010_ (.A(_05137_),
    .B(_05138_),
    .Y(_05139_));
 sky130_fd_sc_hd__o21ai_1 _12011_ (.A1(_05050_),
    .A2(_05054_),
    .B1(_05139_),
    .Y(_05140_));
 sky130_fd_sc_hd__or3_1 _12012_ (.A(_05050_),
    .B(_05054_),
    .C(_05139_),
    .X(_05141_));
 sky130_fd_sc_hd__and2_1 _12013_ (.A(_05140_),
    .B(_05141_),
    .X(_05142_));
 sky130_fd_sc_hd__o22a_1 _12014_ (.A1(net17),
    .A2(net23),
    .B1(net15),
    .B2(net55),
    .X(_05144_));
 sky130_fd_sc_hd__xnor2_1 _12015_ (.A(net69),
    .B(_05144_),
    .Y(_05145_));
 sky130_fd_sc_hd__o22a_1 _12016_ (.A1(net68),
    .A2(net10),
    .B1(net5),
    .B2(net66),
    .X(_05146_));
 sky130_fd_sc_hd__xnor2_1 _12017_ (.A(net20),
    .B(_05146_),
    .Y(_05147_));
 sky130_fd_sc_hd__a22o_1 _12018_ (.A1(net41),
    .A2(_00700_),
    .B1(_01951_),
    .B2(net43),
    .X(_05148_));
 sky130_fd_sc_hd__xnor2_1 _12019_ (.A(net93),
    .B(_05148_),
    .Y(_05149_));
 sky130_fd_sc_hd__nor2_1 _12020_ (.A(_05147_),
    .B(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__and2_1 _12021_ (.A(_05147_),
    .B(_05149_),
    .X(_05151_));
 sky130_fd_sc_hd__or2_1 _12022_ (.A(_05150_),
    .B(_05151_),
    .X(_05152_));
 sky130_fd_sc_hd__nor2_1 _12023_ (.A(_05145_),
    .B(_05152_),
    .Y(_05153_));
 sky130_fd_sc_hd__and2_1 _12024_ (.A(_05145_),
    .B(_05152_),
    .X(_05155_));
 sky130_fd_sc_hd__nor2_1 _12025_ (.A(_05153_),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__o21ai_1 _12026_ (.A1(_05070_),
    .A2(_05073_),
    .B1(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__or3_1 _12027_ (.A(_05070_),
    .B(_05073_),
    .C(_05156_),
    .X(_05158_));
 sky130_fd_sc_hd__nand2_1 _12028_ (.A(_05157_),
    .B(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__a21o_1 _12029_ (.A1(_05058_),
    .A2(_05061_),
    .B1(_05159_),
    .X(_05160_));
 sky130_fd_sc_hd__nand3_1 _12030_ (.A(_05058_),
    .B(_05061_),
    .C(_05159_),
    .Y(_05161_));
 sky130_fd_sc_hd__and2_1 _12031_ (.A(_05160_),
    .B(_05161_),
    .X(_05162_));
 sky130_fd_sc_hd__nand2_1 _12032_ (.A(_05142_),
    .B(_05162_),
    .Y(_05163_));
 sky130_fd_sc_hd__or2_1 _12033_ (.A(_05142_),
    .B(_05162_),
    .X(_05164_));
 sky130_fd_sc_hd__nand2_1 _12034_ (.A(_05163_),
    .B(_05164_),
    .Y(_05166_));
 sky130_fd_sc_hd__a21o_1 _12035_ (.A1(_05075_),
    .A2(_05079_),
    .B1(_05166_),
    .X(_05167_));
 sky130_fd_sc_hd__nand3_1 _12036_ (.A(_05075_),
    .B(_05079_),
    .C(_05166_),
    .Y(_05168_));
 sky130_fd_sc_hd__nand2_1 _12037_ (.A(_05167_),
    .B(_05168_),
    .Y(_05169_));
 sky130_fd_sc_hd__a21oi_2 _12038_ (.A1(_05081_),
    .A2(_05083_),
    .B1(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__inv_2 _12039_ (.A(_05170_),
    .Y(_05171_));
 sky130_fd_sc_hd__and3_1 _12040_ (.A(_05081_),
    .B(_05083_),
    .C(_05169_),
    .X(_05172_));
 sky130_fd_sc_hd__or2_2 _12041_ (.A(_05170_),
    .B(_05172_),
    .X(_05173_));
 sky130_fd_sc_hd__nor2_2 _12042_ (.A(_05001_),
    .B(_05090_),
    .Y(_05174_));
 sky130_fd_sc_hd__nand2_1 _12043_ (.A(_05003_),
    .B(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hd__a21oi_1 _12044_ (.A1(_04998_),
    .A2(_05086_),
    .B1(_05087_),
    .Y(_05177_));
 sky130_fd_sc_hd__a21o_1 _12045_ (.A1(_05006_),
    .A2(_05174_),
    .B1(_05177_),
    .X(_05178_));
 sky130_fd_sc_hd__a31o_1 _12046_ (.A1(_04819_),
    .A2(_05003_),
    .A3(_05174_),
    .B1(_05178_),
    .X(_05179_));
 sky130_fd_sc_hd__a41o_1 _12047_ (.A1(_04416_),
    .A2(_04816_),
    .A3(_05003_),
    .A4(_05174_),
    .B1(_05179_),
    .X(_05180_));
 sky130_fd_sc_hd__xor2_2 _12048_ (.A(_05173_),
    .B(_05180_),
    .X(_05181_));
 sky130_fd_sc_hd__and2_1 _12049_ (.A(_05009_),
    .B(_05098_),
    .X(_05182_));
 sky130_fd_sc_hd__and3_2 _12050_ (.A(_04347_),
    .B(_04955_),
    .C(_05182_),
    .X(_05183_));
 sky130_fd_sc_hd__o21ai_1 _12051_ (.A1(net160),
    .A2(_05183_),
    .B1(_05181_),
    .Y(_05184_));
 sky130_fd_sc_hd__o31a_1 _12052_ (.A1(net160),
    .A2(_05181_),
    .A3(_05183_),
    .B1(_02241_),
    .X(_05185_));
 sky130_fd_sc_hd__a21oi_1 _12053_ (.A1(_05577_),
    .A2(_05106_),
    .B1(_05555_),
    .Y(_05186_));
 sky130_fd_sc_hd__mux2_1 _12054_ (.A0(_06412_),
    .A1(_05186_),
    .S(net285),
    .X(_05188_));
 sky130_fd_sc_hd__a21oi_1 _12055_ (.A1(_05350_),
    .A2(_05188_),
    .B1(net236),
    .Y(_05189_));
 sky130_fd_sc_hd__o21a_1 _12056_ (.A1(_05350_),
    .A2(_05188_),
    .B1(_05189_),
    .X(_05190_));
 sky130_fd_sc_hd__a21oi_1 _12057_ (.A1(net163),
    .A2(_01879_),
    .B1(_01886_),
    .Y(_05191_));
 sky130_fd_sc_hd__a311oi_4 _12058_ (.A1(net163),
    .A2(_01879_),
    .A3(_01886_),
    .B1(_02324_),
    .C1(_05191_),
    .Y(_05192_));
 sky130_fd_sc_hd__o21a_1 _12059_ (.A1(_05113_),
    .A2(_05114_),
    .B1(_05110_),
    .X(_05193_));
 sky130_fd_sc_hd__nor2_1 _12060_ (.A(reg1_val[24]),
    .B(curr_PC[24]),
    .Y(_05194_));
 sky130_fd_sc_hd__nand2_1 _12061_ (.A(reg1_val[24]),
    .B(curr_PC[24]),
    .Y(_05195_));
 sky130_fd_sc_hd__and2b_1 _12062_ (.A_N(_05194_),
    .B(_05195_),
    .X(_05196_));
 sky130_fd_sc_hd__xnor2_1 _12063_ (.A(_05193_),
    .B(_05196_),
    .Y(_05197_));
 sky130_fd_sc_hd__mux2_1 _12064_ (.A0(_03378_),
    .A1(_05197_),
    .S(net249),
    .X(_05199_));
 sky130_fd_sc_hd__or2_1 _12065_ (.A(\div_res[23] ),
    .B(_05117_),
    .X(_05200_));
 sky130_fd_sc_hd__a21oi_1 _12066_ (.A1(net167),
    .A2(_05200_),
    .B1(\div_res[24] ),
    .Y(_05201_));
 sky130_fd_sc_hd__a31o_1 _12067_ (.A1(\div_res[24] ),
    .A2(net167),
    .A3(_05200_),
    .B1(net194),
    .X(_05202_));
 sky130_fd_sc_hd__or2_1 _12068_ (.A(\div_shifter[55] ),
    .B(_05120_),
    .X(_05203_));
 sky130_fd_sc_hd__a21oi_1 _12069_ (.A1(net233),
    .A2(_05203_),
    .B1(\div_shifter[56] ),
    .Y(_05204_));
 sky130_fd_sc_hd__a311o_1 _12070_ (.A1(\div_shifter[56] ),
    .A2(net233),
    .A3(_05203_),
    .B1(_05204_),
    .C1(net192),
    .X(_05205_));
 sky130_fd_sc_hd__mux2_1 _12071_ (.A0(_02325_),
    .A1(_02319_),
    .S(_05328_),
    .X(_05206_));
 sky130_fd_sc_hd__o21a_1 _12072_ (.A1(_02315_),
    .A2(_05206_),
    .B1(_05339_),
    .X(_05207_));
 sky130_fd_sc_hd__a221o_1 _12073_ (.A1(_05317_),
    .A2(net241),
    .B1(_02313_),
    .B2(_03378_),
    .C1(_05207_),
    .X(_05208_));
 sky130_fd_sc_hd__a21oi_1 _12074_ (.A1(net179),
    .A2(_03384_),
    .B1(_05208_),
    .Y(_05210_));
 sky130_fd_sc_hd__o211ai_1 _12075_ (.A1(_05201_),
    .A2(_05202_),
    .B1(_05205_),
    .C1(_05210_),
    .Y(_05211_));
 sky130_fd_sc_hd__a211o_1 _12076_ (.A1(_06475_),
    .A2(_05199_),
    .B1(_05211_),
    .C1(_05192_),
    .X(_05212_));
 sky130_fd_sc_hd__a211o_1 _12077_ (.A1(_05184_),
    .A2(_05185_),
    .B1(_05190_),
    .C1(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__or2_1 _12078_ (.A(curr_PC[24]),
    .B(_05132_),
    .X(_05214_));
 sky130_fd_sc_hd__and2_1 _12079_ (.A(curr_PC[24]),
    .B(_05132_),
    .X(_05215_));
 sky130_fd_sc_hd__nor2_1 _12080_ (.A(net246),
    .B(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__a22o_4 _12081_ (.A1(net246),
    .A2(_05213_),
    .B1(_05214_),
    .B2(_05216_),
    .X(dest_val[24]));
 sky130_fd_sc_hd__o22a_1 _12082_ (.A1(net55),
    .A2(net10),
    .B1(net5),
    .B2(net67),
    .X(_05217_));
 sky130_fd_sc_hd__xnor2_1 _12083_ (.A(net19),
    .B(_05217_),
    .Y(_05218_));
 sky130_fd_sc_hd__nand2b_1 _12084_ (.A_N(_05218_),
    .B(_05137_),
    .Y(_05220_));
 sky130_fd_sc_hd__nand2b_1 _12085_ (.A_N(_05137_),
    .B(_05218_),
    .Y(_05221_));
 sky130_fd_sc_hd__nand2_1 _12086_ (.A(_05220_),
    .B(_05221_),
    .Y(_05222_));
 sky130_fd_sc_hd__nor2_1 _12087_ (.A(net66),
    .B(net19),
    .Y(_05223_));
 sky130_fd_sc_hd__xnor2_1 _12088_ (.A(_05222_),
    .B(_05223_),
    .Y(_05224_));
 sky130_fd_sc_hd__o31ai_2 _12089_ (.A1(net60),
    .A2(net18),
    .A3(_05137_),
    .B1(_05140_),
    .Y(_05225_));
 sky130_fd_sc_hd__o22a_1 _12090_ (.A1(net17),
    .A2(net15),
    .B1(_00699_),
    .B2(net23),
    .X(_05226_));
 sky130_fd_sc_hd__xnor2_1 _12091_ (.A(net70),
    .B(_05226_),
    .Y(_05227_));
 sky130_fd_sc_hd__or2_1 _12092_ (.A(net90),
    .B(_05227_),
    .X(_05228_));
 sky130_fd_sc_hd__nand2_1 _12093_ (.A(net90),
    .B(_05227_),
    .Y(_05229_));
 sky130_fd_sc_hd__and2_1 _12094_ (.A(_05228_),
    .B(_05229_),
    .X(_05231_));
 sky130_fd_sc_hd__a22o_1 _12095_ (.A1(net41),
    .A2(_01951_),
    .B1(_02066_),
    .B2(net43),
    .X(_05232_));
 sky130_fd_sc_hd__xor2_1 _12096_ (.A(net93),
    .B(_05232_),
    .X(_05233_));
 sky130_fd_sc_hd__nand2_1 _12097_ (.A(_05231_),
    .B(_05233_),
    .Y(_05234_));
 sky130_fd_sc_hd__or2_1 _12098_ (.A(_05231_),
    .B(_05233_),
    .X(_05235_));
 sky130_fd_sc_hd__and2_1 _12099_ (.A(_05234_),
    .B(_05235_),
    .X(_05236_));
 sky130_fd_sc_hd__o21a_1 _12100_ (.A1(_05150_),
    .A2(_05153_),
    .B1(_05236_),
    .X(_05237_));
 sky130_fd_sc_hd__nor3_1 _12101_ (.A(_05150_),
    .B(_05153_),
    .C(_05236_),
    .Y(_05238_));
 sky130_fd_sc_hd__nor2_1 _12102_ (.A(_05237_),
    .B(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__xor2_1 _12103_ (.A(_05225_),
    .B(_05239_),
    .X(_05240_));
 sky130_fd_sc_hd__nand2_1 _12104_ (.A(_05224_),
    .B(_05240_),
    .Y(_05242_));
 sky130_fd_sc_hd__or2_1 _12105_ (.A(_05224_),
    .B(_05240_),
    .X(_05243_));
 sky130_fd_sc_hd__nand2_1 _12106_ (.A(_05242_),
    .B(_05243_),
    .Y(_05244_));
 sky130_fd_sc_hd__a21o_1 _12107_ (.A1(_05157_),
    .A2(_05160_),
    .B1(_05244_),
    .X(_05245_));
 sky130_fd_sc_hd__nand3_1 _12108_ (.A(_05157_),
    .B(_05160_),
    .C(_05244_),
    .Y(_05246_));
 sky130_fd_sc_hd__nand2_1 _12109_ (.A(_05245_),
    .B(_05246_),
    .Y(_05247_));
 sky130_fd_sc_hd__a21oi_1 _12110_ (.A1(_05163_),
    .A2(_05167_),
    .B1(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__nand3_1 _12111_ (.A(_05163_),
    .B(_05167_),
    .C(_05247_),
    .Y(_05249_));
 sky130_fd_sc_hd__nand2b_2 _12112_ (.A_N(_05248_),
    .B(_05249_),
    .Y(_05250_));
 sky130_fd_sc_hd__nor2_1 _12113_ (.A(_05090_),
    .B(_05173_),
    .Y(_05251_));
 sky130_fd_sc_hd__nand2_1 _12114_ (.A(_05091_),
    .B(_05251_),
    .Y(_05253_));
 sky130_fd_sc_hd__inv_2 _12115_ (.A(_05253_),
    .Y(_05254_));
 sky130_fd_sc_hd__a21oi_1 _12116_ (.A1(_05086_),
    .A2(_05171_),
    .B1(_05172_),
    .Y(_05255_));
 sky130_fd_sc_hd__a21oi_1 _12117_ (.A1(_05095_),
    .A2(_05251_),
    .B1(_05255_),
    .Y(_05256_));
 sky130_fd_sc_hd__o21ai_1 _12118_ (.A1(_04916_),
    .A2(_05253_),
    .B1(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__a31o_1 _12119_ (.A1(_04526_),
    .A2(_04911_),
    .A3(_05254_),
    .B1(_05257_),
    .X(_05258_));
 sky130_fd_sc_hd__xor2_2 _12120_ (.A(_05250_),
    .B(_05258_),
    .X(_05259_));
 sky130_fd_sc_hd__a21o_1 _12121_ (.A1(_05181_),
    .A2(_05183_),
    .B1(net160),
    .X(_05260_));
 sky130_fd_sc_hd__nand2_1 _12122_ (.A(_05259_),
    .B(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__or2_1 _12123_ (.A(_05259_),
    .B(_05260_),
    .X(_05262_));
 sky130_fd_sc_hd__o21a_1 _12124_ (.A1(_05350_),
    .A2(_05186_),
    .B1(_05328_),
    .X(_05264_));
 sky130_fd_sc_hd__mux2_1 _12125_ (.A0(_06430_),
    .A1(_05264_),
    .S(net286),
    .X(_05265_));
 sky130_fd_sc_hd__a21oi_1 _12126_ (.A1(_05274_),
    .A2(_05265_),
    .B1(net236),
    .Y(_05266_));
 sky130_fd_sc_hd__o21a_1 _12127_ (.A1(_05274_),
    .A2(_05265_),
    .B1(_05266_),
    .X(_05267_));
 sky130_fd_sc_hd__o21ai_1 _12128_ (.A1(net159),
    .A2(_01887_),
    .B1(_01803_),
    .Y(_05268_));
 sky130_fd_sc_hd__or3_1 _12129_ (.A(net159),
    .B(_01803_),
    .C(_01887_),
    .X(_05269_));
 sky130_fd_sc_hd__o21a_1 _12130_ (.A1(_05193_),
    .A2(_05194_),
    .B1(_05195_),
    .X(_05270_));
 sky130_fd_sc_hd__nor2_1 _12131_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .Y(_05271_));
 sky130_fd_sc_hd__nand2_1 _12132_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .Y(_05272_));
 sky130_fd_sc_hd__nand2b_1 _12133_ (.A_N(_05271_),
    .B(_05272_),
    .Y(_05273_));
 sky130_fd_sc_hd__xnor2_1 _12134_ (.A(_05270_),
    .B(_05273_),
    .Y(_05275_));
 sky130_fd_sc_hd__mux2_1 _12135_ (.A0(_03244_),
    .A1(_05275_),
    .S(net250),
    .X(_05276_));
 sky130_fd_sc_hd__or2_1 _12136_ (.A(\div_shifter[56] ),
    .B(_05203_),
    .X(_05277_));
 sky130_fd_sc_hd__a21oi_1 _12137_ (.A1(net233),
    .A2(_05277_),
    .B1(\div_shifter[57] ),
    .Y(_05278_));
 sky130_fd_sc_hd__a31o_1 _12138_ (.A1(\div_shifter[57] ),
    .A2(net233),
    .A3(_05277_),
    .B1(net193),
    .X(_05279_));
 sky130_fd_sc_hd__or2_1 _12139_ (.A(_05278_),
    .B(_05279_),
    .X(_05280_));
 sky130_fd_sc_hd__or2_1 _12140_ (.A(\div_res[24] ),
    .B(_05200_),
    .X(_05281_));
 sky130_fd_sc_hd__a21oi_1 _12141_ (.A1(net166),
    .A2(_05281_),
    .B1(\div_res[25] ),
    .Y(_05282_));
 sky130_fd_sc_hd__a31o_1 _12142_ (.A1(\div_res[25] ),
    .A2(net166),
    .A3(_05281_),
    .B1(net195),
    .X(_05283_));
 sky130_fd_sc_hd__mux2_1 _12143_ (.A0(_02320_),
    .A1(_02326_),
    .S(_05252_),
    .X(_05284_));
 sky130_fd_sc_hd__a21o_1 _12144_ (.A1(net199),
    .A2(_05284_),
    .B1(_05263_),
    .X(_05286_));
 sky130_fd_sc_hd__o221a_1 _12145_ (.A1(_05241_),
    .A2(net209),
    .B1(_02314_),
    .B2(_03244_),
    .C1(_05286_),
    .X(_05287_));
 sky130_fd_sc_hd__a21boi_1 _12146_ (.A1(net179),
    .A2(_03251_),
    .B1_N(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__o211a_1 _12147_ (.A1(_05282_),
    .A2(_05283_),
    .B1(_05288_),
    .C1(_05280_),
    .X(_05289_));
 sky130_fd_sc_hd__o21ai_2 _12148_ (.A1(_06476_),
    .A2(_05276_),
    .B1(_05289_),
    .Y(_05290_));
 sky130_fd_sc_hd__a31o_1 _12149_ (.A1(_02323_),
    .A2(_05268_),
    .A3(_05269_),
    .B1(_05290_),
    .X(_05291_));
 sky130_fd_sc_hd__a311o_1 _12150_ (.A1(_02241_),
    .A2(_05261_),
    .A3(_05262_),
    .B1(_05267_),
    .C1(_05291_),
    .X(_05292_));
 sky130_fd_sc_hd__nor2_1 _12151_ (.A(curr_PC[25]),
    .B(_05215_),
    .Y(_05293_));
 sky130_fd_sc_hd__a31o_1 _12152_ (.A1(curr_PC[24]),
    .A2(curr_PC[25]),
    .A3(_05132_),
    .B1(net246),
    .X(_05294_));
 sky130_fd_sc_hd__a2bb2o_4 _12153_ (.A1_N(_05293_),
    .A2_N(_05294_),
    .B1(net246),
    .B2(_05292_),
    .X(dest_val[25]));
 sky130_fd_sc_hd__a21o_1 _12154_ (.A1(_05225_),
    .A2(_05239_),
    .B1(_05237_),
    .X(_05296_));
 sky130_fd_sc_hd__a21bo_1 _12155_ (.A1(_05221_),
    .A2(_05223_),
    .B1_N(_05220_),
    .X(_05297_));
 sky130_fd_sc_hd__o22a_1 _12156_ (.A1(net15),
    .A2(_00699_),
    .B1(net12),
    .B2(net23),
    .X(_05298_));
 sky130_fd_sc_hd__xnor2_1 _12157_ (.A(net70),
    .B(_05298_),
    .Y(_05299_));
 sky130_fd_sc_hd__nand2_1 _12158_ (.A(_00248_),
    .B(net9),
    .Y(_05300_));
 sky130_fd_sc_hd__a22o_1 _12159_ (.A1(_00250_),
    .A2(net9),
    .B1(_05300_),
    .B2(net92),
    .X(_05301_));
 sky130_fd_sc_hd__and2b_1 _12160_ (.A_N(_05301_),
    .B(_05299_),
    .X(_05302_));
 sky130_fd_sc_hd__and2b_1 _12161_ (.A_N(_05299_),
    .B(_05301_),
    .X(_05303_));
 sky130_fd_sc_hd__nor2_1 _12162_ (.A(_05302_),
    .B(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__a21oi_1 _12163_ (.A1(_05228_),
    .A2(_05234_),
    .B1(_05304_),
    .Y(_05305_));
 sky130_fd_sc_hd__and3_1 _12164_ (.A(_05228_),
    .B(_05234_),
    .C(_05304_),
    .X(_05307_));
 sky130_fd_sc_hd__nor2_1 _12165_ (.A(_05305_),
    .B(_05307_),
    .Y(_05308_));
 sky130_fd_sc_hd__and2_1 _12166_ (.A(_05297_),
    .B(_05308_),
    .X(_05309_));
 sky130_fd_sc_hd__xnor2_1 _12167_ (.A(_05297_),
    .B(_05308_),
    .Y(_05310_));
 sky130_fd_sc_hd__a22o_1 _12168_ (.A1(_00408_),
    .A2(_01967_),
    .B1(_02082_),
    .B2(_00143_),
    .X(_05311_));
 sky130_fd_sc_hd__nor2_1 _12169_ (.A(_06517_),
    .B(net18),
    .Y(_05312_));
 sky130_fd_sc_hd__xnor2_1 _12170_ (.A(_05311_),
    .B(_05312_),
    .Y(_05313_));
 sky130_fd_sc_hd__nor2_1 _12171_ (.A(_05310_),
    .B(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__and2_1 _12172_ (.A(_05310_),
    .B(_05313_),
    .X(_05315_));
 sky130_fd_sc_hd__or2_1 _12173_ (.A(_05314_),
    .B(_05315_),
    .X(_05316_));
 sky130_fd_sc_hd__and2b_1 _12174_ (.A_N(_05316_),
    .B(_05296_),
    .X(_05318_));
 sky130_fd_sc_hd__xor2_1 _12175_ (.A(_05296_),
    .B(_05316_),
    .X(_05319_));
 sky130_fd_sc_hd__a21oi_1 _12176_ (.A1(_05242_),
    .A2(_05245_),
    .B1(_05319_),
    .Y(_05320_));
 sky130_fd_sc_hd__and3_1 _12177_ (.A(_05242_),
    .B(_05245_),
    .C(_05319_),
    .X(_05321_));
 sky130_fd_sc_hd__or2_2 _12178_ (.A(_05320_),
    .B(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__nor2_1 _12179_ (.A(_05173_),
    .B(_05250_),
    .Y(_05323_));
 sky130_fd_sc_hd__o21ai_1 _12180_ (.A1(_05170_),
    .A2(_05248_),
    .B1(_05249_),
    .Y(_05324_));
 sky130_fd_sc_hd__a21bo_1 _12181_ (.A1(_05177_),
    .A2(_05323_),
    .B1_N(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__a31oi_4 _12182_ (.A1(_05008_),
    .A2(_05174_),
    .A3(_05323_),
    .B1(_05325_),
    .Y(_05326_));
 sky130_fd_sc_hd__xnor2_2 _12183_ (.A(_05322_),
    .B(_05326_),
    .Y(_05327_));
 sky130_fd_sc_hd__and2_1 _12184_ (.A(_05181_),
    .B(_05259_),
    .X(_05329_));
 sky130_fd_sc_hd__a41o_1 _12185_ (.A1(_04347_),
    .A2(_04955_),
    .A3(_05182_),
    .A4(_05329_),
    .B1(net160),
    .X(_05330_));
 sky130_fd_sc_hd__a21oi_1 _12186_ (.A1(_05327_),
    .A2(_05330_),
    .B1(_02242_),
    .Y(_05331_));
 sky130_fd_sc_hd__o21a_1 _12187_ (.A1(_05327_),
    .A2(_05330_),
    .B1(_05331_),
    .X(_05332_));
 sky130_fd_sc_hd__o21ba_1 _12188_ (.A1(_05274_),
    .A2(_05264_),
    .B1_N(_05252_),
    .X(_05333_));
 sky130_fd_sc_hd__mux2_1 _12189_ (.A0(_06431_),
    .A1(_05333_),
    .S(net286),
    .X(_05334_));
 sky130_fd_sc_hd__a21oi_1 _12190_ (.A1(_05480_),
    .A2(_05334_),
    .B1(net236),
    .Y(_05335_));
 sky130_fd_sc_hd__o21a_1 _12191_ (.A1(_05480_),
    .A2(_05334_),
    .B1(_05335_),
    .X(_05336_));
 sky130_fd_sc_hd__o21a_1 _12192_ (.A1(_05270_),
    .A2(_05271_),
    .B1(_05272_),
    .X(_05337_));
 sky130_fd_sc_hd__nor2_1 _12193_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .Y(_05338_));
 sky130_fd_sc_hd__nand2_1 _12194_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .Y(_05340_));
 sky130_fd_sc_hd__and2b_1 _12195_ (.A_N(_05338_),
    .B(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__o21ai_1 _12196_ (.A1(_05337_),
    .A2(_05341_),
    .B1(net249),
    .Y(_05342_));
 sky130_fd_sc_hd__a21o_1 _12197_ (.A1(_05337_),
    .A2(_05341_),
    .B1(_05342_),
    .X(_05343_));
 sky130_fd_sc_hd__o211a_1 _12198_ (.A1(net250),
    .A2(_03103_),
    .B1(_05343_),
    .C1(net210),
    .X(_05344_));
 sky130_fd_sc_hd__or2_1 _12199_ (.A(\div_shifter[57] ),
    .B(_05277_),
    .X(_05345_));
 sky130_fd_sc_hd__a21oi_1 _12200_ (.A1(net233),
    .A2(_05345_),
    .B1(\div_shifter[58] ),
    .Y(_05346_));
 sky130_fd_sc_hd__a31o_1 _12201_ (.A1(\div_shifter[58] ),
    .A2(net233),
    .A3(_05345_),
    .B1(net192),
    .X(_05347_));
 sky130_fd_sc_hd__nor2_1 _12202_ (.A(_05346_),
    .B(_05347_),
    .Y(_05348_));
 sky130_fd_sc_hd__or2_1 _12203_ (.A(\div_res[25] ),
    .B(_05281_),
    .X(_05349_));
 sky130_fd_sc_hd__a21oi_1 _12204_ (.A1(net166),
    .A2(_05349_),
    .B1(\div_res[26] ),
    .Y(_05351_));
 sky130_fd_sc_hd__a31o_1 _12205_ (.A1(\div_res[26] ),
    .A2(net166),
    .A3(_05349_),
    .B1(net195),
    .X(_05352_));
 sky130_fd_sc_hd__nor2_1 _12206_ (.A(_05351_),
    .B(_05352_),
    .Y(_05353_));
 sky130_fd_sc_hd__mux2_1 _12207_ (.A0(_02320_),
    .A1(_02326_),
    .S(_05447_),
    .X(_05354_));
 sky130_fd_sc_hd__a21o_1 _12208_ (.A1(net198),
    .A2(_05354_),
    .B1(_05469_),
    .X(_05355_));
 sky130_fd_sc_hd__o21ai_1 _12209_ (.A1(_05436_),
    .A2(net209),
    .B1(_05355_),
    .Y(_05356_));
 sky130_fd_sc_hd__a221o_1 _12210_ (.A1(_02313_),
    .A2(_03103_),
    .B1(_03113_),
    .B2(net179),
    .C1(_05356_),
    .X(_05357_));
 sky130_fd_sc_hd__or4_1 _12211_ (.A(_05344_),
    .B(_05348_),
    .C(_05353_),
    .D(_05357_),
    .X(_05358_));
 sky130_fd_sc_hd__a21o_1 _12212_ (.A1(_01803_),
    .A2(_01887_),
    .B1(net160),
    .X(_05359_));
 sky130_fd_sc_hd__o21ai_1 _12213_ (.A1(_01892_),
    .A2(_05359_),
    .B1(_02323_),
    .Y(_05360_));
 sky130_fd_sc_hd__a21o_1 _12214_ (.A1(_01892_),
    .A2(_05359_),
    .B1(_05360_),
    .X(_05362_));
 sky130_fd_sc_hd__or4b_1 _12215_ (.A(_05332_),
    .B(_05336_),
    .C(_05358_),
    .D_N(_05362_),
    .X(_05363_));
 sky130_fd_sc_hd__and3_1 _12216_ (.A(curr_PC[25]),
    .B(curr_PC[26]),
    .C(_05215_),
    .X(_05364_));
 sky130_fd_sc_hd__a31o_1 _12217_ (.A1(curr_PC[24]),
    .A2(curr_PC[25]),
    .A3(_05132_),
    .B1(curr_PC[26]),
    .X(_05365_));
 sky130_fd_sc_hd__nand2_1 _12218_ (.A(_06457_),
    .B(_05365_),
    .Y(_05366_));
 sky130_fd_sc_hd__a2bb2o_4 _12219_ (.A1_N(_05364_),
    .A2_N(_05366_),
    .B1(net246),
    .B2(_05363_),
    .X(dest_val[26]));
 sky130_fd_sc_hd__xor2_1 _12220_ (.A(curr_PC[27]),
    .B(_05364_),
    .X(_05367_));
 sky130_fd_sc_hd__o22a_1 _12221_ (.A1(_00699_),
    .A2(net11),
    .B1(net6),
    .B2(_00409_),
    .X(_05368_));
 sky130_fd_sc_hd__xnor2_1 _12222_ (.A(net18),
    .B(_05368_),
    .Y(_05369_));
 sky130_fd_sc_hd__or2_1 _12223_ (.A(net92),
    .B(_05369_),
    .X(_05370_));
 sky130_fd_sc_hd__nand2_1 _12224_ (.A(net92),
    .B(_05369_),
    .Y(_05372_));
 sky130_fd_sc_hd__and2_1 _12225_ (.A(_05370_),
    .B(_05372_),
    .X(_05373_));
 sky130_fd_sc_hd__o22a_1 _12226_ (.A1(net15),
    .A2(net12),
    .B1(_02067_),
    .B2(net23),
    .X(_05374_));
 sky130_fd_sc_hd__xnor2_1 _12227_ (.A(net69),
    .B(_05374_),
    .Y(_05375_));
 sky130_fd_sc_hd__inv_2 _12228_ (.A(_05375_),
    .Y(_05376_));
 sky130_fd_sc_hd__nand2_1 _12229_ (.A(_05373_),
    .B(_05376_),
    .Y(_05377_));
 sky130_fd_sc_hd__or2_1 _12230_ (.A(_05373_),
    .B(_05376_),
    .X(_05378_));
 sky130_fd_sc_hd__nand2_1 _12231_ (.A(_05377_),
    .B(_05378_),
    .Y(_05379_));
 sky130_fd_sc_hd__o21a_1 _12232_ (.A1(net67),
    .A2(_05311_),
    .B1(net55),
    .X(_05380_));
 sky130_fd_sc_hd__or4_1 _12233_ (.A(net67),
    .B(net55),
    .C(net18),
    .D(_05311_),
    .X(_05381_));
 sky130_fd_sc_hd__or3b_1 _12234_ (.A(net18),
    .B(_05380_),
    .C_N(_05381_),
    .X(_05383_));
 sky130_fd_sc_hd__xor2_1 _12235_ (.A(_05302_),
    .B(_05383_),
    .X(_05384_));
 sky130_fd_sc_hd__and3_1 _12236_ (.A(_05377_),
    .B(_05378_),
    .C(_05384_),
    .X(_05385_));
 sky130_fd_sc_hd__xnor2_1 _12237_ (.A(_05379_),
    .B(_05384_),
    .Y(_05386_));
 sky130_fd_sc_hd__o21a_1 _12238_ (.A1(_05305_),
    .A2(_05309_),
    .B1(_05386_),
    .X(_05387_));
 sky130_fd_sc_hd__nor3_1 _12239_ (.A(_05305_),
    .B(_05309_),
    .C(_05386_),
    .Y(_05388_));
 sky130_fd_sc_hd__nor2_1 _12240_ (.A(_05387_),
    .B(_05388_),
    .Y(_05389_));
 sky130_fd_sc_hd__o21ai_2 _12241_ (.A1(_05314_),
    .A2(_05318_),
    .B1(_05389_),
    .Y(_05390_));
 sky130_fd_sc_hd__inv_2 _12242_ (.A(_05390_),
    .Y(_05391_));
 sky130_fd_sc_hd__or3_1 _12243_ (.A(_05314_),
    .B(_05318_),
    .C(_05389_),
    .X(_05392_));
 sky130_fd_sc_hd__nand2_2 _12244_ (.A(_05390_),
    .B(_05392_),
    .Y(_05394_));
 sky130_fd_sc_hd__nor2_1 _12245_ (.A(_05250_),
    .B(_05322_),
    .Y(_05395_));
 sky130_fd_sc_hd__o21ba_1 _12246_ (.A1(_05248_),
    .A2(_05320_),
    .B1_N(_05321_),
    .X(_05396_));
 sky130_fd_sc_hd__a21o_1 _12247_ (.A1(_05255_),
    .A2(_05395_),
    .B1(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__a31oi_4 _12248_ (.A1(_05097_),
    .A2(_05251_),
    .A3(_05395_),
    .B1(_05397_),
    .Y(_05398_));
 sky130_fd_sc_hd__xnor2_2 _12249_ (.A(_05394_),
    .B(_05398_),
    .Y(_05399_));
 sky130_fd_sc_hd__a31o_1 _12250_ (.A1(_05183_),
    .A2(_05327_),
    .A3(_05329_),
    .B1(net160),
    .X(_05400_));
 sky130_fd_sc_hd__a21oi_1 _12251_ (.A1(_05399_),
    .A2(_05400_),
    .B1(_02242_),
    .Y(_05401_));
 sky130_fd_sc_hd__o21a_1 _12252_ (.A1(_05399_),
    .A2(_05400_),
    .B1(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__o211a_1 _12253_ (.A1(_05480_),
    .A2(_05333_),
    .B1(net286),
    .C1(_05458_),
    .X(_05403_));
 sky130_fd_sc_hd__a21o_1 _12254_ (.A1(instruction[7]),
    .A2(_06432_),
    .B1(_05403_),
    .X(_05405_));
 sky130_fd_sc_hd__a21oi_1 _12255_ (.A1(_05198_),
    .A2(_05405_),
    .B1(net236),
    .Y(_05406_));
 sky130_fd_sc_hd__o21a_1 _12256_ (.A1(_05198_),
    .A2(_05405_),
    .B1(_05406_),
    .X(_05407_));
 sky130_fd_sc_hd__o21ai_1 _12257_ (.A1(net159),
    .A2(_01893_),
    .B1(_01894_),
    .Y(_05408_));
 sky130_fd_sc_hd__or3_1 _12258_ (.A(net159),
    .B(_01893_),
    .C(_01894_),
    .X(_05409_));
 sky130_fd_sc_hd__o21a_1 _12259_ (.A1(_05337_),
    .A2(_05338_),
    .B1(_05340_),
    .X(_05410_));
 sky130_fd_sc_hd__nor2_1 _12260_ (.A(reg1_val[27]),
    .B(curr_PC[27]),
    .Y(_05411_));
 sky130_fd_sc_hd__nand2_1 _12261_ (.A(reg1_val[27]),
    .B(curr_PC[27]),
    .Y(_05412_));
 sky130_fd_sc_hd__and2b_1 _12262_ (.A_N(_05411_),
    .B(_05412_),
    .X(_05413_));
 sky130_fd_sc_hd__o21ai_1 _12263_ (.A1(_05410_),
    .A2(_05413_),
    .B1(net249),
    .Y(_05414_));
 sky130_fd_sc_hd__a21o_1 _12264_ (.A1(_05410_),
    .A2(_05413_),
    .B1(_05414_),
    .X(_05416_));
 sky130_fd_sc_hd__o211a_1 _12265_ (.A1(net250),
    .A2(_02968_),
    .B1(_05416_),
    .C1(net210),
    .X(_05417_));
 sky130_fd_sc_hd__or2_1 _12266_ (.A(\div_res[26] ),
    .B(_05349_),
    .X(_05418_));
 sky130_fd_sc_hd__a21oi_1 _12267_ (.A1(net166),
    .A2(_05418_),
    .B1(\div_res[27] ),
    .Y(_05419_));
 sky130_fd_sc_hd__a31o_1 _12268_ (.A1(\div_res[27] ),
    .A2(net166),
    .A3(_05418_),
    .B1(net194),
    .X(_05420_));
 sky130_fd_sc_hd__nor2_1 _12269_ (.A(_05419_),
    .B(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__or2_1 _12270_ (.A(\div_shifter[58] ),
    .B(_05345_),
    .X(_05422_));
 sky130_fd_sc_hd__a21oi_1 _12271_ (.A1(net234),
    .A2(_05422_),
    .B1(\div_shifter[59] ),
    .Y(_05423_));
 sky130_fd_sc_hd__a311o_1 _12272_ (.A1(\div_shifter[59] ),
    .A2(net233),
    .A3(_05422_),
    .B1(_05423_),
    .C1(net192),
    .X(_05424_));
 sky130_fd_sc_hd__a21oi_1 _12273_ (.A1(_05187_),
    .A2(_02319_),
    .B1(_02315_),
    .Y(_05425_));
 sky130_fd_sc_hd__o221a_1 _12274_ (.A1(_05165_),
    .A2(net209),
    .B1(net196),
    .B2(_05187_),
    .C1(net246),
    .X(_05427_));
 sky130_fd_sc_hd__o21ai_1 _12275_ (.A1(_05176_),
    .A2(_05425_),
    .B1(_05427_),
    .Y(_05428_));
 sky130_fd_sc_hd__a221o_1 _12276_ (.A1(_02313_),
    .A2(_02968_),
    .B1(_02974_),
    .B2(net179),
    .C1(_05428_),
    .X(_05429_));
 sky130_fd_sc_hd__or4b_2 _12277_ (.A(_05417_),
    .B(_05421_),
    .C(_05429_),
    .D_N(_05424_),
    .X(_05430_));
 sky130_fd_sc_hd__a31o_1 _12278_ (.A1(_02323_),
    .A2(_05408_),
    .A3(_05409_),
    .B1(_05430_),
    .X(_05431_));
 sky130_fd_sc_hd__o32a_4 _12279_ (.A1(_05402_),
    .A2(_05407_),
    .A3(_05431_),
    .B1(_05367_),
    .B2(net246),
    .X(dest_val[27]));
 sky130_fd_sc_hd__o31a_1 _12280_ (.A1(net18),
    .A2(_05302_),
    .A3(_05380_),
    .B1(_05381_),
    .X(_05432_));
 sky130_fd_sc_hd__o22a_1 _12281_ (.A1(net12),
    .A2(net10),
    .B1(net5),
    .B2(_00699_),
    .X(_05433_));
 sky130_fd_sc_hd__xnor2_1 _12282_ (.A(net18),
    .B(_05433_),
    .Y(_05434_));
 sky130_fd_sc_hd__a21oi_1 _12283_ (.A1(_05370_),
    .A2(_05377_),
    .B1(_05434_),
    .Y(_05435_));
 sky130_fd_sc_hd__and3_1 _12284_ (.A(_05370_),
    .B(_05377_),
    .C(_05434_),
    .X(_05437_));
 sky130_fd_sc_hd__nor2_1 _12285_ (.A(_05435_),
    .B(_05437_),
    .Y(_05438_));
 sky130_fd_sc_hd__nor2_1 _12286_ (.A(_00409_),
    .B(net18),
    .Y(_05439_));
 sky130_fd_sc_hd__xnor2_1 _12287_ (.A(_05438_),
    .B(_05439_),
    .Y(_05440_));
 sky130_fd_sc_hd__o21a_1 _12288_ (.A1(net15),
    .A2(net7),
    .B1(_00678_),
    .X(_05441_));
 sky130_fd_sc_hd__a31o_1 _12289_ (.A1(net70),
    .A2(_00686_),
    .A3(net9),
    .B1(_05441_),
    .X(_05442_));
 sky130_fd_sc_hd__nor2_1 _12290_ (.A(_05440_),
    .B(_05442_),
    .Y(_05443_));
 sky130_fd_sc_hd__and2_1 _12291_ (.A(_05440_),
    .B(_05442_),
    .X(_05444_));
 sky130_fd_sc_hd__nor3_1 _12292_ (.A(_05432_),
    .B(_05443_),
    .C(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__o21a_1 _12293_ (.A1(_05443_),
    .A2(_05444_),
    .B1(_05432_),
    .X(_05446_));
 sky130_fd_sc_hd__nor2_1 _12294_ (.A(_05445_),
    .B(_05446_),
    .Y(_05448_));
 sky130_fd_sc_hd__o21ai_2 _12295_ (.A1(_05385_),
    .A2(_05387_),
    .B1(_05448_),
    .Y(_05449_));
 sky130_fd_sc_hd__nor3_1 _12296_ (.A(_05385_),
    .B(_05387_),
    .C(_05448_),
    .Y(_05450_));
 sky130_fd_sc_hd__inv_2 _12297_ (.A(_05450_),
    .Y(_05451_));
 sky130_fd_sc_hd__nand2_2 _12298_ (.A(_05449_),
    .B(_05451_),
    .Y(_05452_));
 sky130_fd_sc_hd__or2_1 _12299_ (.A(_05322_),
    .B(_05394_),
    .X(_05453_));
 sky130_fd_sc_hd__or3_1 _12300_ (.A(_05173_),
    .B(_05250_),
    .C(_05453_),
    .X(_05454_));
 sky130_fd_sc_hd__o21ai_1 _12301_ (.A1(_05320_),
    .A2(_05391_),
    .B1(_05392_),
    .Y(_05455_));
 sky130_fd_sc_hd__nand2_1 _12302_ (.A(_05178_),
    .B(_05323_),
    .Y(_05456_));
 sky130_fd_sc_hd__a21o_1 _12303_ (.A1(_05324_),
    .A2(_05456_),
    .B1(_05453_),
    .X(_05457_));
 sky130_fd_sc_hd__o311a_1 _12304_ (.A1(_04821_),
    .A2(_05175_),
    .A3(_05454_),
    .B1(_05455_),
    .C1(_05457_),
    .X(_05459_));
 sky130_fd_sc_hd__xnor2_2 _12305_ (.A(_05452_),
    .B(_05459_),
    .Y(_05460_));
 sky130_fd_sc_hd__and3_1 _12306_ (.A(_05327_),
    .B(_05329_),
    .C(_05399_),
    .X(_05461_));
 sky130_fd_sc_hd__a21o_1 _12307_ (.A1(_05183_),
    .A2(_05461_),
    .B1(net160),
    .X(_05462_));
 sky130_fd_sc_hd__a21oi_1 _12308_ (.A1(_05460_),
    .A2(_05462_),
    .B1(_02242_),
    .Y(_05463_));
 sky130_fd_sc_hd__o21a_1 _12309_ (.A1(_05460_),
    .A2(_05462_),
    .B1(_05463_),
    .X(_05464_));
 sky130_fd_sc_hd__a21o_1 _12310_ (.A1(_05187_),
    .A2(_05458_),
    .B1(_05176_),
    .X(_05465_));
 sky130_fd_sc_hd__o31ai_2 _12311_ (.A1(_05198_),
    .A2(_05480_),
    .A3(_05333_),
    .B1(_05465_),
    .Y(_05466_));
 sky130_fd_sc_hd__mux2_1 _12312_ (.A0(_06433_),
    .A1(_05466_),
    .S(net286),
    .X(_05467_));
 sky130_fd_sc_hd__nand2_1 _12313_ (.A(_05056_),
    .B(_05467_),
    .Y(_05468_));
 sky130_fd_sc_hd__o211a_1 _12314_ (.A1(_05056_),
    .A2(_05467_),
    .B1(_05468_),
    .C1(_02317_),
    .X(_05470_));
 sky130_fd_sc_hd__o21ai_1 _12315_ (.A1(net159),
    .A2(_01895_),
    .B1(_01901_),
    .Y(_05471_));
 sky130_fd_sc_hd__o311a_1 _12316_ (.A1(net159),
    .A2(_01895_),
    .A3(_01901_),
    .B1(_02323_),
    .C1(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__o21ai_2 _12317_ (.A1(_05410_),
    .A2(_05411_),
    .B1(_05412_),
    .Y(_05473_));
 sky130_fd_sc_hd__xor2_1 _12318_ (.A(reg1_val[28]),
    .B(_05473_),
    .X(_05474_));
 sky130_fd_sc_hd__or2_1 _12319_ (.A(net250),
    .B(_02830_),
    .X(_05475_));
 sky130_fd_sc_hd__o211a_1 _12320_ (.A1(_06331_),
    .A2(_05474_),
    .B1(_05475_),
    .C1(_06475_),
    .X(_05476_));
 sky130_fd_sc_hd__or2_1 _12321_ (.A(\div_res[27] ),
    .B(_05418_),
    .X(_05477_));
 sky130_fd_sc_hd__a21oi_1 _12322_ (.A1(net167),
    .A2(_05477_),
    .B1(\div_res[28] ),
    .Y(_05478_));
 sky130_fd_sc_hd__a31o_1 _12323_ (.A1(\div_res[28] ),
    .A2(net166),
    .A3(_05477_),
    .B1(net194),
    .X(_05479_));
 sky130_fd_sc_hd__or2_1 _12324_ (.A(\div_shifter[59] ),
    .B(_05422_),
    .X(_05481_));
 sky130_fd_sc_hd__a21oi_1 _12325_ (.A1(net233),
    .A2(_05481_),
    .B1(\div_shifter[60] ),
    .Y(_05482_));
 sky130_fd_sc_hd__a311o_1 _12326_ (.A1(\div_shifter[60] ),
    .A2(net233),
    .A3(_05481_),
    .B1(_05482_),
    .C1(net192),
    .X(_05483_));
 sky130_fd_sc_hd__o21ai_1 _12327_ (.A1(_05035_),
    .A2(_02320_),
    .B1(net198),
    .Y(_05484_));
 sky130_fd_sc_hd__a221o_1 _12328_ (.A1(_05035_),
    .A2(_02325_),
    .B1(_05484_),
    .B2(_05045_),
    .C1(net241),
    .X(_05485_));
 sky130_fd_sc_hd__a221oi_2 _12329_ (.A1(net179),
    .A2(_02820_),
    .B1(_02830_),
    .B2(_02313_),
    .C1(_05485_),
    .Y(_05486_));
 sky130_fd_sc_hd__o211a_1 _12330_ (.A1(_05478_),
    .A2(_05479_),
    .B1(_05483_),
    .C1(_05486_),
    .X(_05487_));
 sky130_fd_sc_hd__or4b_1 _12331_ (.A(_05470_),
    .B(_05472_),
    .C(_05476_),
    .D_N(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__o221a_4 _12332_ (.A1(_05024_),
    .A2(_06488_),
    .B1(_05464_),
    .B2(_05488_),
    .C1(net246),
    .X(dest_val[28]));
 sky130_fd_sc_hd__o22a_1 _12333_ (.A1(net10),
    .A2(net7),
    .B1(net5),
    .B2(net12),
    .X(_05489_));
 sky130_fd_sc_hd__xnor2_1 _12334_ (.A(net18),
    .B(_05489_),
    .Y(_05491_));
 sky130_fd_sc_hd__nor2_1 _12335_ (.A(_00699_),
    .B(net18),
    .Y(_05492_));
 sky130_fd_sc_hd__xnor2_1 _12336_ (.A(net69),
    .B(_05492_),
    .Y(_05493_));
 sky130_fd_sc_hd__nor2_1 _12337_ (.A(_05491_),
    .B(_05493_),
    .Y(_05494_));
 sky130_fd_sc_hd__and2_1 _12338_ (.A(_05491_),
    .B(_05493_),
    .X(_05495_));
 sky130_fd_sc_hd__nor2_1 _12339_ (.A(_05494_),
    .B(_05495_),
    .Y(_05496_));
 sky130_fd_sc_hd__nand2_1 _12340_ (.A(_05442_),
    .B(_05496_),
    .Y(_05497_));
 sky130_fd_sc_hd__or2_1 _12341_ (.A(_05442_),
    .B(_05496_),
    .X(_05498_));
 sky130_fd_sc_hd__nand2_1 _12342_ (.A(_05497_),
    .B(_05498_),
    .Y(_05499_));
 sky130_fd_sc_hd__a31o_1 _12343_ (.A1(_00408_),
    .A2(net22),
    .A3(_05438_),
    .B1(_05435_),
    .X(_05500_));
 sky130_fd_sc_hd__nand2b_1 _12344_ (.A_N(_05499_),
    .B(_05500_),
    .Y(_05502_));
 sky130_fd_sc_hd__xnor2_1 _12345_ (.A(_05499_),
    .B(_05500_),
    .Y(_05503_));
 sky130_fd_sc_hd__nor3_1 _12346_ (.A(_05443_),
    .B(_05445_),
    .C(_05503_),
    .Y(_05504_));
 sky130_fd_sc_hd__o21a_1 _12347_ (.A1(_05443_),
    .A2(_05445_),
    .B1(_05503_),
    .X(_05505_));
 sky130_fd_sc_hd__or2_2 _12348_ (.A(_05504_),
    .B(_05505_),
    .X(_05506_));
 sky130_fd_sc_hd__nor2_1 _12349_ (.A(_05394_),
    .B(_05452_),
    .Y(_05507_));
 sky130_fd_sc_hd__nand2_1 _12350_ (.A(_05395_),
    .B(_05507_),
    .Y(_05508_));
 sky130_fd_sc_hd__a21o_1 _12351_ (.A1(_05390_),
    .A2(_05449_),
    .B1(_05450_),
    .X(_05509_));
 sky130_fd_sc_hd__o2bb2a_1 _12352_ (.A1_N(_05396_),
    .A2_N(_05507_),
    .B1(_05508_),
    .B2(_05256_),
    .X(_05510_));
 sky130_fd_sc_hd__o311a_1 _12353_ (.A1(_04917_),
    .A2(_05253_),
    .A3(_05508_),
    .B1(_05509_),
    .C1(_05510_),
    .X(_05511_));
 sky130_fd_sc_hd__xnor2_2 _12354_ (.A(_05506_),
    .B(_05511_),
    .Y(_05513_));
 sky130_fd_sc_hd__a31o_1 _12355_ (.A1(_05183_),
    .A2(_05460_),
    .A3(_05461_),
    .B1(net160),
    .X(_05514_));
 sky130_fd_sc_hd__o21ai_1 _12356_ (.A1(_05513_),
    .A2(_05514_),
    .B1(net200),
    .Y(_05515_));
 sky130_fd_sc_hd__a21oi_1 _12357_ (.A1(_05513_),
    .A2(_05514_),
    .B1(_05515_),
    .Y(_05516_));
 sky130_fd_sc_hd__a21o_1 _12358_ (.A1(_05045_),
    .A2(_05466_),
    .B1(_05035_),
    .X(_05517_));
 sky130_fd_sc_hd__nand2_1 _12359_ (.A(net295),
    .B(_06434_),
    .Y(_05518_));
 sky130_fd_sc_hd__o21a_1 _12360_ (.A1(net295),
    .A2(_05517_),
    .B1(_05518_),
    .X(_05519_));
 sky130_fd_sc_hd__o21ai_1 _12361_ (.A1(_04969_),
    .A2(_05519_),
    .B1(_02317_),
    .Y(_05520_));
 sky130_fd_sc_hd__a21oi_1 _12362_ (.A1(_04969_),
    .A2(_05519_),
    .B1(_05520_),
    .Y(_05521_));
 sky130_fd_sc_hd__a21bo_1 _12363_ (.A1(net163),
    .A2(_01902_),
    .B1_N(_01802_),
    .X(_05522_));
 sky130_fd_sc_hd__or3b_1 _12364_ (.A(net159),
    .B(_01802_),
    .C_N(_01902_),
    .X(_05524_));
 sky130_fd_sc_hd__and3_1 _12365_ (.A(_02323_),
    .B(_05522_),
    .C(_05524_),
    .X(_05525_));
 sky130_fd_sc_hd__and3_1 _12366_ (.A(reg1_val[28]),
    .B(reg1_val[29]),
    .C(_05473_),
    .X(_05526_));
 sky130_fd_sc_hd__a21oi_1 _12367_ (.A1(reg1_val[28]),
    .A2(_05473_),
    .B1(reg1_val[29]),
    .Y(_05527_));
 sky130_fd_sc_hd__o21a_1 _12368_ (.A1(_05526_),
    .A2(_05527_),
    .B1(net250),
    .X(_05528_));
 sky130_fd_sc_hd__a211o_1 _12369_ (.A1(_06331_),
    .A2(_02651_),
    .B1(_05528_),
    .C1(_06476_),
    .X(_05529_));
 sky130_fd_sc_hd__or2_1 _12370_ (.A(\div_res[28] ),
    .B(_05477_),
    .X(_05530_));
 sky130_fd_sc_hd__a21oi_1 _12371_ (.A1(net166),
    .A2(_05530_),
    .B1(\div_res[29] ),
    .Y(_05531_));
 sky130_fd_sc_hd__a31o_1 _12372_ (.A1(\div_res[29] ),
    .A2(net166),
    .A3(_05530_),
    .B1(net194),
    .X(_05532_));
 sky130_fd_sc_hd__nor2_1 _12373_ (.A(_05531_),
    .B(_05532_),
    .Y(_05533_));
 sky130_fd_sc_hd__or2_1 _12374_ (.A(\div_shifter[60] ),
    .B(_05481_),
    .X(_05535_));
 sky130_fd_sc_hd__a21oi_1 _12375_ (.A1(net233),
    .A2(_05535_),
    .B1(\div_shifter[61] ),
    .Y(_05536_));
 sky130_fd_sc_hd__a311o_1 _12376_ (.A1(\div_shifter[61] ),
    .A2(net233),
    .A3(_05535_),
    .B1(_05536_),
    .C1(net192),
    .X(_05537_));
 sky130_fd_sc_hd__o21ai_1 _12377_ (.A1(_04948_),
    .A2(net197),
    .B1(net198),
    .Y(_05538_));
 sky130_fd_sc_hd__a221o_1 _12378_ (.A1(_04948_),
    .A2(_02325_),
    .B1(_05538_),
    .B2(_04958_),
    .C1(net241),
    .X(_05539_));
 sky130_fd_sc_hd__a221o_1 _12379_ (.A1(_02313_),
    .A2(_02652_),
    .B1(_02666_),
    .B2(net179),
    .C1(_05539_),
    .X(_05540_));
 sky130_fd_sc_hd__or3b_1 _12380_ (.A(_05533_),
    .B(_05540_),
    .C_N(_05537_),
    .X(_05541_));
 sky130_fd_sc_hd__or4b_1 _12381_ (.A(_05521_),
    .B(_05525_),
    .C(_05541_),
    .D_N(_05529_),
    .X(_05542_));
 sky130_fd_sc_hd__o221a_4 _12382_ (.A1(_04937_),
    .A2(_06488_),
    .B1(_05516_),
    .B2(_05542_),
    .C1(net246),
    .X(dest_val[29]));
 sky130_fd_sc_hd__a21o_1 _12383_ (.A1(net69),
    .A2(_05492_),
    .B1(_05494_),
    .X(_05543_));
 sky130_fd_sc_hd__o21ai_1 _12384_ (.A1(_01965_),
    .A2(net7),
    .B1(net18),
    .Y(_05545_));
 sky130_fd_sc_hd__or2_1 _12385_ (.A(net7),
    .B(_02080_),
    .X(_05546_));
 sky130_fd_sc_hd__o21ai_1 _12386_ (.A1(_01951_),
    .A2(_05546_),
    .B1(_05545_),
    .Y(_05547_));
 sky130_fd_sc_hd__a31o_1 _12387_ (.A1(_01951_),
    .A2(net22),
    .A3(_05546_),
    .B1(_05547_),
    .X(_05548_));
 sky130_fd_sc_hd__nand2_1 _12388_ (.A(_05543_),
    .B(_05548_),
    .Y(_05549_));
 sky130_fd_sc_hd__or2_1 _12389_ (.A(_05543_),
    .B(_05548_),
    .X(_05550_));
 sky130_fd_sc_hd__nand2_1 _12390_ (.A(_05549_),
    .B(_05550_),
    .Y(_05551_));
 sky130_fd_sc_hd__and3_1 _12391_ (.A(_05497_),
    .B(_05502_),
    .C(_05551_),
    .X(_05552_));
 sky130_fd_sc_hd__inv_2 _12392_ (.A(_05552_),
    .Y(_05553_));
 sky130_fd_sc_hd__a21oi_1 _12393_ (.A1(_05497_),
    .A2(_05502_),
    .B1(_05551_),
    .Y(_05554_));
 sky130_fd_sc_hd__or2_1 _12394_ (.A(_05552_),
    .B(_05554_),
    .X(_05556_));
 sky130_fd_sc_hd__o21ba_1 _12395_ (.A1(_05449_),
    .A2(_05504_),
    .B1_N(_05505_),
    .X(_05557_));
 sky130_fd_sc_hd__o31a_1 _12396_ (.A1(_05452_),
    .A2(_05455_),
    .A3(_05506_),
    .B1(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__o41a_1 _12397_ (.A1(_05326_),
    .A2(_05452_),
    .A3(_05453_),
    .A4(_05506_),
    .B1(_05558_),
    .X(_05559_));
 sky130_fd_sc_hd__xnor2_2 _12398_ (.A(_05556_),
    .B(_05559_),
    .Y(_05560_));
 sky130_fd_sc_hd__and2_1 _12399_ (.A(_05460_),
    .B(_05513_),
    .X(_05561_));
 sky130_fd_sc_hd__a31o_1 _12400_ (.A1(_05183_),
    .A2(_05461_),
    .A3(_05561_),
    .B1(net160),
    .X(_05562_));
 sky130_fd_sc_hd__o21ai_1 _12401_ (.A1(_05560_),
    .A2(_05562_),
    .B1(_02241_),
    .Y(_05563_));
 sky130_fd_sc_hd__a21oi_1 _12402_ (.A1(_05560_),
    .A2(_05562_),
    .B1(_05563_),
    .Y(_05564_));
 sky130_fd_sc_hd__a21oi_1 _12403_ (.A1(_04958_),
    .A2(_05517_),
    .B1(_04948_),
    .Y(_05565_));
 sky130_fd_sc_hd__mux2_1 _12404_ (.A0(_06435_),
    .A1(_05565_),
    .S(net286),
    .X(_05567_));
 sky130_fd_sc_hd__a21oi_1 _12405_ (.A1(_05133_),
    .A2(_05567_),
    .B1(net236),
    .Y(_05568_));
 sky130_fd_sc_hd__or2_1 _12406_ (.A(_05133_),
    .B(_05565_),
    .X(_05569_));
 sky130_fd_sc_hd__o21a_1 _12407_ (.A1(_05133_),
    .A2(_05567_),
    .B1(_05568_),
    .X(_05570_));
 sky130_fd_sc_hd__a21o_1 _12408_ (.A1(_01895_),
    .A2(_01903_),
    .B1(net159),
    .X(_05571_));
 sky130_fd_sc_hd__a21oi_1 _12409_ (.A1(_02015_),
    .A2(_05571_),
    .B1(_02324_),
    .Y(_05572_));
 sky130_fd_sc_hd__o21a_1 _12410_ (.A1(_02015_),
    .A2(_05571_),
    .B1(_05572_),
    .X(_05573_));
 sky130_fd_sc_hd__xor2_1 _12411_ (.A(reg1_val[30]),
    .B(_05526_),
    .X(_05574_));
 sky130_fd_sc_hd__nand2_1 _12412_ (.A(_06331_),
    .B(_02529_),
    .Y(_05575_));
 sky130_fd_sc_hd__o211a_1 _12413_ (.A1(_06331_),
    .A2(_05574_),
    .B1(_05575_),
    .C1(net210),
    .X(_05576_));
 sky130_fd_sc_hd__or2_1 _12414_ (.A(\div_shifter[61] ),
    .B(_05535_),
    .X(_05578_));
 sky130_fd_sc_hd__a21oi_1 _12415_ (.A1(net233),
    .A2(_05578_),
    .B1(\div_shifter[62] ),
    .Y(_05579_));
 sky130_fd_sc_hd__a311o_1 _12416_ (.A1(\div_shifter[62] ),
    .A2(net233),
    .A3(_05578_),
    .B1(_05579_),
    .C1(net193),
    .X(_05580_));
 sky130_fd_sc_hd__or2_1 _12417_ (.A(\div_res[29] ),
    .B(_05530_),
    .X(_05581_));
 sky130_fd_sc_hd__a21oi_1 _12418_ (.A1(net166),
    .A2(_05581_),
    .B1(\div_res[30] ),
    .Y(_05582_));
 sky130_fd_sc_hd__a31o_1 _12419_ (.A1(\div_res[30] ),
    .A2(net166),
    .A3(_05581_),
    .B1(net194),
    .X(_05583_));
 sky130_fd_sc_hd__mux2_1 _12420_ (.A0(net197),
    .A1(net196),
    .S(_05111_),
    .X(_05584_));
 sky130_fd_sc_hd__a21oi_1 _12421_ (.A1(net198),
    .A2(_05584_),
    .B1(_05122_),
    .Y(_05585_));
 sky130_fd_sc_hd__nor2_1 _12422_ (.A(net241),
    .B(_05585_),
    .Y(_05586_));
 sky130_fd_sc_hd__o221a_1 _12423_ (.A1(net177),
    .A2(_02500_),
    .B1(_02529_),
    .B2(_02314_),
    .C1(_05586_),
    .X(_05587_));
 sky130_fd_sc_hd__o211a_1 _12424_ (.A1(_05582_),
    .A2(_05583_),
    .B1(_05587_),
    .C1(_05580_),
    .X(_05589_));
 sky130_fd_sc_hd__or4b_1 _12425_ (.A(_05570_),
    .B(_05573_),
    .C(_05576_),
    .D_N(_05589_),
    .X(_05590_));
 sky130_fd_sc_hd__o221a_4 _12426_ (.A1(_05100_),
    .A2(_06488_),
    .B1(_05564_),
    .B2(_05590_),
    .C1(net246),
    .X(dest_val[30]));
 sky130_fd_sc_hd__a41o_1 _12427_ (.A1(_05183_),
    .A2(_05461_),
    .A3(_05560_),
    .A4(_05561_),
    .B1(net160),
    .X(_05591_));
 sky130_fd_sc_hd__nand2_1 _12428_ (.A(net7),
    .B(_02078_),
    .Y(_05592_));
 sky130_fd_sc_hd__or2_1 _12429_ (.A(_05506_),
    .B(_05556_),
    .X(_05593_));
 sky130_fd_sc_hd__or3_1 _12430_ (.A(_05394_),
    .B(_05452_),
    .C(_05593_),
    .X(_05594_));
 sky130_fd_sc_hd__a21oi_1 _12431_ (.A1(_05505_),
    .A2(_05553_),
    .B1(_05554_),
    .Y(_05595_));
 sky130_fd_sc_hd__o221a_1 _12432_ (.A1(_05509_),
    .A2(_05593_),
    .B1(_05594_),
    .B2(_05398_),
    .C1(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__xnor2_1 _12433_ (.A(_05592_),
    .B(_05596_),
    .Y(_05597_));
 sky130_fd_sc_hd__mux2_1 _12434_ (.A0(_05549_),
    .A1(_05543_),
    .S(_05547_),
    .X(_05599_));
 sky130_fd_sc_hd__xnor2_1 _12435_ (.A(_05597_),
    .B(_05599_),
    .Y(_05600_));
 sky130_fd_sc_hd__o21ai_1 _12436_ (.A1(_05591_),
    .A2(_05600_),
    .B1(_02241_),
    .Y(_05601_));
 sky130_fd_sc_hd__a21oi_1 _12437_ (.A1(_05591_),
    .A2(_05600_),
    .B1(_05601_),
    .Y(_05602_));
 sky130_fd_sc_hd__nor2_1 _12438_ (.A(net294),
    .B(_05111_),
    .Y(_05603_));
 sky130_fd_sc_hd__a22o_1 _12439_ (.A1(net294),
    .A2(_06436_),
    .B1(_05569_),
    .B2(_05603_),
    .X(_05604_));
 sky130_fd_sc_hd__a21oi_1 _12440_ (.A1(_05404_),
    .A2(_05604_),
    .B1(_02318_),
    .Y(_05605_));
 sky130_fd_sc_hd__o21a_1 _12441_ (.A1(_05404_),
    .A2(_05604_),
    .B1(_05605_),
    .X(_05606_));
 sky130_fd_sc_hd__o21ai_1 _12442_ (.A1(net159),
    .A2(_02016_),
    .B1(_02131_),
    .Y(_05607_));
 sky130_fd_sc_hd__o31a_1 _12443_ (.A1(net159),
    .A2(_02016_),
    .A3(_02131_),
    .B1(_02323_),
    .X(_05608_));
 sky130_fd_sc_hd__nand3_1 _12444_ (.A(reg1_val[30]),
    .B(net250),
    .C(_05526_),
    .Y(_05610_));
 sky130_fd_sc_hd__nand2_1 _12445_ (.A(_02343_),
    .B(_05610_),
    .Y(_05611_));
 sky130_fd_sc_hd__o211a_1 _12446_ (.A1(_02343_),
    .A2(_05610_),
    .B1(_05611_),
    .C1(net210),
    .X(_05612_));
 sky130_fd_sc_hd__o21ai_1 _12447_ (.A1(\div_res[30] ),
    .A2(_05581_),
    .B1(net166),
    .Y(_05613_));
 sky130_fd_sc_hd__xnor2_1 _12448_ (.A(\div_res[31] ),
    .B(_05613_),
    .Y(_05614_));
 sky130_fd_sc_hd__o21a_1 _12449_ (.A1(\div_shifter[62] ),
    .A2(_05578_),
    .B1(net233),
    .X(_05615_));
 sky130_fd_sc_hd__o21ai_1 _12450_ (.A1(\div_shifter[63] ),
    .A2(_05615_),
    .B1(_02330_),
    .Y(_05616_));
 sky130_fd_sc_hd__a21oi_1 _12451_ (.A1(\div_shifter[63] ),
    .A2(_05615_),
    .B1(_05616_),
    .Y(_05617_));
 sky130_fd_sc_hd__o21a_1 _12452_ (.A1(reg1_val[31]),
    .A2(_05382_),
    .B1(_02315_),
    .X(_05618_));
 sky130_fd_sc_hd__a311o_1 _12453_ (.A1(reg1_val[31]),
    .A2(_05382_),
    .A3(_02325_),
    .B1(_05618_),
    .C1(net241),
    .X(_05619_));
 sky130_fd_sc_hd__a221o_1 _12454_ (.A1(_05393_),
    .A2(_02319_),
    .B1(_02344_),
    .B2(_02313_),
    .C1(_05619_),
    .X(_05621_));
 sky130_fd_sc_hd__a211o_1 _12455_ (.A1(_02244_),
    .A2(_02308_),
    .B1(_05617_),
    .C1(_05621_),
    .X(_05622_));
 sky130_fd_sc_hd__a21o_1 _12456_ (.A1(_02328_),
    .A2(_05614_),
    .B1(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__a211o_1 _12457_ (.A1(_05607_),
    .A2(_05608_),
    .B1(_05612_),
    .C1(_05623_),
    .X(_05624_));
 sky130_fd_sc_hd__o21a_1 _12458_ (.A1(_05382_),
    .A2(net209),
    .B1(net247),
    .X(_05625_));
 sky130_fd_sc_hd__o31a_4 _12459_ (.A1(_05602_),
    .A2(_05606_),
    .A3(_05624_),
    .B1(_05625_),
    .X(dest_val[31]));
 sky130_fd_sc_hd__mux2_1 _12460_ (.A0(net293),
    .A1(curr_PC[0]),
    .S(net244),
    .X(_05626_));
 sky130_fd_sc_hd__nand2_1 _12461_ (.A(_04828_),
    .B(_05626_),
    .Y(_05627_));
 sky130_fd_sc_hd__or2_1 _12462_ (.A(_04828_),
    .B(_05626_),
    .X(_05628_));
 sky130_fd_sc_hd__and2_4 _12463_ (.A(_05627_),
    .B(_05628_),
    .X(new_PC[0]));
 sky130_fd_sc_hd__mux2_1 _12464_ (.A0(net289),
    .A1(curr_PC[1]),
    .S(net243),
    .X(_05630_));
 sky130_fd_sc_hd__nand2_1 _12465_ (.A(_05962_),
    .B(_05630_),
    .Y(_05631_));
 sky130_fd_sc_hd__or2_1 _12466_ (.A(_05962_),
    .B(_05630_),
    .X(_05632_));
 sky130_fd_sc_hd__nand2_1 _12467_ (.A(_05631_),
    .B(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__or2_1 _12468_ (.A(_05627_),
    .B(_05633_),
    .X(_05634_));
 sky130_fd_sc_hd__nand2_1 _12469_ (.A(_05627_),
    .B(_05633_),
    .Y(_05635_));
 sky130_fd_sc_hd__and2_4 _12470_ (.A(_05634_),
    .B(_05635_),
    .X(new_PC[1]));
 sky130_fd_sc_hd__mux2_1 _12471_ (.A0(reg1_val[2]),
    .A1(curr_PC[2]),
    .S(net243),
    .X(_05636_));
 sky130_fd_sc_hd__nand2_1 _12472_ (.A(_05916_),
    .B(_05636_),
    .Y(_05637_));
 sky130_fd_sc_hd__or2_1 _12473_ (.A(_05916_),
    .B(_05636_),
    .X(_05638_));
 sky130_fd_sc_hd__nand2_1 _12474_ (.A(_05637_),
    .B(_05638_),
    .Y(_05640_));
 sky130_fd_sc_hd__a21o_1 _12475_ (.A1(_05631_),
    .A2(_05634_),
    .B1(_05640_),
    .X(_05641_));
 sky130_fd_sc_hd__nand3_1 _12476_ (.A(_05631_),
    .B(_05634_),
    .C(_05640_),
    .Y(_05642_));
 sky130_fd_sc_hd__and2_4 _12477_ (.A(_05641_),
    .B(_05642_),
    .X(new_PC[2]));
 sky130_fd_sc_hd__mux2_1 _12478_ (.A0(reg1_val[3]),
    .A1(curr_PC[3]),
    .S(net244),
    .X(_05643_));
 sky130_fd_sc_hd__nand2_1 _12479_ (.A(_05854_),
    .B(_05643_),
    .Y(_05644_));
 sky130_fd_sc_hd__or2_1 _12480_ (.A(_05854_),
    .B(_05643_),
    .X(_05645_));
 sky130_fd_sc_hd__nand2_1 _12481_ (.A(_05644_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__a21o_1 _12482_ (.A1(_05637_),
    .A2(_05641_),
    .B1(_05646_),
    .X(_05647_));
 sky130_fd_sc_hd__nand3_1 _12483_ (.A(_05637_),
    .B(_05641_),
    .C(_05646_),
    .Y(_05648_));
 sky130_fd_sc_hd__and2_4 _12484_ (.A(_05647_),
    .B(_05648_),
    .X(new_PC[3]));
 sky130_fd_sc_hd__mux2_1 _12485_ (.A0(reg1_val[4]),
    .A1(curr_PC[4]),
    .S(net244),
    .X(_05650_));
 sky130_fd_sc_hd__nand2_1 _12486_ (.A(_05791_),
    .B(_05650_),
    .Y(_05651_));
 sky130_fd_sc_hd__or2_1 _12487_ (.A(_05791_),
    .B(_05650_),
    .X(_05652_));
 sky130_fd_sc_hd__nand2_1 _12488_ (.A(_05651_),
    .B(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__a21o_1 _12489_ (.A1(_05644_),
    .A2(_05647_),
    .B1(_05653_),
    .X(_05654_));
 sky130_fd_sc_hd__nand3_1 _12490_ (.A(_05644_),
    .B(_05647_),
    .C(_05653_),
    .Y(_05655_));
 sky130_fd_sc_hd__and2_4 _12491_ (.A(_05654_),
    .B(_05655_),
    .X(new_PC[4]));
 sky130_fd_sc_hd__mux2_1 _12492_ (.A0(reg1_val[5]),
    .A1(curr_PC[5]),
    .S(net244),
    .X(_05656_));
 sky130_fd_sc_hd__nand2_1 _12493_ (.A(_05649_),
    .B(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__or2_1 _12494_ (.A(_05649_),
    .B(_05656_),
    .X(_05659_));
 sky130_fd_sc_hd__nand2_1 _12495_ (.A(_05657_),
    .B(_05659_),
    .Y(_05660_));
 sky130_fd_sc_hd__a21o_1 _12496_ (.A1(_05651_),
    .A2(_05654_),
    .B1(_05660_),
    .X(_05661_));
 sky130_fd_sc_hd__nand3_1 _12497_ (.A(_05651_),
    .B(_05654_),
    .C(_05660_),
    .Y(_05662_));
 sky130_fd_sc_hd__and2_4 _12498_ (.A(_05661_),
    .B(_05662_),
    .X(new_PC[5]));
 sky130_fd_sc_hd__mux2_1 _12499_ (.A0(reg1_val[6]),
    .A1(curr_PC[6]),
    .S(net244),
    .X(_05663_));
 sky130_fd_sc_hd__nand2_1 _12500_ (.A(_05706_),
    .B(_05663_),
    .Y(_05664_));
 sky130_fd_sc_hd__or2_1 _12501_ (.A(_05706_),
    .B(_05663_),
    .X(_05665_));
 sky130_fd_sc_hd__nand2_1 _12502_ (.A(_05664_),
    .B(_05665_),
    .Y(_05666_));
 sky130_fd_sc_hd__a21o_1 _12503_ (.A1(_05657_),
    .A2(_05661_),
    .B1(_05666_),
    .X(_05667_));
 sky130_fd_sc_hd__nand3_1 _12504_ (.A(_05657_),
    .B(_05661_),
    .C(_05666_),
    .Y(_05669_));
 sky130_fd_sc_hd__and2_4 _12505_ (.A(_05667_),
    .B(_05669_),
    .X(new_PC[6]));
 sky130_fd_sc_hd__mux2_1 _12506_ (.A0(reg1_val[7]),
    .A1(curr_PC[7]),
    .S(net244),
    .X(_05670_));
 sky130_fd_sc_hd__nand2_1 _12507_ (.A(_05588_),
    .B(_05670_),
    .Y(_05671_));
 sky130_fd_sc_hd__or2_1 _12508_ (.A(_05588_),
    .B(_05670_),
    .X(_05672_));
 sky130_fd_sc_hd__nand2_1 _12509_ (.A(_05671_),
    .B(_05672_),
    .Y(_05673_));
 sky130_fd_sc_hd__a21o_1 _12510_ (.A1(_05664_),
    .A2(_05667_),
    .B1(_05673_),
    .X(_05674_));
 sky130_fd_sc_hd__nand3_1 _12511_ (.A(_05664_),
    .B(_05667_),
    .C(_05673_),
    .Y(_05675_));
 sky130_fd_sc_hd__and2_4 _12512_ (.A(_05674_),
    .B(_05675_),
    .X(new_PC[7]));
 sky130_fd_sc_hd__mux2_1 _12513_ (.A0(reg1_val[8]),
    .A1(curr_PC[8]),
    .S(net244),
    .X(_05676_));
 sky130_fd_sc_hd__nand2_1 _12514_ (.A(_05523_),
    .B(_05676_),
    .Y(_05678_));
 sky130_fd_sc_hd__or2_1 _12515_ (.A(_05523_),
    .B(_05676_),
    .X(_05679_));
 sky130_fd_sc_hd__nand2_1 _12516_ (.A(_05678_),
    .B(_05679_),
    .Y(_05680_));
 sky130_fd_sc_hd__a21o_1 _12517_ (.A1(_05671_),
    .A2(_05674_),
    .B1(_05680_),
    .X(_05681_));
 sky130_fd_sc_hd__nand3_1 _12518_ (.A(_05671_),
    .B(_05674_),
    .C(_05680_),
    .Y(_05682_));
 sky130_fd_sc_hd__and2_4 _12519_ (.A(_05681_),
    .B(_05682_),
    .X(new_PC[8]));
 sky130_fd_sc_hd__mux2_1 _12520_ (.A0(reg1_val[9]),
    .A1(curr_PC[9]),
    .S(net244),
    .X(_05683_));
 sky130_fd_sc_hd__nand2_1 _12521_ (.A(_05285_),
    .B(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__or2_1 _12522_ (.A(_05285_),
    .B(_05683_),
    .X(_05685_));
 sky130_fd_sc_hd__nand2_1 _12523_ (.A(_05684_),
    .B(_05685_),
    .Y(_05686_));
 sky130_fd_sc_hd__a21o_1 _12524_ (.A1(_05678_),
    .A2(_05681_),
    .B1(_05686_),
    .X(_05688_));
 sky130_fd_sc_hd__nand3_1 _12525_ (.A(_05678_),
    .B(_05681_),
    .C(_05686_),
    .Y(_05689_));
 sky130_fd_sc_hd__and2_4 _12526_ (.A(_05688_),
    .B(_05689_),
    .X(new_PC[9]));
 sky130_fd_sc_hd__mux2_1 _12527_ (.A0(reg1_val[10]),
    .A1(curr_PC[10]),
    .S(net245),
    .X(_05690_));
 sky130_fd_sc_hd__nand2_1 _12528_ (.A(_05219_),
    .B(_05690_),
    .Y(_05691_));
 sky130_fd_sc_hd__or2_1 _12529_ (.A(_05219_),
    .B(_05690_),
    .X(_05692_));
 sky130_fd_sc_hd__nand2_1 _12530_ (.A(_05691_),
    .B(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__a21o_1 _12531_ (.A1(_05684_),
    .A2(_05688_),
    .B1(_05693_),
    .X(_05694_));
 sky130_fd_sc_hd__nand3_1 _12532_ (.A(_05684_),
    .B(_05688_),
    .C(_05693_),
    .Y(_05695_));
 sky130_fd_sc_hd__and2_4 _12533_ (.A(_05694_),
    .B(_05695_),
    .X(new_PC[10]));
 sky130_fd_sc_hd__mux2_1 _12534_ (.A0(reg1_val[11]),
    .A1(curr_PC[11]),
    .S(net245),
    .X(_05697_));
 sky130_fd_sc_hd__nand2_1 _12535_ (.A(_05415_),
    .B(_05697_),
    .Y(_05698_));
 sky130_fd_sc_hd__or2_1 _12536_ (.A(_05415_),
    .B(_05697_),
    .X(_05699_));
 sky130_fd_sc_hd__nand2_1 _12537_ (.A(_05698_),
    .B(_05699_),
    .Y(_05700_));
 sky130_fd_sc_hd__a21o_1 _12538_ (.A1(_05691_),
    .A2(_05694_),
    .B1(_05700_),
    .X(_05701_));
 sky130_fd_sc_hd__nand3_1 _12539_ (.A(_05691_),
    .B(_05694_),
    .C(_05700_),
    .Y(_05702_));
 sky130_fd_sc_hd__and2_4 _12540_ (.A(_05701_),
    .B(_05702_),
    .X(new_PC[11]));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(reg1_val[12]),
    .A1(curr_PC[12]),
    .S(net245),
    .X(_05703_));
 sky130_fd_sc_hd__nand2_1 _12542_ (.A(_05143_),
    .B(_05703_),
    .Y(_05704_));
 sky130_fd_sc_hd__or2_1 _12543_ (.A(_05143_),
    .B(_05703_),
    .X(_05705_));
 sky130_fd_sc_hd__nand2_1 _12544_ (.A(_05704_),
    .B(_05705_),
    .Y(_05707_));
 sky130_fd_sc_hd__a21o_1 _12545_ (.A1(_05698_),
    .A2(_05701_),
    .B1(_05707_),
    .X(_05708_));
 sky130_fd_sc_hd__nand3_1 _12546_ (.A(_05698_),
    .B(_05701_),
    .C(_05707_),
    .Y(_05709_));
 sky130_fd_sc_hd__and2_4 _12547_ (.A(_05708_),
    .B(_05709_),
    .X(new_PC[12]));
 sky130_fd_sc_hd__mux2_1 _12548_ (.A0(reg1_val[13]),
    .A1(curr_PC[13]),
    .S(net245),
    .X(_05710_));
 sky130_fd_sc_hd__nand2_1 _12549_ (.A(_04991_),
    .B(_05710_),
    .Y(_05711_));
 sky130_fd_sc_hd__or2_1 _12550_ (.A(_04991_),
    .B(_05710_),
    .X(_05712_));
 sky130_fd_sc_hd__nand2_1 _12551_ (.A(_05711_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__a21o_1 _12552_ (.A1(_05704_),
    .A2(_05708_),
    .B1(_05713_),
    .X(_05714_));
 sky130_fd_sc_hd__nand3_1 _12553_ (.A(_05704_),
    .B(_05708_),
    .C(_05713_),
    .Y(_05715_));
 sky130_fd_sc_hd__and2_4 _12554_ (.A(_05714_),
    .B(_05715_),
    .X(new_PC[13]));
 sky130_fd_sc_hd__mux2_1 _12555_ (.A0(net291),
    .A1(curr_PC[14]),
    .S(net245),
    .X(_05717_));
 sky130_fd_sc_hd__nand2_1 _12556_ (.A(_04904_),
    .B(_05717_),
    .Y(_05718_));
 sky130_fd_sc_hd__or2_1 _12557_ (.A(_04904_),
    .B(_05717_),
    .X(_05719_));
 sky130_fd_sc_hd__nand2_1 _12558_ (.A(_05718_),
    .B(_05719_),
    .Y(_05720_));
 sky130_fd_sc_hd__a21o_1 _12559_ (.A1(_05711_),
    .A2(_05714_),
    .B1(_05720_),
    .X(_05721_));
 sky130_fd_sc_hd__nand3_1 _12560_ (.A(_05711_),
    .B(_05714_),
    .C(_05720_),
    .Y(_05722_));
 sky130_fd_sc_hd__and2_4 _12561_ (.A(_05721_),
    .B(_05722_),
    .X(new_PC[14]));
 sky130_fd_sc_hd__mux2_1 _12562_ (.A0(net290),
    .A1(curr_PC[15]),
    .S(net245),
    .X(_05723_));
 sky130_fd_sc_hd__nand2_1 _12563_ (.A(_05067_),
    .B(_05723_),
    .Y(_05724_));
 sky130_fd_sc_hd__or2_1 _12564_ (.A(_05067_),
    .B(_05723_),
    .X(_05726_));
 sky130_fd_sc_hd__nand2_1 _12565_ (.A(_05724_),
    .B(_05726_),
    .Y(_05727_));
 sky130_fd_sc_hd__a21o_1 _12566_ (.A1(_05718_),
    .A2(_05721_),
    .B1(_05727_),
    .X(_05728_));
 sky130_fd_sc_hd__nand3_1 _12567_ (.A(_05718_),
    .B(_05721_),
    .C(_05727_),
    .Y(_05729_));
 sky130_fd_sc_hd__and2_4 _12568_ (.A(_05728_),
    .B(_05729_),
    .X(new_PC[15]));
 sky130_fd_sc_hd__mux2_1 _12569_ (.A0(reg1_val[16]),
    .A1(curr_PC[16]),
    .S(net245),
    .X(_05730_));
 sky130_fd_sc_hd__xnor2_1 _12570_ (.A(net264),
    .B(_05730_),
    .Y(_05731_));
 sky130_fd_sc_hd__a21o_1 _12571_ (.A1(_05724_),
    .A2(_05728_),
    .B1(_05731_),
    .X(_05732_));
 sky130_fd_sc_hd__nand3_1 _12572_ (.A(_05724_),
    .B(_05728_),
    .C(_05731_),
    .Y(_05733_));
 sky130_fd_sc_hd__and2_4 _12573_ (.A(_05732_),
    .B(_05733_),
    .X(new_PC[16]));
 sky130_fd_sc_hd__mux2_2 _12574_ (.A0(reg1_val[17]),
    .A1(curr_PC[17]),
    .S(net245),
    .X(_05735_));
 sky130_fd_sc_hd__xnor2_4 _12575_ (.A(net264),
    .B(_05735_),
    .Y(_05736_));
 sky130_fd_sc_hd__a21bo_1 _12576_ (.A1(net264),
    .A2(_05730_),
    .B1_N(_05732_),
    .X(_05737_));
 sky130_fd_sc_hd__xnor2_4 _12577_ (.A(_05736_),
    .B(_05737_),
    .Y(new_PC[17]));
 sky130_fd_sc_hd__mux2_1 _12578_ (.A0(reg1_val[18]),
    .A1(curr_PC[18]),
    .S(net245),
    .X(_05738_));
 sky130_fd_sc_hd__nand2_1 _12579_ (.A(net263),
    .B(_05738_),
    .Y(_05739_));
 sky130_fd_sc_hd__or2_1 _12580_ (.A(net263),
    .B(_05738_),
    .X(_05740_));
 sky130_fd_sc_hd__nand2_1 _12581_ (.A(_05739_),
    .B(_05740_),
    .Y(_05741_));
 sky130_fd_sc_hd__or2_1 _12582_ (.A(_05732_),
    .B(_05736_),
    .X(_05742_));
 sky130_fd_sc_hd__o21ai_1 _12583_ (.A1(_05730_),
    .A2(_05735_),
    .B1(net264),
    .Y(_05743_));
 sky130_fd_sc_hd__a21o_1 _12584_ (.A1(_05742_),
    .A2(_05743_),
    .B1(_05741_),
    .X(_05745_));
 sky130_fd_sc_hd__nand3_1 _12585_ (.A(_05741_),
    .B(_05742_),
    .C(_05743_),
    .Y(_05746_));
 sky130_fd_sc_hd__and2_4 _12586_ (.A(_05745_),
    .B(_05746_),
    .X(new_PC[18]));
 sky130_fd_sc_hd__mux2_1 _12587_ (.A0(reg1_val[19]),
    .A1(curr_PC[19]),
    .S(net245),
    .X(_05747_));
 sky130_fd_sc_hd__nand2_1 _12588_ (.A(net263),
    .B(_05747_),
    .Y(_05748_));
 sky130_fd_sc_hd__or2_1 _12589_ (.A(net263),
    .B(_05747_),
    .X(_05749_));
 sky130_fd_sc_hd__nand2_2 _12590_ (.A(_05748_),
    .B(_05749_),
    .Y(_05750_));
 sky130_fd_sc_hd__nand2_2 _12591_ (.A(_05739_),
    .B(_05745_),
    .Y(_05751_));
 sky130_fd_sc_hd__xnor2_4 _12592_ (.A(_05750_),
    .B(_05751_),
    .Y(new_PC[19]));
 sky130_fd_sc_hd__mux2_1 _12593_ (.A0(reg1_val[20]),
    .A1(curr_PC[20]),
    .S(net245),
    .X(_05752_));
 sky130_fd_sc_hd__nand2_1 _12594_ (.A(net263),
    .B(_05752_),
    .Y(_05754_));
 sky130_fd_sc_hd__or2_1 _12595_ (.A(net263),
    .B(_05752_),
    .X(_05755_));
 sky130_fd_sc_hd__nand2_2 _12596_ (.A(_05754_),
    .B(_05755_),
    .Y(_05756_));
 sky130_fd_sc_hd__or3_1 _12597_ (.A(_05741_),
    .B(_05742_),
    .C(_05750_),
    .X(_05757_));
 sky130_fd_sc_hd__and3_1 _12598_ (.A(_05739_),
    .B(_05743_),
    .C(_05748_),
    .X(_05758_));
 sky130_fd_sc_hd__nand2_2 _12599_ (.A(_05757_),
    .B(_05758_),
    .Y(_05759_));
 sky130_fd_sc_hd__inv_2 _12600_ (.A(_05759_),
    .Y(_05760_));
 sky130_fd_sc_hd__xnor2_4 _12601_ (.A(_05756_),
    .B(_05759_),
    .Y(new_PC[20]));
 sky130_fd_sc_hd__mux2_2 _12602_ (.A0(reg1_val[21]),
    .A1(curr_PC[21]),
    .S(net246),
    .X(_05761_));
 sky130_fd_sc_hd__xnor2_4 _12603_ (.A(net263),
    .B(_05761_),
    .Y(_05762_));
 sky130_fd_sc_hd__o21ai_2 _12604_ (.A1(_05756_),
    .A2(_05760_),
    .B1(_05754_),
    .Y(_05764_));
 sky130_fd_sc_hd__xnor2_4 _12605_ (.A(_05762_),
    .B(_05764_),
    .Y(new_PC[21]));
 sky130_fd_sc_hd__mux2_1 _12606_ (.A0(reg1_val[22]),
    .A1(curr_PC[22]),
    .S(net246),
    .X(_05765_));
 sky130_fd_sc_hd__and2_1 _12607_ (.A(net263),
    .B(_05765_),
    .X(_05766_));
 sky130_fd_sc_hd__or2_1 _12608_ (.A(net263),
    .B(_05765_),
    .X(_05767_));
 sky130_fd_sc_hd__nand2b_2 _12609_ (.A_N(_05766_),
    .B(_05767_),
    .Y(_05768_));
 sky130_fd_sc_hd__o21ai_2 _12610_ (.A1(_05752_),
    .A2(_05761_),
    .B1(net263),
    .Y(_05769_));
 sky130_fd_sc_hd__nor2_1 _12611_ (.A(_05756_),
    .B(_05762_),
    .Y(_05770_));
 sky130_fd_sc_hd__inv_2 _12612_ (.A(_05770_),
    .Y(_05771_));
 sky130_fd_sc_hd__o21ai_4 _12613_ (.A1(_05760_),
    .A2(_05771_),
    .B1(_05769_),
    .Y(_05772_));
 sky130_fd_sc_hd__xnor2_4 _12614_ (.A(_05768_),
    .B(_05772_),
    .Y(new_PC[22]));
 sky130_fd_sc_hd__mux2_2 _12615_ (.A0(reg1_val[23]),
    .A1(curr_PC[23]),
    .S(net245),
    .X(_05774_));
 sky130_fd_sc_hd__xnor2_4 _12616_ (.A(net263),
    .B(_05774_),
    .Y(_05775_));
 sky130_fd_sc_hd__a21o_1 _12617_ (.A1(_05767_),
    .A2(_05772_),
    .B1(_05766_),
    .X(_05776_));
 sky130_fd_sc_hd__xnor2_4 _12618_ (.A(_05775_),
    .B(_05776_),
    .Y(new_PC[23]));
 sky130_fd_sc_hd__mux2_2 _12619_ (.A0(reg1_val[24]),
    .A1(curr_PC[24]),
    .S(net245),
    .X(_05777_));
 sky130_fd_sc_hd__xnor2_4 _12620_ (.A(net264),
    .B(_05777_),
    .Y(_05778_));
 sky130_fd_sc_hd__or4_1 _12621_ (.A(_05757_),
    .B(_05768_),
    .C(_05771_),
    .D(_05775_),
    .X(_05779_));
 sky130_fd_sc_hd__o21ai_1 _12622_ (.A1(_05765_),
    .A2(_05774_),
    .B1(net263),
    .Y(_05780_));
 sky130_fd_sc_hd__and4_2 _12623_ (.A(_05758_),
    .B(_05769_),
    .C(_05779_),
    .D(_05780_),
    .X(_05781_));
 sky130_fd_sc_hd__xor2_4 _12624_ (.A(_05778_),
    .B(_05781_),
    .X(new_PC[24]));
 sky130_fd_sc_hd__mux2_1 _12625_ (.A0(reg1_val[25]),
    .A1(curr_PC[25]),
    .S(net245),
    .X(_05783_));
 sky130_fd_sc_hd__and2_1 _12626_ (.A(net264),
    .B(_05783_),
    .X(_05784_));
 sky130_fd_sc_hd__nor2_1 _12627_ (.A(net263),
    .B(_05783_),
    .Y(_05785_));
 sky130_fd_sc_hd__nor2_2 _12628_ (.A(_05784_),
    .B(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__o2bb2a_2 _12629_ (.A1_N(net263),
    .A2_N(_05777_),
    .B1(_05778_),
    .B2(_05781_),
    .X(_05787_));
 sky130_fd_sc_hd__xnor2_4 _12630_ (.A(_05786_),
    .B(_05787_),
    .Y(new_PC[25]));
 sky130_fd_sc_hd__mux2_1 _12631_ (.A0(reg1_val[26]),
    .A1(curr_PC[26]),
    .S(net246),
    .X(_05788_));
 sky130_fd_sc_hd__and2_1 _12632_ (.A(net263),
    .B(_05788_),
    .X(_05789_));
 sky130_fd_sc_hd__nor2_1 _12633_ (.A(net263),
    .B(_05788_),
    .Y(_05790_));
 sky130_fd_sc_hd__nor2_2 _12634_ (.A(_05789_),
    .B(_05790_),
    .Y(_05792_));
 sky130_fd_sc_hd__o21ba_2 _12635_ (.A1(_05785_),
    .A2(_05787_),
    .B1_N(_05784_),
    .X(_05793_));
 sky130_fd_sc_hd__xnor2_4 _12636_ (.A(_05792_),
    .B(_05793_),
    .Y(new_PC[26]));
 sky130_fd_sc_hd__o21ba_1 _12637_ (.A1(_05790_),
    .A2(_05793_),
    .B1_N(_05789_),
    .X(_05794_));
 sky130_fd_sc_hd__mux2_2 _12638_ (.A0(reg1_val[27]),
    .A1(curr_PC[27]),
    .S(net245),
    .X(_05795_));
 sky130_fd_sc_hd__xor2_2 _12639_ (.A(net264),
    .B(_05795_),
    .X(_05796_));
 sky130_fd_sc_hd__xnor2_4 _12640_ (.A(_05794_),
    .B(_05796_),
    .Y(new_PC[27]));
 sky130_fd_sc_hd__nand2_2 _12641_ (.A(net292),
    .B(_04828_),
    .Y(_05797_));
 sky130_fd_sc_hd__or2_1 _12642_ (.A(net292),
    .B(_04828_),
    .X(_05798_));
 sky130_fd_sc_hd__and2_4 _12643_ (.A(_05797_),
    .B(_05798_),
    .X(loadstore_address[0]));
 sky130_fd_sc_hd__or2_1 _12644_ (.A(net289),
    .B(_05962_),
    .X(_05800_));
 sky130_fd_sc_hd__nand2_1 _12645_ (.A(reg1_val[1]),
    .B(_05962_),
    .Y(_05801_));
 sky130_fd_sc_hd__nand2_2 _12646_ (.A(_05800_),
    .B(_05801_),
    .Y(_05802_));
 sky130_fd_sc_hd__xor2_4 _12647_ (.A(_05797_),
    .B(_05802_),
    .X(loadstore_address[1]));
 sky130_fd_sc_hd__o21a_2 _12648_ (.A1(_05797_),
    .A2(_05802_),
    .B1(_05801_),
    .X(_05803_));
 sky130_fd_sc_hd__nor2_1 _12649_ (.A(reg1_val[2]),
    .B(_05916_),
    .Y(_05804_));
 sky130_fd_sc_hd__nand2_1 _12650_ (.A(reg1_val[2]),
    .B(_05916_),
    .Y(_05805_));
 sky130_fd_sc_hd__and2b_1 _12651_ (.A_N(_05804_),
    .B(_05805_),
    .X(_05806_));
 sky130_fd_sc_hd__xnor2_4 _12652_ (.A(_05803_),
    .B(_05806_),
    .Y(loadstore_address[2]));
 sky130_fd_sc_hd__o21a_2 _12653_ (.A1(_05803_),
    .A2(_05804_),
    .B1(_05805_),
    .X(_05807_));
 sky130_fd_sc_hd__nor2_1 _12654_ (.A(reg1_val[3]),
    .B(_05854_),
    .Y(_05809_));
 sky130_fd_sc_hd__nand2_1 _12655_ (.A(reg1_val[3]),
    .B(_05854_),
    .Y(_05810_));
 sky130_fd_sc_hd__and2b_1 _12656_ (.A_N(_05809_),
    .B(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__xnor2_4 _12657_ (.A(_05807_),
    .B(_05811_),
    .Y(loadstore_address[3]));
 sky130_fd_sc_hd__o21a_2 _12658_ (.A1(_05807_),
    .A2(_05809_),
    .B1(_05810_),
    .X(_05812_));
 sky130_fd_sc_hd__nor2_1 _12659_ (.A(reg1_val[4]),
    .B(_05791_),
    .Y(_05813_));
 sky130_fd_sc_hd__nand2_1 _12660_ (.A(reg1_val[4]),
    .B(_05791_),
    .Y(_05814_));
 sky130_fd_sc_hd__and2b_1 _12661_ (.A_N(_05813_),
    .B(_05814_),
    .X(_05815_));
 sky130_fd_sc_hd__xnor2_4 _12662_ (.A(_05812_),
    .B(_05815_),
    .Y(loadstore_address[4]));
 sky130_fd_sc_hd__o21a_2 _12663_ (.A1(_05812_),
    .A2(_05813_),
    .B1(_05814_),
    .X(_05816_));
 sky130_fd_sc_hd__nor2_1 _12664_ (.A(reg1_val[5]),
    .B(_05649_),
    .Y(_05818_));
 sky130_fd_sc_hd__nand2_1 _12665_ (.A(reg1_val[5]),
    .B(_05649_),
    .Y(_05819_));
 sky130_fd_sc_hd__nand2b_2 _12666_ (.A_N(_05818_),
    .B(_05819_),
    .Y(_05820_));
 sky130_fd_sc_hd__xor2_4 _12667_ (.A(_05816_),
    .B(_05820_),
    .X(loadstore_address[5]));
 sky130_fd_sc_hd__o21a_2 _12668_ (.A1(_05816_),
    .A2(_05818_),
    .B1(_05819_),
    .X(_05821_));
 sky130_fd_sc_hd__nor2_1 _12669_ (.A(reg1_val[6]),
    .B(_05706_),
    .Y(_05822_));
 sky130_fd_sc_hd__and2_1 _12670_ (.A(reg1_val[6]),
    .B(_05706_),
    .X(_05823_));
 sky130_fd_sc_hd__or2_2 _12671_ (.A(_05822_),
    .B(_05823_),
    .X(_05824_));
 sky130_fd_sc_hd__xor2_4 _12672_ (.A(_05821_),
    .B(_05824_),
    .X(loadstore_address[6]));
 sky130_fd_sc_hd__o21ba_2 _12673_ (.A1(_05821_),
    .A2(_05822_),
    .B1_N(_05823_),
    .X(_05825_));
 sky130_fd_sc_hd__nor2_1 _12674_ (.A(reg1_val[7]),
    .B(_05588_),
    .Y(_05827_));
 sky130_fd_sc_hd__nand2_1 _12675_ (.A(reg1_val[7]),
    .B(_05588_),
    .Y(_05828_));
 sky130_fd_sc_hd__nand2b_2 _12676_ (.A_N(_05827_),
    .B(_05828_),
    .Y(_05829_));
 sky130_fd_sc_hd__xor2_4 _12677_ (.A(_05825_),
    .B(_05829_),
    .X(loadstore_address[7]));
 sky130_fd_sc_hd__o21a_2 _12678_ (.A1(_05825_),
    .A2(_05827_),
    .B1(_05828_),
    .X(_05830_));
 sky130_fd_sc_hd__nor2_1 _12679_ (.A(reg1_val[8]),
    .B(_05523_),
    .Y(_05831_));
 sky130_fd_sc_hd__nand2_1 _12680_ (.A(reg1_val[8]),
    .B(_05523_),
    .Y(_05832_));
 sky130_fd_sc_hd__nand2b_2 _12681_ (.A_N(_05831_),
    .B(_05832_),
    .Y(_05833_));
 sky130_fd_sc_hd__xor2_4 _12682_ (.A(_05830_),
    .B(_05833_),
    .X(loadstore_address[8]));
 sky130_fd_sc_hd__o21a_2 _12683_ (.A1(_05830_),
    .A2(_05831_),
    .B1(_05832_),
    .X(_05834_));
 sky130_fd_sc_hd__or2_1 _12684_ (.A(reg1_val[9]),
    .B(_05285_),
    .X(_05836_));
 sky130_fd_sc_hd__nand2_1 _12685_ (.A(reg1_val[9]),
    .B(_05285_),
    .Y(_05837_));
 sky130_fd_sc_hd__nand2_2 _12686_ (.A(_05836_),
    .B(_05837_),
    .Y(_05838_));
 sky130_fd_sc_hd__xor2_4 _12687_ (.A(_05834_),
    .B(_05838_),
    .X(loadstore_address[9]));
 sky130_fd_sc_hd__nand2_1 _12688_ (.A(reg1_val[10]),
    .B(_05219_),
    .Y(_05839_));
 sky130_fd_sc_hd__or2_1 _12689_ (.A(reg1_val[10]),
    .B(_05219_),
    .X(_05840_));
 sky130_fd_sc_hd__nand2_1 _12690_ (.A(_05839_),
    .B(_05840_),
    .Y(_05841_));
 sky130_fd_sc_hd__nand2b_1 _12691_ (.A_N(_05834_),
    .B(_05836_),
    .Y(_05842_));
 sky130_fd_sc_hd__a21o_1 _12692_ (.A1(_05837_),
    .A2(_05842_),
    .B1(_05841_),
    .X(_05843_));
 sky130_fd_sc_hd__nand3_1 _12693_ (.A(_05837_),
    .B(_05841_),
    .C(_05842_),
    .Y(_05844_));
 sky130_fd_sc_hd__and2_4 _12694_ (.A(_05843_),
    .B(_05844_),
    .X(loadstore_address[10]));
 sky130_fd_sc_hd__nand2_1 _12695_ (.A(reg1_val[11]),
    .B(_05415_),
    .Y(_05846_));
 sky130_fd_sc_hd__or2_1 _12696_ (.A(reg1_val[11]),
    .B(_05415_),
    .X(_05847_));
 sky130_fd_sc_hd__nand2_1 _12697_ (.A(_05846_),
    .B(_05847_),
    .Y(_05848_));
 sky130_fd_sc_hd__a21o_1 _12698_ (.A1(_05839_),
    .A2(_05843_),
    .B1(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__nand3_1 _12699_ (.A(_05839_),
    .B(_05843_),
    .C(_05848_),
    .Y(_05850_));
 sky130_fd_sc_hd__and2_4 _12700_ (.A(_05849_),
    .B(_05850_),
    .X(loadstore_address[11]));
 sky130_fd_sc_hd__nand2_1 _12701_ (.A(reg1_val[12]),
    .B(_05143_),
    .Y(_05851_));
 sky130_fd_sc_hd__or2_1 _12702_ (.A(reg1_val[12]),
    .B(_05143_),
    .X(_05852_));
 sky130_fd_sc_hd__nand2_1 _12703_ (.A(_05851_),
    .B(_05852_),
    .Y(_05853_));
 sky130_fd_sc_hd__a21o_1 _12704_ (.A1(_05846_),
    .A2(_05849_),
    .B1(_05853_),
    .X(_05855_));
 sky130_fd_sc_hd__nand3_1 _12705_ (.A(_05846_),
    .B(_05849_),
    .C(_05853_),
    .Y(_05856_));
 sky130_fd_sc_hd__and2_4 _12706_ (.A(_05855_),
    .B(_05856_),
    .X(loadstore_address[12]));
 sky130_fd_sc_hd__nand2_1 _12707_ (.A(reg1_val[13]),
    .B(_04991_),
    .Y(_05857_));
 sky130_fd_sc_hd__or2_1 _12708_ (.A(reg1_val[13]),
    .B(_04991_),
    .X(_05858_));
 sky130_fd_sc_hd__nand2_1 _12709_ (.A(_05857_),
    .B(_05858_),
    .Y(_05859_));
 sky130_fd_sc_hd__a21o_1 _12710_ (.A1(_05851_),
    .A2(_05855_),
    .B1(_05859_),
    .X(_05860_));
 sky130_fd_sc_hd__nand3_1 _12711_ (.A(_05851_),
    .B(_05855_),
    .C(_05859_),
    .Y(_05861_));
 sky130_fd_sc_hd__and2_4 _12712_ (.A(_05860_),
    .B(_05861_),
    .X(loadstore_address[13]));
 sky130_fd_sc_hd__nand2_2 _12713_ (.A(reg1_val[14]),
    .B(_04904_),
    .Y(_05862_));
 sky130_fd_sc_hd__or2_1 _12714_ (.A(reg1_val[14]),
    .B(_04904_),
    .X(_05864_));
 sky130_fd_sc_hd__nand2_1 _12715_ (.A(_05862_),
    .B(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__a21o_1 _12716_ (.A1(_05857_),
    .A2(_05860_),
    .B1(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__nand3_1 _12717_ (.A(_05857_),
    .B(_05860_),
    .C(_05865_),
    .Y(_05867_));
 sky130_fd_sc_hd__and2_4 _12718_ (.A(_05866_),
    .B(_05867_),
    .X(loadstore_address[14]));
 sky130_fd_sc_hd__xnor2_2 _12719_ (.A(reg1_val[15]),
    .B(_05067_),
    .Y(_05868_));
 sky130_fd_sc_hd__a21oi_4 _12720_ (.A1(_05862_),
    .A2(_05866_),
    .B1(_05868_),
    .Y(_05869_));
 sky130_fd_sc_hd__and3_2 _12721_ (.A(_05862_),
    .B(_05866_),
    .C(_05868_),
    .X(_05870_));
 sky130_fd_sc_hd__nor2_8 _12722_ (.A(_05869_),
    .B(_05870_),
    .Y(loadstore_address[15]));
 sky130_fd_sc_hd__xor2_4 _12723_ (.A(reg1_val[16]),
    .B(net265),
    .X(_05871_));
 sky130_fd_sc_hd__a21o_2 _12724_ (.A1(reg1_val[15]),
    .A2(_05067_),
    .B1(_05869_),
    .X(_05873_));
 sky130_fd_sc_hd__nand2_1 _12725_ (.A(_05871_),
    .B(_05873_),
    .Y(_05874_));
 sky130_fd_sc_hd__xor2_4 _12726_ (.A(_05871_),
    .B(_05873_),
    .X(loadstore_address[16]));
 sky130_fd_sc_hd__a21bo_1 _12727_ (.A1(reg1_val[16]),
    .A2(net265),
    .B1_N(_05874_),
    .X(_05875_));
 sky130_fd_sc_hd__xnor2_4 _12728_ (.A(reg1_val[17]),
    .B(net265),
    .Y(_05876_));
 sky130_fd_sc_hd__xnor2_4 _12729_ (.A(_05875_),
    .B(_05876_),
    .Y(loadstore_address[17]));
 sky130_fd_sc_hd__nand2_2 _12730_ (.A(reg1_val[18]),
    .B(net265),
    .Y(_05877_));
 sky130_fd_sc_hd__or2_1 _12731_ (.A(reg1_val[18]),
    .B(net265),
    .X(_05878_));
 sky130_fd_sc_hd__nand2_4 _12732_ (.A(_05877_),
    .B(_05878_),
    .Y(_05879_));
 sky130_fd_sc_hd__o2bb2a_2 _12733_ (.A1_N(net265),
    .A2_N(_00200_),
    .B1(_05874_),
    .B2(_05876_),
    .X(_05880_));
 sky130_fd_sc_hd__xor2_4 _12734_ (.A(_05879_),
    .B(_05880_),
    .X(loadstore_address[18]));
 sky130_fd_sc_hd__o21ai_4 _12735_ (.A1(_05879_),
    .A2(_05880_),
    .B1(_05877_),
    .Y(_05882_));
 sky130_fd_sc_hd__xnor2_4 _12736_ (.A(reg1_val[19]),
    .B(net265),
    .Y(_05883_));
 sky130_fd_sc_hd__xnor2_4 _12737_ (.A(_05882_),
    .B(_05883_),
    .Y(loadstore_address[19]));
 sky130_fd_sc_hd__xnor2_2 _12738_ (.A(reg1_val[20]),
    .B(net265),
    .Y(_05884_));
 sky130_fd_sc_hd__or4_2 _12739_ (.A(_05874_),
    .B(_05876_),
    .C(_05879_),
    .D(_05883_),
    .X(_05885_));
 sky130_fd_sc_hd__nand2_1 _12740_ (.A(net265),
    .B(_00201_),
    .Y(_05886_));
 sky130_fd_sc_hd__a21oi_4 _12741_ (.A1(_05885_),
    .A2(_05886_),
    .B1(_05884_),
    .Y(_05887_));
 sky130_fd_sc_hd__and3_2 _12742_ (.A(_05884_),
    .B(_05885_),
    .C(_05886_),
    .X(_05888_));
 sky130_fd_sc_hd__nor2_8 _12743_ (.A(_05887_),
    .B(_05888_),
    .Y(loadstore_address[20]));
 sky130_fd_sc_hd__nor2_1 _12744_ (.A(reg1_val[21]),
    .B(net265),
    .Y(_05890_));
 sky130_fd_sc_hd__nand2_1 _12745_ (.A(reg1_val[21]),
    .B(net265),
    .Y(_05891_));
 sky130_fd_sc_hd__nand2b_2 _12746_ (.A_N(_05890_),
    .B(_05891_),
    .Y(_05892_));
 sky130_fd_sc_hd__a21oi_4 _12747_ (.A1(reg1_val[20]),
    .A2(net265),
    .B1(_05887_),
    .Y(_05893_));
 sky130_fd_sc_hd__xor2_4 _12748_ (.A(_05892_),
    .B(_05893_),
    .X(loadstore_address[21]));
 sky130_fd_sc_hd__nand2_2 _12749_ (.A(reg1_val[22]),
    .B(net265),
    .Y(_05894_));
 sky130_fd_sc_hd__or2_1 _12750_ (.A(reg1_val[22]),
    .B(net265),
    .X(_05895_));
 sky130_fd_sc_hd__nand2_4 _12751_ (.A(_05894_),
    .B(_05895_),
    .Y(_05896_));
 sky130_fd_sc_hd__o21a_2 _12752_ (.A1(_05890_),
    .A2(_05893_),
    .B1(_05891_),
    .X(_05897_));
 sky130_fd_sc_hd__xor2_4 _12753_ (.A(_05896_),
    .B(_05897_),
    .X(loadstore_address[22]));
 sky130_fd_sc_hd__o21ai_4 _12754_ (.A1(_05896_),
    .A2(_05897_),
    .B1(_05894_),
    .Y(_05899_));
 sky130_fd_sc_hd__xnor2_4 _12755_ (.A(reg1_val[23]),
    .B(net265),
    .Y(_05900_));
 sky130_fd_sc_hd__xnor2_4 _12756_ (.A(_05899_),
    .B(_05900_),
    .Y(loadstore_address[23]));
 sky130_fd_sc_hd__nand2_1 _12757_ (.A(reg1_val[24]),
    .B(net266),
    .Y(_05901_));
 sky130_fd_sc_hd__or2_1 _12758_ (.A(reg1_val[24]),
    .B(net266),
    .X(_05902_));
 sky130_fd_sc_hd__nand2_2 _12759_ (.A(_05901_),
    .B(_05902_),
    .Y(_05903_));
 sky130_fd_sc_hd__or4_1 _12760_ (.A(_05884_),
    .B(_05892_),
    .C(_05896_),
    .D(_05900_),
    .X(_05904_));
 sky130_fd_sc_hd__a2bb2o_2 _12761_ (.A1_N(_05885_),
    .A2_N(_05904_),
    .B1(net265),
    .B2(_00232_),
    .X(_05905_));
 sky130_fd_sc_hd__nand2b_1 _12762_ (.A_N(_05903_),
    .B(_05905_),
    .Y(_05906_));
 sky130_fd_sc_hd__xnor2_4 _12763_ (.A(_05903_),
    .B(_05905_),
    .Y(loadstore_address[24]));
 sky130_fd_sc_hd__nand2_2 _12764_ (.A(_05901_),
    .B(_05906_),
    .Y(_05908_));
 sky130_fd_sc_hd__xnor2_4 _12765_ (.A(reg1_val[25]),
    .B(net266),
    .Y(_05909_));
 sky130_fd_sc_hd__xnor2_4 _12766_ (.A(_05908_),
    .B(_05909_),
    .Y(loadstore_address[25]));
 sky130_fd_sc_hd__and2_1 _12767_ (.A(reg1_val[26]),
    .B(net266),
    .X(_05910_));
 sky130_fd_sc_hd__or2_1 _12768_ (.A(reg1_val[26]),
    .B(net266),
    .X(_05911_));
 sky130_fd_sc_hd__nand2b_2 _12769_ (.A_N(_05910_),
    .B(_05911_),
    .Y(_05912_));
 sky130_fd_sc_hd__or2_1 _12770_ (.A(_05906_),
    .B(_05909_),
    .X(_05913_));
 sky130_fd_sc_hd__a21bo_2 _12771_ (.A1(net266),
    .A2(_00234_),
    .B1_N(_05913_),
    .X(_05914_));
 sky130_fd_sc_hd__xnor2_4 _12772_ (.A(_05912_),
    .B(_05914_),
    .Y(loadstore_address[26]));
 sky130_fd_sc_hd__a21o_1 _12773_ (.A1(_05911_),
    .A2(_05914_),
    .B1(_05910_),
    .X(_05915_));
 sky130_fd_sc_hd__xnor2_4 _12774_ (.A(reg1_val[27]),
    .B(net266),
    .Y(_05917_));
 sky130_fd_sc_hd__xnor2_4 _12775_ (.A(_05915_),
    .B(_05917_),
    .Y(loadstore_address[27]));
 sky130_fd_sc_hd__and2_1 _12776_ (.A(reg1_val[28]),
    .B(net266),
    .X(_05918_));
 sky130_fd_sc_hd__nor2_1 _12777_ (.A(reg1_val[28]),
    .B(net266),
    .Y(_05919_));
 sky130_fd_sc_hd__or2_1 _12778_ (.A(_05918_),
    .B(_05919_),
    .X(_05920_));
 sky130_fd_sc_hd__nand2_1 _12779_ (.A(net266),
    .B(_00449_),
    .Y(_05921_));
 sky130_fd_sc_hd__or3_1 _12780_ (.A(_05912_),
    .B(_05913_),
    .C(_05917_),
    .X(_05922_));
 sky130_fd_sc_hd__a21oi_2 _12781_ (.A1(_05921_),
    .A2(_05922_),
    .B1(_05920_),
    .Y(_05923_));
 sky130_fd_sc_hd__and3_2 _12782_ (.A(_05920_),
    .B(_05921_),
    .C(_05922_),
    .X(_05924_));
 sky130_fd_sc_hd__nor2_8 _12783_ (.A(_05923_),
    .B(_05924_),
    .Y(loadstore_address[28]));
 sky130_fd_sc_hd__or2_1 _12784_ (.A(reg1_val[29]),
    .B(net266),
    .X(_05926_));
 sky130_fd_sc_hd__nand2_1 _12785_ (.A(reg1_val[29]),
    .B(net266),
    .Y(_05927_));
 sky130_fd_sc_hd__nand2_2 _12786_ (.A(_05926_),
    .B(_05927_),
    .Y(_05928_));
 sky130_fd_sc_hd__or2_2 _12787_ (.A(_05918_),
    .B(_05923_),
    .X(_05929_));
 sky130_fd_sc_hd__xnor2_4 _12788_ (.A(_05928_),
    .B(_05929_),
    .Y(loadstore_address[29]));
 sky130_fd_sc_hd__and2_1 _12789_ (.A(reg1_val[30]),
    .B(net266),
    .X(_05930_));
 sky130_fd_sc_hd__or2_1 _12790_ (.A(reg1_val[30]),
    .B(net266),
    .X(_05931_));
 sky130_fd_sc_hd__nand2b_2 _12791_ (.A_N(_05930_),
    .B(_05931_),
    .Y(_05932_));
 sky130_fd_sc_hd__a21bo_2 _12792_ (.A1(_05926_),
    .A2(_05929_),
    .B1_N(_05927_),
    .X(_05933_));
 sky130_fd_sc_hd__xnor2_4 _12793_ (.A(_05932_),
    .B(_05933_),
    .Y(loadstore_address[30]));
 sky130_fd_sc_hd__a21oi_1 _12794_ (.A1(_05931_),
    .A2(_05933_),
    .B1(_05930_),
    .Y(_05935_));
 sky130_fd_sc_hd__xnor2_2 _12795_ (.A(_04531_),
    .B(_05935_),
    .Y(_05936_));
 sky130_fd_sc_hd__xnor2_4 _12796_ (.A(_04795_),
    .B(_05936_),
    .Y(loadstore_address[31]));
 sky130_fd_sc_hd__nand2_1 _12797_ (.A(net462),
    .B(net435),
    .Y(_05937_));
 sky130_fd_sc_hd__nand3_1 _12798_ (.A(net422),
    .B(net462),
    .C(net435),
    .Y(_05938_));
 sky130_fd_sc_hd__and4_1 _12799_ (.A(net361),
    .B(net495),
    .C(net593),
    .D(\div_counter[0] ),
    .X(_05939_));
 sky130_fd_sc_hd__inv_2 _12800_ (.A(net362),
    .Y(_05940_));
 sky130_fd_sc_hd__nand2_1 _12801_ (.A(net298),
    .B(net362),
    .Y(_05941_));
 sky130_fd_sc_hd__nor2_1 _12802_ (.A(net254),
    .B(net363),
    .Y(_05942_));
 sky130_fd_sc_hd__nor3_1 _12803_ (.A(rst),
    .B(_06465_),
    .C(_05942_),
    .Y(_00000_));
 sky130_fd_sc_hd__nor2_2 _12804_ (.A(net256),
    .B(_06464_),
    .Y(_05944_));
 sky130_fd_sc_hd__nand2_4 _12805_ (.A(net254),
    .B(_06463_),
    .Y(_05945_));
 sky130_fd_sc_hd__or2_1 _12806_ (.A(net304),
    .B(net175),
    .X(_05946_));
 sky130_fd_sc_hd__o211a_1 _12807_ (.A1(_02078_),
    .A2(net171),
    .B1(net305),
    .C1(net282),
    .X(_00001_));
 sky130_fd_sc_hd__nand2_1 _12808_ (.A(net216),
    .B(net172),
    .Y(_05947_));
 sky130_fd_sc_hd__o211a_1 _12809_ (.A1(net306),
    .A2(net172),
    .B1(_05947_),
    .C1(net280),
    .X(_00002_));
 sky130_fd_sc_hd__or2_1 _12810_ (.A(net449),
    .B(net172),
    .X(_05948_));
 sky130_fd_sc_hd__o211a_1 _12811_ (.A1(_00240_),
    .A2(net168),
    .B1(net450),
    .C1(net280),
    .X(_00003_));
 sky130_fd_sc_hd__or2_1 _12812_ (.A(net365),
    .B(net172),
    .X(_05949_));
 sky130_fd_sc_hd__o211a_1 _12813_ (.A1(_00265_),
    .A2(net168),
    .B1(net366),
    .C1(net279),
    .X(_00004_));
 sky130_fd_sc_hd__or2_1 _12814_ (.A(net387),
    .B(net172),
    .X(_05951_));
 sky130_fd_sc_hd__o211a_1 _12815_ (.A1(_00258_),
    .A2(net168),
    .B1(net388),
    .C1(net279),
    .X(_00005_));
 sky130_fd_sc_hd__or2_1 _12816_ (.A(net406),
    .B(_05944_),
    .X(_05952_));
 sky130_fd_sc_hd__o211a_1 _12817_ (.A1(_00226_),
    .A2(_05945_),
    .B1(net407),
    .C1(net279),
    .X(_00006_));
 sky130_fd_sc_hd__or2_1 _12818_ (.A(net349),
    .B(net172),
    .X(_05953_));
 sky130_fd_sc_hd__o211a_1 _12819_ (.A1(_00213_),
    .A2(net168),
    .B1(net350),
    .C1(net279),
    .X(_00007_));
 sky130_fd_sc_hd__or2_1 _12820_ (.A(net313),
    .B(net172),
    .X(_05954_));
 sky130_fd_sc_hd__o211a_1 _12821_ (.A1(_00374_),
    .A2(net168),
    .B1(net314),
    .C1(net279),
    .X(_00008_));
 sky130_fd_sc_hd__or2_1 _12822_ (.A(net341),
    .B(net173),
    .X(_05955_));
 sky130_fd_sc_hd__o211a_1 _12823_ (.A1(net113),
    .A2(net168),
    .B1(net342),
    .C1(net279),
    .X(_00009_));
 sky130_fd_sc_hd__or2_1 _12824_ (.A(net325),
    .B(net173),
    .X(_05957_));
 sky130_fd_sc_hd__o211a_1 _12825_ (.A1(_00308_),
    .A2(net169),
    .B1(net326),
    .C1(net283),
    .X(_00010_));
 sky130_fd_sc_hd__or2_1 _12826_ (.A(net327),
    .B(net173),
    .X(_05958_));
 sky130_fd_sc_hd__o211a_1 _12827_ (.A1(_00330_),
    .A2(net168),
    .B1(net328),
    .C1(net279),
    .X(_00011_));
 sky130_fd_sc_hd__or2_1 _12828_ (.A(net317),
    .B(net175),
    .X(_05959_));
 sky130_fd_sc_hd__o211a_1 _12829_ (.A1(_00324_),
    .A2(net171),
    .B1(net318),
    .C1(net282),
    .X(_00012_));
 sky130_fd_sc_hd__or2_1 _12830_ (.A(net380),
    .B(net174),
    .X(_05960_));
 sky130_fd_sc_hd__o211a_1 _12831_ (.A1(_00291_),
    .A2(net170),
    .B1(net381),
    .C1(net282),
    .X(_00013_));
 sky130_fd_sc_hd__or2_1 _12832_ (.A(net389),
    .B(net174),
    .X(_05961_));
 sky130_fd_sc_hd__o211a_1 _12833_ (.A1(_00287_),
    .A2(net170),
    .B1(net390),
    .C1(net277),
    .X(_00014_));
 sky130_fd_sc_hd__or2_1 _12834_ (.A(net401),
    .B(net174),
    .X(_05963_));
 sky130_fd_sc_hd__o211a_1 _12835_ (.A1(_00366_),
    .A2(net170),
    .B1(net402),
    .C1(net276),
    .X(_00015_));
 sky130_fd_sc_hd__or2_1 _12836_ (.A(net345),
    .B(net174),
    .X(_05964_));
 sky130_fd_sc_hd__o211a_1 _12837_ (.A1(_00361_),
    .A2(net170),
    .B1(net346),
    .C1(net276),
    .X(_00016_));
 sky130_fd_sc_hd__or2_1 _12838_ (.A(net315),
    .B(net174),
    .X(_05965_));
 sky130_fd_sc_hd__o211a_1 _12839_ (.A1(_00354_),
    .A2(net170),
    .B1(net316),
    .C1(net276),
    .X(_00017_));
 sky130_fd_sc_hd__or2_1 _12840_ (.A(net331),
    .B(net174),
    .X(_05966_));
 sky130_fd_sc_hd__o211a_1 _12841_ (.A1(_00348_),
    .A2(net170),
    .B1(net332),
    .C1(net274),
    .X(_00018_));
 sky130_fd_sc_hd__or2_1 _12842_ (.A(net382),
    .B(net174),
    .X(_05967_));
 sky130_fd_sc_hd__o211a_1 _12843_ (.A1(_00189_),
    .A2(net170),
    .B1(net383),
    .C1(net274),
    .X(_00019_));
 sky130_fd_sc_hd__or2_1 _12844_ (.A(net416),
    .B(net174),
    .X(_05969_));
 sky130_fd_sc_hd__o211a_1 _12845_ (.A1(_00179_),
    .A2(net170),
    .B1(net417),
    .C1(net274),
    .X(_00020_));
 sky130_fd_sc_hd__or2_1 _12846_ (.A(net391),
    .B(net174),
    .X(_05970_));
 sky130_fd_sc_hd__o211a_1 _12847_ (.A1(_00172_),
    .A2(net170),
    .B1(net392),
    .C1(net275),
    .X(_00021_));
 sky130_fd_sc_hd__or2_1 _12848_ (.A(net347),
    .B(net174),
    .X(_05971_));
 sky130_fd_sc_hd__o211a_1 _12849_ (.A1(_00163_),
    .A2(net170),
    .B1(net348),
    .C1(net274),
    .X(_00022_));
 sky130_fd_sc_hd__or2_1 _12850_ (.A(net329),
    .B(net174),
    .X(_05972_));
 sky130_fd_sc_hd__o211a_1 _12851_ (.A1(_06547_),
    .A2(net170),
    .B1(net330),
    .C1(net274),
    .X(_00023_));
 sky130_fd_sc_hd__or2_1 _12852_ (.A(net357),
    .B(net174),
    .X(_05973_));
 sky130_fd_sc_hd__o211a_1 _12853_ (.A1(_06540_),
    .A2(net170),
    .B1(net358),
    .C1(net274),
    .X(_00024_));
 sky130_fd_sc_hd__or2_1 _12854_ (.A(net319),
    .B(net174),
    .X(_05975_));
 sky130_fd_sc_hd__o211a_1 _12855_ (.A1(_06563_),
    .A2(net170),
    .B1(net320),
    .C1(net276),
    .X(_00025_));
 sky130_fd_sc_hd__or2_1 _12856_ (.A(net372),
    .B(net175),
    .X(_05976_));
 sky130_fd_sc_hd__o211a_1 _12857_ (.A1(_06559_),
    .A2(net170),
    .B1(net373),
    .C1(net276),
    .X(_00026_));
 sky130_fd_sc_hd__or2_1 _12858_ (.A(net359),
    .B(net174),
    .X(_05977_));
 sky130_fd_sc_hd__o211a_1 _12859_ (.A1(_06525_),
    .A2(net171),
    .B1(net360),
    .C1(net276),
    .X(_00027_));
 sky130_fd_sc_hd__or2_1 _12860_ (.A(net339),
    .B(net174),
    .X(_05978_));
 sky130_fd_sc_hd__o211a_1 _12861_ (.A1(_06517_),
    .A2(net170),
    .B1(net340),
    .C1(net276),
    .X(_00028_));
 sky130_fd_sc_hd__or2_1 _12862_ (.A(net355),
    .B(net174),
    .X(_05979_));
 sky130_fd_sc_hd__o211a_1 _12863_ (.A1(_00143_),
    .A2(net170),
    .B1(net356),
    .C1(net282),
    .X(_00029_));
 sky130_fd_sc_hd__or2_1 _12864_ (.A(net353),
    .B(net175),
    .X(_05981_));
 sky130_fd_sc_hd__o211a_1 _12865_ (.A1(_00408_),
    .A2(net171),
    .B1(net354),
    .C1(net282),
    .X(_00030_));
 sky130_fd_sc_hd__or2_1 _12866_ (.A(net323),
    .B(net175),
    .X(_05982_));
 sky130_fd_sc_hd__o211a_1 _12867_ (.A1(_00700_),
    .A2(net171),
    .B1(net324),
    .C1(net282),
    .X(_00031_));
 sky130_fd_sc_hd__or2_1 _12868_ (.A(net321),
    .B(net175),
    .X(_05983_));
 sky130_fd_sc_hd__o211a_1 _12869_ (.A1(_01951_),
    .A2(net171),
    .B1(net322),
    .C1(net282),
    .X(_00032_));
 sky130_fd_sc_hd__or2_1 _12870_ (.A(net343),
    .B(net175),
    .X(_05984_));
 sky130_fd_sc_hd__o211a_1 _12871_ (.A1(_02066_),
    .A2(net171),
    .B1(net344),
    .C1(net282),
    .X(_00033_));
 sky130_fd_sc_hd__and2b_1 _12872_ (.A_N(net321),
    .B(\div_shifter[61] ),
    .X(_05985_));
 sky130_fd_sc_hd__and2b_1 _12873_ (.A_N(\div_shifter[61] ),
    .B(net321),
    .X(_05986_));
 sky130_fd_sc_hd__nor2_1 _12874_ (.A(_05985_),
    .B(_05986_),
    .Y(_05988_));
 sky130_fd_sc_hd__nand2b_1 _12875_ (.A_N(\div_shifter[60] ),
    .B(net323),
    .Y(_05989_));
 sky130_fd_sc_hd__and2b_1 _12876_ (.A_N(net353),
    .B(net577),
    .X(_05990_));
 sky130_fd_sc_hd__nand2b_1 _12877_ (.A_N(net579),
    .B(net355),
    .Y(_05991_));
 sky130_fd_sc_hd__and2b_1 _12878_ (.A_N(net339),
    .B(net571),
    .X(_05992_));
 sky130_fd_sc_hd__nand2b_1 _12879_ (.A_N(net571),
    .B(net339),
    .Y(_05993_));
 sky130_fd_sc_hd__nand2b_1 _12880_ (.A_N(_05992_),
    .B(_05993_),
    .Y(_05994_));
 sky130_fd_sc_hd__nand2b_1 _12881_ (.A_N(net573),
    .B(net359),
    .Y(_05995_));
 sky130_fd_sc_hd__and2b_1 _12882_ (.A_N(net372),
    .B(net549),
    .X(_05996_));
 sky130_fd_sc_hd__nand2b_1 _12883_ (.A_N(net561),
    .B(net319),
    .Y(_05997_));
 sky130_fd_sc_hd__and2b_1 _12884_ (.A_N(net357),
    .B(\div_shifter[53] ),
    .X(_05999_));
 sky130_fd_sc_hd__nand2b_1 _12885_ (.A_N(\div_shifter[52] ),
    .B(net329),
    .Y(_06000_));
 sky130_fd_sc_hd__and2b_1 _12886_ (.A_N(net347),
    .B(net557),
    .X(_06001_));
 sky130_fd_sc_hd__nand2b_1 _12887_ (.A_N(net559),
    .B(net391),
    .Y(_06002_));
 sky130_fd_sc_hd__and2b_1 _12888_ (.A_N(net416),
    .B(net541),
    .X(_06003_));
 sky130_fd_sc_hd__nand2b_1 _12889_ (.A_N(net541),
    .B(net416),
    .Y(_06004_));
 sky130_fd_sc_hd__nand2b_1 _12890_ (.A_N(\div_shifter[48] ),
    .B(net382),
    .Y(_06005_));
 sky130_fd_sc_hd__nand2b_1 _12891_ (.A_N(net570),
    .B(net331),
    .Y(_06006_));
 sky130_fd_sc_hd__nand2b_1 _12892_ (.A_N(net567),
    .B(net315),
    .Y(_06007_));
 sky130_fd_sc_hd__nand2b_1 _12893_ (.A_N(net565),
    .B(net345),
    .Y(_06008_));
 sky130_fd_sc_hd__nand2b_1 _12894_ (.A_N(\div_shifter[44] ),
    .B(net401),
    .Y(_06010_));
 sky130_fd_sc_hd__nand2b_1 _12895_ (.A_N(\div_shifter[43] ),
    .B(net389),
    .Y(_06011_));
 sky130_fd_sc_hd__nand2b_1 _12896_ (.A_N(net574),
    .B(net380),
    .Y(_06012_));
 sky130_fd_sc_hd__nand2b_1 _12897_ (.A_N(\div_shifter[41] ),
    .B(net317),
    .Y(_06013_));
 sky130_fd_sc_hd__nand2b_1 _12898_ (.A_N(net547),
    .B(net327),
    .Y(_06014_));
 sky130_fd_sc_hd__nand2b_1 _12899_ (.A_N(net576),
    .B(net325),
    .Y(_06015_));
 sky130_fd_sc_hd__nand2b_1 _12900_ (.A_N(net555),
    .B(net341),
    .Y(_06016_));
 sky130_fd_sc_hd__nand2b_1 _12901_ (.A_N(net543),
    .B(net313),
    .Y(_06017_));
 sky130_fd_sc_hd__and2b_1 _12902_ (.A_N(net349),
    .B(\div_shifter[36] ),
    .X(_06018_));
 sky130_fd_sc_hd__nand2b_1 _12903_ (.A_N(\div_shifter[36] ),
    .B(net349),
    .Y(_06019_));
 sky130_fd_sc_hd__nand2b_1 _12904_ (.A_N(_06018_),
    .B(_06019_),
    .Y(_06021_));
 sky130_fd_sc_hd__and2b_1 _12905_ (.A_N(net406),
    .B(net551),
    .X(_06022_));
 sky130_fd_sc_hd__nand2b_1 _12906_ (.A_N(net551),
    .B(net406),
    .Y(_06023_));
 sky130_fd_sc_hd__nand2b_1 _12907_ (.A_N(_06022_),
    .B(_06023_),
    .Y(_06024_));
 sky130_fd_sc_hd__nand2b_1 _12908_ (.A_N(\div_shifter[34] ),
    .B(net387),
    .Y(_06025_));
 sky130_fd_sc_hd__nand2b_1 _12909_ (.A_N(net530),
    .B(net365),
    .Y(_06026_));
 sky130_fd_sc_hd__and2b_1 _12910_ (.A_N(net449),
    .B(net540),
    .X(_06027_));
 sky130_fd_sc_hd__xnor2_1 _12911_ (.A(net540),
    .B(net449),
    .Y(_06028_));
 sky130_fd_sc_hd__nand2b_1 _12912_ (.A_N(net311),
    .B(net306),
    .Y(_06029_));
 sky130_fd_sc_hd__a21o_1 _12913_ (.A1(_06028_),
    .A2(_06029_),
    .B1(_06027_),
    .X(_06030_));
 sky130_fd_sc_hd__nand2b_1 _12914_ (.A_N(net365),
    .B(net530),
    .Y(_06032_));
 sky130_fd_sc_hd__a21bo_1 _12915_ (.A1(_06026_),
    .A2(_06030_),
    .B1_N(_06032_),
    .X(_06033_));
 sky130_fd_sc_hd__nand2b_1 _12916_ (.A_N(net387),
    .B(\div_shifter[34] ),
    .Y(_06034_));
 sky130_fd_sc_hd__a21bo_1 _12917_ (.A1(_06025_),
    .A2(_06033_),
    .B1_N(_06034_),
    .X(_06035_));
 sky130_fd_sc_hd__a21o_1 _12918_ (.A1(_06023_),
    .A2(_06035_),
    .B1(_06022_),
    .X(_06036_));
 sky130_fd_sc_hd__a21o_1 _12919_ (.A1(_06019_),
    .A2(_06036_),
    .B1(_06018_),
    .X(_06037_));
 sky130_fd_sc_hd__nand2b_1 _12920_ (.A_N(net313),
    .B(net543),
    .Y(_06038_));
 sky130_fd_sc_hd__a21bo_1 _12921_ (.A1(_06017_),
    .A2(_06037_),
    .B1_N(_06038_),
    .X(_06039_));
 sky130_fd_sc_hd__nand2b_1 _12922_ (.A_N(net341),
    .B(net555),
    .Y(_06040_));
 sky130_fd_sc_hd__a21bo_1 _12923_ (.A1(_06016_),
    .A2(_06039_),
    .B1_N(_06040_),
    .X(_06041_));
 sky130_fd_sc_hd__nand2b_1 _12924_ (.A_N(net325),
    .B(net576),
    .Y(_06043_));
 sky130_fd_sc_hd__a21bo_1 _12925_ (.A1(_06015_),
    .A2(_06041_),
    .B1_N(_06043_),
    .X(_06044_));
 sky130_fd_sc_hd__nand2b_1 _12926_ (.A_N(net327),
    .B(net547),
    .Y(_06045_));
 sky130_fd_sc_hd__a21bo_1 _12927_ (.A1(_06014_),
    .A2(_06044_),
    .B1_N(_06045_),
    .X(_06046_));
 sky130_fd_sc_hd__nand2b_1 _12928_ (.A_N(net317),
    .B(\div_shifter[41] ),
    .Y(_06047_));
 sky130_fd_sc_hd__a21bo_1 _12929_ (.A1(_06013_),
    .A2(_06046_),
    .B1_N(_06047_),
    .X(_06048_));
 sky130_fd_sc_hd__nand2b_1 _12930_ (.A_N(net380),
    .B(net574),
    .Y(_06049_));
 sky130_fd_sc_hd__a21bo_1 _12931_ (.A1(_06012_),
    .A2(_06048_),
    .B1_N(_06049_),
    .X(_06050_));
 sky130_fd_sc_hd__nand2b_1 _12932_ (.A_N(net389),
    .B(\div_shifter[43] ),
    .Y(_06051_));
 sky130_fd_sc_hd__a21bo_1 _12933_ (.A1(_06011_),
    .A2(_06050_),
    .B1_N(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__nand2b_1 _12934_ (.A_N(net401),
    .B(\div_shifter[44] ),
    .Y(_06054_));
 sky130_fd_sc_hd__a21bo_1 _12935_ (.A1(_06010_),
    .A2(_06052_),
    .B1_N(_06054_),
    .X(_06055_));
 sky130_fd_sc_hd__nand2b_1 _12936_ (.A_N(net345),
    .B(net565),
    .Y(_06056_));
 sky130_fd_sc_hd__a21bo_1 _12937_ (.A1(_06008_),
    .A2(_06055_),
    .B1_N(_06056_),
    .X(_06057_));
 sky130_fd_sc_hd__nand2b_1 _12938_ (.A_N(net315),
    .B(net567),
    .Y(_06058_));
 sky130_fd_sc_hd__a21bo_1 _12939_ (.A1(_06007_),
    .A2(_06057_),
    .B1_N(_06058_),
    .X(_06059_));
 sky130_fd_sc_hd__nand2b_1 _12940_ (.A_N(net331),
    .B(net570),
    .Y(_06060_));
 sky130_fd_sc_hd__a21bo_1 _12941_ (.A1(_06006_),
    .A2(_06059_),
    .B1_N(_06060_),
    .X(_06061_));
 sky130_fd_sc_hd__nand2b_1 _12942_ (.A_N(net382),
    .B(\div_shifter[48] ),
    .Y(_06062_));
 sky130_fd_sc_hd__a21bo_1 _12943_ (.A1(_06005_),
    .A2(_06061_),
    .B1_N(_06062_),
    .X(_06063_));
 sky130_fd_sc_hd__a21o_1 _12944_ (.A1(_06004_),
    .A2(_06063_),
    .B1(_06003_),
    .X(_06065_));
 sky130_fd_sc_hd__nand2b_1 _12945_ (.A_N(net391),
    .B(net559),
    .Y(_06066_));
 sky130_fd_sc_hd__a21bo_1 _12946_ (.A1(_06002_),
    .A2(_06065_),
    .B1_N(_06066_),
    .X(_06067_));
 sky130_fd_sc_hd__nand2b_1 _12947_ (.A_N(net557),
    .B(net347),
    .Y(_06068_));
 sky130_fd_sc_hd__nand2b_1 _12948_ (.A_N(_06001_),
    .B(_06068_),
    .Y(_06069_));
 sky130_fd_sc_hd__a21o_1 _12949_ (.A1(_06067_),
    .A2(_06068_),
    .B1(_06001_),
    .X(_06070_));
 sky130_fd_sc_hd__nand2b_1 _12950_ (.A_N(net329),
    .B(\div_shifter[52] ),
    .Y(_06071_));
 sky130_fd_sc_hd__a21bo_1 _12951_ (.A1(_06000_),
    .A2(_06070_),
    .B1_N(_06071_),
    .X(_06072_));
 sky130_fd_sc_hd__nand2b_1 _12952_ (.A_N(\div_shifter[53] ),
    .B(net357),
    .Y(_06073_));
 sky130_fd_sc_hd__nand2b_1 _12953_ (.A_N(_05999_),
    .B(_06073_),
    .Y(_06074_));
 sky130_fd_sc_hd__a21o_1 _12954_ (.A1(_06072_),
    .A2(_06073_),
    .B1(_05999_),
    .X(_06076_));
 sky130_fd_sc_hd__nand2b_1 _12955_ (.A_N(net319),
    .B(net561),
    .Y(_06077_));
 sky130_fd_sc_hd__a21bo_1 _12956_ (.A1(_05997_),
    .A2(_06076_),
    .B1_N(_06077_),
    .X(_06078_));
 sky130_fd_sc_hd__nand2b_1 _12957_ (.A_N(net549),
    .B(net372),
    .Y(_06079_));
 sky130_fd_sc_hd__nand2b_1 _12958_ (.A_N(_05996_),
    .B(_06079_),
    .Y(_06080_));
 sky130_fd_sc_hd__a21o_1 _12959_ (.A1(_06078_),
    .A2(_06079_),
    .B1(_05996_),
    .X(_06081_));
 sky130_fd_sc_hd__nand2b_1 _12960_ (.A_N(net359),
    .B(net573),
    .Y(_06082_));
 sky130_fd_sc_hd__a21bo_1 _12961_ (.A1(_05995_),
    .A2(_06081_),
    .B1_N(_06082_),
    .X(_06083_));
 sky130_fd_sc_hd__a21o_1 _12962_ (.A1(_05993_),
    .A2(_06083_),
    .B1(_05992_),
    .X(_06084_));
 sky130_fd_sc_hd__nand2b_1 _12963_ (.A_N(net355),
    .B(net579),
    .Y(_06085_));
 sky130_fd_sc_hd__a21bo_1 _12964_ (.A1(_05991_),
    .A2(_06084_),
    .B1_N(_06085_),
    .X(_06087_));
 sky130_fd_sc_hd__nand2b_1 _12965_ (.A_N(net577),
    .B(net353),
    .Y(_06088_));
 sky130_fd_sc_hd__nand2b_1 _12966_ (.A_N(_05990_),
    .B(_06088_),
    .Y(_06089_));
 sky130_fd_sc_hd__a21o_1 _12967_ (.A1(_06087_),
    .A2(_06088_),
    .B1(_05990_),
    .X(_06090_));
 sky130_fd_sc_hd__nand2b_1 _12968_ (.A_N(net323),
    .B(\div_shifter[60] ),
    .Y(_06091_));
 sky130_fd_sc_hd__a21boi_1 _12969_ (.A1(_05989_),
    .A2(_06090_),
    .B1_N(_06091_),
    .Y(_06092_));
 sky130_fd_sc_hd__o21ba_1 _12970_ (.A1(_05986_),
    .A2(_06092_),
    .B1_N(_05985_),
    .X(_06093_));
 sky130_fd_sc_hd__nor2_1 _12971_ (.A(net343),
    .B(_06093_),
    .Y(_06094_));
 sky130_fd_sc_hd__a21boi_1 _12972_ (.A1(net343),
    .A2(_06093_),
    .B1_N(net545),
    .Y(_06095_));
 sky130_fd_sc_hd__or2_2 _12973_ (.A(_06094_),
    .B(_06095_),
    .X(_06096_));
 sky130_fd_sc_hd__a22o_1 _12974_ (.A1(net588),
    .A2(net188),
    .B1(net2),
    .B2(net257),
    .X(_06098_));
 sky130_fd_sc_hd__and2_1 _12975_ (.A(net278),
    .B(_06098_),
    .X(_00034_));
 sky130_fd_sc_hd__a22o_1 _12976_ (.A1(\div_res[0] ),
    .A2(net257),
    .B1(net188),
    .B2(net538),
    .X(_06099_));
 sky130_fd_sc_hd__and2_1 _12977_ (.A(net278),
    .B(net539),
    .X(_00035_));
 sky130_fd_sc_hd__a22o_1 _12978_ (.A1(net596),
    .A2(net257),
    .B1(net188),
    .B2(net532),
    .X(_06100_));
 sky130_fd_sc_hd__and2_1 _12979_ (.A(net278),
    .B(net533),
    .X(_00036_));
 sky130_fd_sc_hd__a22o_1 _12980_ (.A1(\div_res[2] ),
    .A2(net257),
    .B1(net188),
    .B2(net516),
    .X(_06101_));
 sky130_fd_sc_hd__and2_1 _12981_ (.A(net278),
    .B(net517),
    .X(_00037_));
 sky130_fd_sc_hd__a22o_1 _12982_ (.A1(net516),
    .A2(net257),
    .B1(net188),
    .B2(net534),
    .X(_06102_));
 sky130_fd_sc_hd__and2_1 _12983_ (.A(net278),
    .B(net535),
    .X(_00038_));
 sky130_fd_sc_hd__a22o_1 _12984_ (.A1(net595),
    .A2(net257),
    .B1(net188),
    .B2(net491),
    .X(_06104_));
 sky130_fd_sc_hd__and2_1 _12985_ (.A(net278),
    .B(net492),
    .X(_00039_));
 sky130_fd_sc_hd__a22o_1 _12986_ (.A1(net491),
    .A2(net257),
    .B1(net188),
    .B2(net506),
    .X(_06105_));
 sky130_fd_sc_hd__and2_1 _12987_ (.A(net278),
    .B(net507),
    .X(_00040_));
 sky130_fd_sc_hd__a22o_1 _12988_ (.A1(net506),
    .A2(net257),
    .B1(net188),
    .B2(net510),
    .X(_06106_));
 sky130_fd_sc_hd__and2_1 _12989_ (.A(net278),
    .B(net511),
    .X(_00041_));
 sky130_fd_sc_hd__a22o_1 _12990_ (.A1(net510),
    .A2(net257),
    .B1(net188),
    .B2(net512),
    .X(_06107_));
 sky130_fd_sc_hd__and2_1 _12991_ (.A(net278),
    .B(net513),
    .X(_00042_));
 sky130_fd_sc_hd__a22o_1 _12992_ (.A1(\div_res[8] ),
    .A2(net257),
    .B1(net188),
    .B2(net503),
    .X(_06108_));
 sky130_fd_sc_hd__and2_1 _12993_ (.A(net278),
    .B(net504),
    .X(_00043_));
 sky130_fd_sc_hd__a22o_1 _12994_ (.A1(net503),
    .A2(net257),
    .B1(net188),
    .B2(net508),
    .X(_06110_));
 sky130_fd_sc_hd__and2_1 _12995_ (.A(net278),
    .B(net509),
    .X(_00044_));
 sky130_fd_sc_hd__a22o_1 _12996_ (.A1(\div_res[10] ),
    .A2(net257),
    .B1(net188),
    .B2(net480),
    .X(_06111_));
 sky130_fd_sc_hd__and2_1 _12997_ (.A(net278),
    .B(net481),
    .X(_00045_));
 sky130_fd_sc_hd__a22o_1 _12998_ (.A1(net480),
    .A2(net257),
    .B1(net188),
    .B2(net464),
    .X(_06112_));
 sky130_fd_sc_hd__and2_1 _12999_ (.A(net278),
    .B(net494),
    .X(_00046_));
 sky130_fd_sc_hd__a22o_1 _13000_ (.A1(net464),
    .A2(net257),
    .B1(net188),
    .B2(\div_res[13] ),
    .X(_06113_));
 sky130_fd_sc_hd__and2_1 _13001_ (.A(net278),
    .B(net465),
    .X(_00047_));
 sky130_fd_sc_hd__a22o_1 _13002_ (.A1(\div_res[13] ),
    .A2(net258),
    .B1(net189),
    .B2(net488),
    .X(_06114_));
 sky130_fd_sc_hd__and2_1 _13003_ (.A(net275),
    .B(net489),
    .X(_00048_));
 sky130_fd_sc_hd__a22o_1 _13004_ (.A1(\div_res[14] ),
    .A2(net258),
    .B1(net189),
    .B2(net477),
    .X(_06116_));
 sky130_fd_sc_hd__and2_1 _13005_ (.A(net275),
    .B(net478),
    .X(_00049_));
 sky130_fd_sc_hd__a22o_1 _13006_ (.A1(net477),
    .A2(net258),
    .B1(net189),
    .B2(net499),
    .X(_06117_));
 sky130_fd_sc_hd__and2_1 _13007_ (.A(net275),
    .B(net500),
    .X(_00050_));
 sky130_fd_sc_hd__a22o_1 _13008_ (.A1(\div_res[16] ),
    .A2(net258),
    .B1(net189),
    .B2(net472),
    .X(_06118_));
 sky130_fd_sc_hd__and2_1 _13009_ (.A(net275),
    .B(net473),
    .X(_00051_));
 sky130_fd_sc_hd__a22o_1 _13010_ (.A1(net472),
    .A2(net258),
    .B1(net189),
    .B2(net475),
    .X(_06119_));
 sky130_fd_sc_hd__and2_1 _13011_ (.A(net274),
    .B(net487),
    .X(_00052_));
 sky130_fd_sc_hd__a22o_1 _13012_ (.A1(net475),
    .A2(net258),
    .B1(net189),
    .B2(net467),
    .X(_06120_));
 sky130_fd_sc_hd__and2_1 _13013_ (.A(net274),
    .B(net476),
    .X(_00053_));
 sky130_fd_sc_hd__a22o_1 _13014_ (.A1(net467),
    .A2(net258),
    .B1(net189),
    .B2(\div_res[20] ),
    .X(_06122_));
 sky130_fd_sc_hd__and2_1 _13015_ (.A(net275),
    .B(net468),
    .X(_00054_));
 sky130_fd_sc_hd__a22o_1 _13016_ (.A1(\div_res[20] ),
    .A2(net258),
    .B1(net189),
    .B2(net483),
    .X(_06123_));
 sky130_fd_sc_hd__and2_1 _13017_ (.A(net275),
    .B(net484),
    .X(_00055_));
 sky130_fd_sc_hd__a22o_1 _13018_ (.A1(net483),
    .A2(net258),
    .B1(net189),
    .B2(net514),
    .X(_06124_));
 sky130_fd_sc_hd__and2_1 _13019_ (.A(net275),
    .B(net515),
    .X(_00056_));
 sky130_fd_sc_hd__a22o_1 _13020_ (.A1(\div_res[22] ),
    .A2(net258),
    .B1(net189),
    .B2(net496),
    .X(_06125_));
 sky130_fd_sc_hd__and2_1 _13021_ (.A(net277),
    .B(net497),
    .X(_00057_));
 sky130_fd_sc_hd__a22o_1 _13022_ (.A1(net496),
    .A2(net258),
    .B1(net189),
    .B2(net457),
    .X(_06126_));
 sky130_fd_sc_hd__and2_1 _13023_ (.A(net276),
    .B(net502),
    .X(_00058_));
 sky130_fd_sc_hd__a22o_1 _13024_ (.A1(net457),
    .A2(net258),
    .B1(net190),
    .B2(\div_res[25] ),
    .X(_06128_));
 sky130_fd_sc_hd__and2_1 _13025_ (.A(net276),
    .B(net458),
    .X(_00059_));
 sky130_fd_sc_hd__a22o_1 _13026_ (.A1(\div_res[25] ),
    .A2(net258),
    .B1(net189),
    .B2(net524),
    .X(_06129_));
 sky130_fd_sc_hd__and2_1 _13027_ (.A(net277),
    .B(net525),
    .X(_00060_));
 sky130_fd_sc_hd__a22o_1 _13028_ (.A1(\div_res[26] ),
    .A2(net259),
    .B1(net189),
    .B2(net519),
    .X(_06130_));
 sky130_fd_sc_hd__and2_1 _13029_ (.A(net277),
    .B(net520),
    .X(_00061_));
 sky130_fd_sc_hd__a22o_1 _13030_ (.A1(net519),
    .A2(net260),
    .B1(net191),
    .B2(net522),
    .X(_06131_));
 sky130_fd_sc_hd__and2_1 _13031_ (.A(net277),
    .B(net523),
    .X(_00062_));
 sky130_fd_sc_hd__a22o_1 _13032_ (.A1(net522),
    .A2(net260),
    .B1(net191),
    .B2(net536),
    .X(_06132_));
 sky130_fd_sc_hd__and2_1 _13033_ (.A(net282),
    .B(net537),
    .X(_00063_));
 sky130_fd_sc_hd__a22o_1 _13034_ (.A1(\div_res[29] ),
    .A2(net260),
    .B1(net191),
    .B2(net527),
    .X(_06134_));
 sky130_fd_sc_hd__and2_1 _13035_ (.A(net283),
    .B(net528),
    .X(_00064_));
 sky130_fd_sc_hd__a22o_1 _13036_ (.A1(\div_res[30] ),
    .A2(net260),
    .B1(net191),
    .B2(net432),
    .X(_06135_));
 sky130_fd_sc_hd__and2_1 _13037_ (.A(net282),
    .B(net433),
    .X(_00065_));
 sky130_fd_sc_hd__a22o_1 _13038_ (.A1(net414),
    .A2(net187),
    .B1(net172),
    .B2(net292),
    .X(_06136_));
 sky130_fd_sc_hd__and2_1 _13039_ (.A(net280),
    .B(net415),
    .X(_00066_));
 sky130_fd_sc_hd__o221a_1 _13040_ (.A1(net414),
    .A2(net253),
    .B1(net185),
    .B2(net420),
    .C1(net280),
    .X(_06137_));
 sky130_fd_sc_hd__o21a_1 _13041_ (.A1(net240),
    .A2(net168),
    .B1(net421),
    .X(_00067_));
 sky130_fd_sc_hd__o221a_1 _13042_ (.A1(net420),
    .A2(net253),
    .B1(net185),
    .B2(net460),
    .C1(net280),
    .X(_06138_));
 sky130_fd_sc_hd__a21boi_1 _13043_ (.A1(_06552_),
    .A2(net172),
    .B1_N(net461),
    .Y(_00068_));
 sky130_fd_sc_hd__a221o_1 _13044_ (.A1(_04454_),
    .A2(net255),
    .B1(net187),
    .B2(net334),
    .C1(rst),
    .X(_06140_));
 sky130_fd_sc_hd__a21oi_1 _13045_ (.A1(net205),
    .A2(net172),
    .B1(net335),
    .Y(_00069_));
 sky130_fd_sc_hd__a221o_1 _13046_ (.A1(net334),
    .A2(net255),
    .B1(net187),
    .B2(net338),
    .C1(rst),
    .X(_06141_));
 sky130_fd_sc_hd__a21oi_1 _13047_ (.A1(_06535_),
    .A2(net172),
    .B1(_06141_),
    .Y(_00070_));
 sky130_fd_sc_hd__a21oi_1 _13048_ (.A1(_04433_),
    .A2(net255),
    .B1(rst),
    .Y(_06142_));
 sky130_fd_sc_hd__o221a_1 _13049_ (.A1(net296),
    .A2(net185),
    .B1(_06532_),
    .B2(net168),
    .C1(_06142_),
    .X(_00071_));
 sky130_fd_sc_hd__o221a_1 _13050_ (.A1(net296),
    .A2(net253),
    .B1(net185),
    .B2(net451),
    .C1(net281),
    .X(_06143_));
 sky130_fd_sc_hd__a21boi_1 _13051_ (.A1(_00157_),
    .A2(net172),
    .B1_N(net452),
    .Y(_00072_));
 sky130_fd_sc_hd__o221a_1 _13052_ (.A1(\div_shifter[6] ),
    .A2(net253),
    .B1(net185),
    .B2(net442),
    .C1(net281),
    .X(_06144_));
 sky130_fd_sc_hd__a21boi_1 _13053_ (.A1(net203),
    .A2(net172),
    .B1_N(net443),
    .Y(_00073_));
 sky130_fd_sc_hd__o221a_1 _13054_ (.A1(net442),
    .A2(net253),
    .B1(net185),
    .B2(net445),
    .C1(net281),
    .X(_06146_));
 sky130_fd_sc_hd__a21boi_1 _13055_ (.A1(_00181_),
    .A2(net172),
    .B1_N(net454),
    .Y(_00074_));
 sky130_fd_sc_hd__o221a_1 _13056_ (.A1(net445),
    .A2(net253),
    .B1(net185),
    .B2(net440),
    .C1(net281),
    .X(_06147_));
 sky130_fd_sc_hd__a21boi_1 _13057_ (.A1(net182),
    .A2(net173),
    .B1_N(net446),
    .Y(_00075_));
 sky130_fd_sc_hd__o221a_1 _13058_ (.A1(net440),
    .A2(net253),
    .B1(net185),
    .B2(net393),
    .C1(net280),
    .X(_06148_));
 sky130_fd_sc_hd__a21boi_1 _13059_ (.A1(_00387_),
    .A2(net173),
    .B1_N(net441),
    .Y(_00076_));
 sky130_fd_sc_hd__o221a_1 _13060_ (.A1(net393),
    .A2(net253),
    .B1(net185),
    .B2(net377),
    .C1(net281),
    .X(_06149_));
 sky130_fd_sc_hd__o21a_1 _13061_ (.A1(_00342_),
    .A2(net168),
    .B1(net394),
    .X(_00077_));
 sky130_fd_sc_hd__o221a_1 _13062_ (.A1(net377),
    .A2(net253),
    .B1(net185),
    .B2(\div_shifter[12] ),
    .C1(net281),
    .X(_06150_));
 sky130_fd_sc_hd__a21boi_1 _13063_ (.A1(_00344_),
    .A2(net173),
    .B1_N(net378),
    .Y(_00078_));
 sky130_fd_sc_hd__o221a_1 _13064_ (.A1(\div_shifter[12] ),
    .A2(net253),
    .B1(net185),
    .B2(net425),
    .C1(net281),
    .X(_06152_));
 sky130_fd_sc_hd__o21a_1 _13065_ (.A1(_00339_),
    .A2(net168),
    .B1(net426),
    .X(_00079_));
 sky130_fd_sc_hd__o221a_1 _13066_ (.A1(net425),
    .A2(net253),
    .B1(net185),
    .B2(net430),
    .C1(net280),
    .X(_06153_));
 sky130_fd_sc_hd__a21boi_1 _13067_ (.A1(_00357_),
    .A2(net173),
    .B1_N(net448),
    .Y(_00080_));
 sky130_fd_sc_hd__o221a_1 _13068_ (.A1(net430),
    .A2(net254),
    .B1(net185),
    .B2(net374),
    .C1(net280),
    .X(_06154_));
 sky130_fd_sc_hd__a21boi_1 _13069_ (.A1(net121),
    .A2(net173),
    .B1_N(net431),
    .Y(_00081_));
 sky130_fd_sc_hd__o221a_1 _13070_ (.A1(net374),
    .A2(net254),
    .B1(net186),
    .B2(\div_shifter[16] ),
    .C1(net280),
    .X(_06155_));
 sky130_fd_sc_hd__a21boi_1 _13071_ (.A1(_00280_),
    .A2(net173),
    .B1_N(net375),
    .Y(_00082_));
 sky130_fd_sc_hd__o221a_1 _13072_ (.A1(\div_shifter[16] ),
    .A2(net254),
    .B1(net186),
    .B2(net395),
    .C1(net280),
    .X(_06156_));
 sky130_fd_sc_hd__o21a_1 _13073_ (.A1(net126),
    .A2(net169),
    .B1(net396),
    .X(_00083_));
 sky130_fd_sc_hd__o221a_1 _13074_ (.A1(net395),
    .A2(net254),
    .B1(net186),
    .B2(net428),
    .C1(net283),
    .X(_06158_));
 sky130_fd_sc_hd__a21boi_1 _13075_ (.A1(_00320_),
    .A2(net173),
    .B1_N(net429),
    .Y(_00084_));
 sky130_fd_sc_hd__o221a_1 _13076_ (.A1(\div_shifter[18] ),
    .A2(net254),
    .B1(net185),
    .B2(net408),
    .C1(net281),
    .X(_06159_));
 sky130_fd_sc_hd__o21a_1 _13077_ (.A1(net89),
    .A2(net168),
    .B1(net409),
    .X(_00085_));
 sky130_fd_sc_hd__o221a_1 _13078_ (.A1(\div_shifter[19] ),
    .A2(net254),
    .B1(net186),
    .B2(net398),
    .C1(net281),
    .X(_06160_));
 sky130_fd_sc_hd__o21a_1 _13079_ (.A1(_00302_),
    .A2(net169),
    .B1(net399),
    .X(_00086_));
 sky130_fd_sc_hd__o221a_1 _13080_ (.A1(\div_shifter[20] ),
    .A2(net254),
    .B1(net186),
    .B2(net384),
    .C1(net281),
    .X(_06161_));
 sky130_fd_sc_hd__o21a_1 _13081_ (.A1(_00216_),
    .A2(net169),
    .B1(net385),
    .X(_00087_));
 sky130_fd_sc_hd__o221a_1 _13082_ (.A1(net384),
    .A2(net253),
    .B1(net186),
    .B2(net418),
    .C1(net283),
    .X(_06162_));
 sky130_fd_sc_hd__o21a_1 _13083_ (.A1(_00220_),
    .A2(net169),
    .B1(net419),
    .X(_00088_));
 sky130_fd_sc_hd__o221a_1 _13084_ (.A1(\div_shifter[22] ),
    .A2(net253),
    .B1(net186),
    .B2(net403),
    .C1(net281),
    .X(_06164_));
 sky130_fd_sc_hd__o21a_1 _13085_ (.A1(net95),
    .A2(net169),
    .B1(net404),
    .X(_00089_));
 sky130_fd_sc_hd__o221a_1 _13086_ (.A1(\div_shifter[23] ),
    .A2(net253),
    .B1(net186),
    .B2(net367),
    .C1(net281),
    .X(_06165_));
 sky130_fd_sc_hd__o21a_1 _13087_ (.A1(_00259_),
    .A2(net169),
    .B1(net368),
    .X(_00090_));
 sky130_fd_sc_hd__o221a_1 _13088_ (.A1(net367),
    .A2(net253),
    .B1(net186),
    .B2(net308),
    .C1(net280),
    .X(_06166_));
 sky130_fd_sc_hd__o21a_1 _13089_ (.A1(net91),
    .A2(net169),
    .B1(net371),
    .X(_00091_));
 sky130_fd_sc_hd__o221a_1 _13090_ (.A1(net308),
    .A2(net254),
    .B1(net186),
    .B2(\div_shifter[26] ),
    .C1(net280),
    .X(_06167_));
 sky130_fd_sc_hd__o21a_1 _13091_ (.A1(_00246_),
    .A2(net168),
    .B1(net309),
    .X(_00092_));
 sky130_fd_sc_hd__o221a_1 _13092_ (.A1(\div_shifter[26] ),
    .A2(net254),
    .B1(net186),
    .B2(net411),
    .C1(net280),
    .X(_06168_));
 sky130_fd_sc_hd__o21a_1 _13093_ (.A1(net92),
    .A2(net168),
    .B1(net412),
    .X(_00093_));
 sky130_fd_sc_hd__o221a_1 _13094_ (.A1(net411),
    .A2(net253),
    .B1(net185),
    .B2(net351),
    .C1(net280),
    .X(_06170_));
 sky130_fd_sc_hd__o21a_1 _13095_ (.A1(_00451_),
    .A2(net168),
    .B1(net439),
    .X(_00094_));
 sky130_fd_sc_hd__a221o_1 _13096_ (.A1(net352),
    .A2(net255),
    .B1(net187),
    .B2(net301),
    .C1(rst),
    .X(_06171_));
 sky130_fd_sc_hd__a21oi_1 _13097_ (.A1(net71),
    .A2(net172),
    .B1(_06171_),
    .Y(_00095_));
 sky130_fd_sc_hd__a221o_1 _13098_ (.A1(net301),
    .A2(net255),
    .B1(net187),
    .B2(_04400_),
    .C1(rst),
    .X(_06172_));
 sky130_fd_sc_hd__a21oi_1 _13099_ (.A1(_01964_),
    .A2(net172),
    .B1(net302),
    .Y(_00096_));
 sky130_fd_sc_hd__a21oi_1 _13100_ (.A1(_04400_),
    .A2(net255),
    .B1(rst),
    .Y(_06173_));
 sky130_fd_sc_hd__o221a_1 _13101_ (.A1(net311),
    .A2(net185),
    .B1(net22),
    .B2(net168),
    .C1(_06173_),
    .X(_00097_));
 sky130_fd_sc_hd__nand3_1 _13102_ (.A(net311),
    .B(net306),
    .C(net2),
    .Y(_06174_));
 sky130_fd_sc_hd__a21o_1 _13103_ (.A1(net306),
    .A2(net2),
    .B1(net311),
    .X(_06175_));
 sky130_fd_sc_hd__a32o_1 _13104_ (.A1(net256),
    .A2(net598),
    .A3(_06175_),
    .B1(net187),
    .B2(net540),
    .X(_06177_));
 sky130_fd_sc_hd__and2_1 _13105_ (.A(net279),
    .B(net599),
    .X(_00098_));
 sky130_fd_sc_hd__xor2_1 _13106_ (.A(_06028_),
    .B(_06029_),
    .X(_06178_));
 sky130_fd_sc_hd__mux2_1 _13107_ (.A0(\div_shifter[32] ),
    .A1(_06178_),
    .S(net2),
    .X(_06179_));
 sky130_fd_sc_hd__a22o_1 _13108_ (.A1(net530),
    .A2(net187),
    .B1(_06179_),
    .B2(net255),
    .X(_06180_));
 sky130_fd_sc_hd__and2_1 _13109_ (.A(net279),
    .B(net531),
    .X(_00099_));
 sky130_fd_sc_hd__nand2_1 _13110_ (.A(_06026_),
    .B(_06032_),
    .Y(_06181_));
 sky130_fd_sc_hd__xnor2_1 _13111_ (.A(_06030_),
    .B(_06181_),
    .Y(_06182_));
 sky130_fd_sc_hd__mux2_1 _13112_ (.A0(net530),
    .A1(_06182_),
    .S(net2),
    .X(_06183_));
 sky130_fd_sc_hd__a22o_1 _13113_ (.A1(net590),
    .A2(net187),
    .B1(_06183_),
    .B2(net255),
    .X(_06184_));
 sky130_fd_sc_hd__and2_1 _13114_ (.A(net279),
    .B(_06184_),
    .X(_00100_));
 sky130_fd_sc_hd__nand2_1 _13115_ (.A(_06025_),
    .B(_06034_),
    .Y(_06186_));
 sky130_fd_sc_hd__xnor2_1 _13116_ (.A(_06033_),
    .B(_06186_),
    .Y(_06187_));
 sky130_fd_sc_hd__mux2_1 _13117_ (.A0(\div_shifter[34] ),
    .A1(_06187_),
    .S(net2),
    .X(_06188_));
 sky130_fd_sc_hd__a22o_1 _13118_ (.A1(net551),
    .A2(net187),
    .B1(_06188_),
    .B2(net255),
    .X(_06189_));
 sky130_fd_sc_hd__and2_1 _13119_ (.A(net279),
    .B(net552),
    .X(_00101_));
 sky130_fd_sc_hd__xnor2_1 _13120_ (.A(_06024_),
    .B(_06035_),
    .Y(_06190_));
 sky130_fd_sc_hd__mux2_1 _13121_ (.A0(net551),
    .A1(_06190_),
    .S(net2),
    .X(_06191_));
 sky130_fd_sc_hd__a22o_1 _13122_ (.A1(net585),
    .A2(net187),
    .B1(_06191_),
    .B2(net255),
    .X(_06192_));
 sky130_fd_sc_hd__and2_1 _13123_ (.A(net279),
    .B(net586),
    .X(_00102_));
 sky130_fd_sc_hd__xnor2_1 _13124_ (.A(_06021_),
    .B(_06036_),
    .Y(_06194_));
 sky130_fd_sc_hd__mux2_1 _13125_ (.A0(\div_shifter[36] ),
    .A1(_06194_),
    .S(net2),
    .X(_06195_));
 sky130_fd_sc_hd__a22o_1 _13126_ (.A1(net543),
    .A2(net187),
    .B1(_06195_),
    .B2(net255),
    .X(_06196_));
 sky130_fd_sc_hd__and2_1 _13127_ (.A(net279),
    .B(net544),
    .X(_00103_));
 sky130_fd_sc_hd__nand2_1 _13128_ (.A(_06017_),
    .B(_06038_),
    .Y(_06197_));
 sky130_fd_sc_hd__xnor2_1 _13129_ (.A(_06037_),
    .B(_06197_),
    .Y(_06198_));
 sky130_fd_sc_hd__mux2_1 _13130_ (.A0(net543),
    .A1(_06198_),
    .S(net2),
    .X(_06199_));
 sky130_fd_sc_hd__a22o_1 _13131_ (.A1(net555),
    .A2(net187),
    .B1(_06199_),
    .B2(net255),
    .X(_06200_));
 sky130_fd_sc_hd__and2_1 _13132_ (.A(net279),
    .B(net556),
    .X(_00104_));
 sky130_fd_sc_hd__nand2_1 _13133_ (.A(_06016_),
    .B(_06040_),
    .Y(_06201_));
 sky130_fd_sc_hd__xnor2_1 _13134_ (.A(_06039_),
    .B(_06201_),
    .Y(_06203_));
 sky130_fd_sc_hd__mux2_1 _13135_ (.A0(net555),
    .A1(_06203_),
    .S(net2),
    .X(_06204_));
 sky130_fd_sc_hd__a22o_1 _13136_ (.A1(net576),
    .A2(net187),
    .B1(_06204_),
    .B2(net255),
    .X(_06205_));
 sky130_fd_sc_hd__and2_1 _13137_ (.A(net279),
    .B(_06205_),
    .X(_00105_));
 sky130_fd_sc_hd__nand2_1 _13138_ (.A(_06015_),
    .B(_06043_),
    .Y(_06206_));
 sky130_fd_sc_hd__xnor2_1 _13139_ (.A(_06041_),
    .B(_06206_),
    .Y(_06207_));
 sky130_fd_sc_hd__mux2_1 _13140_ (.A0(\div_shifter[39] ),
    .A1(_06207_),
    .S(net2),
    .X(_06208_));
 sky130_fd_sc_hd__a22o_1 _13141_ (.A1(net547),
    .A2(net187),
    .B1(_06208_),
    .B2(net256),
    .X(_06209_));
 sky130_fd_sc_hd__and2_1 _13142_ (.A(net283),
    .B(net548),
    .X(_00106_));
 sky130_fd_sc_hd__nand2_1 _13143_ (.A(_06014_),
    .B(_06045_),
    .Y(_06210_));
 sky130_fd_sc_hd__xnor2_1 _13144_ (.A(_06044_),
    .B(_06210_),
    .Y(_06212_));
 sky130_fd_sc_hd__mux2_1 _13145_ (.A0(net547),
    .A1(_06212_),
    .S(net2),
    .X(_06213_));
 sky130_fd_sc_hd__a22o_1 _13146_ (.A1(net589),
    .A2(_06465_),
    .B1(_06213_),
    .B2(net256),
    .X(_06214_));
 sky130_fd_sc_hd__and2_1 _13147_ (.A(net279),
    .B(_06214_),
    .X(_00107_));
 sky130_fd_sc_hd__nand2_1 _13148_ (.A(_06013_),
    .B(_06047_),
    .Y(_06215_));
 sky130_fd_sc_hd__xnor2_1 _13149_ (.A(_06046_),
    .B(_06215_),
    .Y(_06216_));
 sky130_fd_sc_hd__mux2_1 _13150_ (.A0(\div_shifter[41] ),
    .A1(_06216_),
    .S(net1),
    .X(_06217_));
 sky130_fd_sc_hd__a22o_1 _13151_ (.A1(net574),
    .A2(net191),
    .B1(_06217_),
    .B2(net260),
    .X(_06218_));
 sky130_fd_sc_hd__and2_1 _13152_ (.A(net282),
    .B(net575),
    .X(_00108_));
 sky130_fd_sc_hd__nand2_1 _13153_ (.A(_06012_),
    .B(_06049_),
    .Y(_06219_));
 sky130_fd_sc_hd__xnor2_1 _13154_ (.A(_06048_),
    .B(_06219_),
    .Y(_06221_));
 sky130_fd_sc_hd__mux2_1 _13155_ (.A0(net574),
    .A1(_06221_),
    .S(_06096_),
    .X(_06222_));
 sky130_fd_sc_hd__a22o_1 _13156_ (.A1(net583),
    .A2(net191),
    .B1(_06222_),
    .B2(net260),
    .X(_06223_));
 sky130_fd_sc_hd__and2_1 _13157_ (.A(net282),
    .B(net584),
    .X(_00109_));
 sky130_fd_sc_hd__nand2_1 _13158_ (.A(_06011_),
    .B(_06051_),
    .Y(_06224_));
 sky130_fd_sc_hd__xnor2_1 _13159_ (.A(_06050_),
    .B(_06224_),
    .Y(_06225_));
 sky130_fd_sc_hd__mux2_1 _13160_ (.A0(\div_shifter[43] ),
    .A1(_06225_),
    .S(net2),
    .X(_06226_));
 sky130_fd_sc_hd__a22o_1 _13161_ (.A1(net580),
    .A2(net189),
    .B1(_06226_),
    .B2(net258),
    .X(_06227_));
 sky130_fd_sc_hd__and2_1 _13162_ (.A(net277),
    .B(net581),
    .X(_00110_));
 sky130_fd_sc_hd__nand2_1 _13163_ (.A(_06010_),
    .B(_06054_),
    .Y(_06228_));
 sky130_fd_sc_hd__xnor2_1 _13164_ (.A(_06052_),
    .B(_06228_),
    .Y(_06230_));
 sky130_fd_sc_hd__mux2_1 _13165_ (.A0(\div_shifter[44] ),
    .A1(_06230_),
    .S(net2),
    .X(_06231_));
 sky130_fd_sc_hd__a22o_1 _13166_ (.A1(net565),
    .A2(net189),
    .B1(_06231_),
    .B2(net258),
    .X(_06232_));
 sky130_fd_sc_hd__and2_1 _13167_ (.A(net276),
    .B(net566),
    .X(_00111_));
 sky130_fd_sc_hd__nand2_1 _13168_ (.A(_06008_),
    .B(_06056_),
    .Y(_06233_));
 sky130_fd_sc_hd__xnor2_1 _13169_ (.A(_06055_),
    .B(_06233_),
    .Y(_06234_));
 sky130_fd_sc_hd__mux2_1 _13170_ (.A0(net565),
    .A1(_06234_),
    .S(net1),
    .X(_06235_));
 sky130_fd_sc_hd__a22o_1 _13171_ (.A1(net567),
    .A2(net190),
    .B1(_06235_),
    .B2(net258),
    .X(_06236_));
 sky130_fd_sc_hd__and2_1 _13172_ (.A(net276),
    .B(net568),
    .X(_00112_));
 sky130_fd_sc_hd__nand2_1 _13173_ (.A(_06007_),
    .B(_06058_),
    .Y(_06237_));
 sky130_fd_sc_hd__xnor2_1 _13174_ (.A(_06057_),
    .B(_06237_),
    .Y(_06239_));
 sky130_fd_sc_hd__mux2_1 _13175_ (.A0(net567),
    .A1(_06239_),
    .S(net1),
    .X(_06240_));
 sky130_fd_sc_hd__a22o_1 _13176_ (.A1(net570),
    .A2(net190),
    .B1(_06240_),
    .B2(net259),
    .X(_06241_));
 sky130_fd_sc_hd__and2_1 _13177_ (.A(net274),
    .B(_06241_),
    .X(_00113_));
 sky130_fd_sc_hd__nand2_1 _13178_ (.A(_06006_),
    .B(_06060_),
    .Y(_06242_));
 sky130_fd_sc_hd__xnor2_1 _13179_ (.A(_06059_),
    .B(_06242_),
    .Y(_06243_));
 sky130_fd_sc_hd__mux2_1 _13180_ (.A0(net570),
    .A1(_06243_),
    .S(net1),
    .X(_06244_));
 sky130_fd_sc_hd__a22o_1 _13181_ (.A1(net587),
    .A2(net190),
    .B1(_06244_),
    .B2(net259),
    .X(_06245_));
 sky130_fd_sc_hd__and2_1 _13182_ (.A(net274),
    .B(_06245_),
    .X(_00114_));
 sky130_fd_sc_hd__nand2_1 _13183_ (.A(_06005_),
    .B(_06062_),
    .Y(_06246_));
 sky130_fd_sc_hd__xnor2_1 _13184_ (.A(_06061_),
    .B(_06246_),
    .Y(_06248_));
 sky130_fd_sc_hd__mux2_1 _13185_ (.A0(\div_shifter[48] ),
    .A1(_06248_),
    .S(net1),
    .X(_06249_));
 sky130_fd_sc_hd__a22o_1 _13186_ (.A1(net541),
    .A2(net190),
    .B1(_06249_),
    .B2(net259),
    .X(_06250_));
 sky130_fd_sc_hd__and2_1 _13187_ (.A(net274),
    .B(net542),
    .X(_00115_));
 sky130_fd_sc_hd__nand2b_1 _13188_ (.A_N(_06003_),
    .B(_06004_),
    .Y(_06251_));
 sky130_fd_sc_hd__xnor2_1 _13189_ (.A(_06063_),
    .B(_06251_),
    .Y(_06252_));
 sky130_fd_sc_hd__mux2_1 _13190_ (.A0(net541),
    .A1(_06252_),
    .S(net1),
    .X(_06253_));
 sky130_fd_sc_hd__a22o_1 _13191_ (.A1(net559),
    .A2(net190),
    .B1(_06253_),
    .B2(net259),
    .X(_06254_));
 sky130_fd_sc_hd__and2_1 _13192_ (.A(net274),
    .B(net560),
    .X(_00116_));
 sky130_fd_sc_hd__nand2_1 _13193_ (.A(_06002_),
    .B(_06066_),
    .Y(_06255_));
 sky130_fd_sc_hd__xnor2_1 _13194_ (.A(_06065_),
    .B(_06255_),
    .Y(_06257_));
 sky130_fd_sc_hd__mux2_1 _13195_ (.A0(\div_shifter[50] ),
    .A1(_06257_),
    .S(net1),
    .X(_06258_));
 sky130_fd_sc_hd__a22o_1 _13196_ (.A1(net557),
    .A2(net190),
    .B1(_06258_),
    .B2(net259),
    .X(_06259_));
 sky130_fd_sc_hd__and2_1 _13197_ (.A(net274),
    .B(net558),
    .X(_00117_));
 sky130_fd_sc_hd__xnor2_1 _13198_ (.A(_06067_),
    .B(_06069_),
    .Y(_06260_));
 sky130_fd_sc_hd__mux2_1 _13199_ (.A0(net557),
    .A1(_06260_),
    .S(net1),
    .X(_06261_));
 sky130_fd_sc_hd__a22o_1 _13200_ (.A1(net569),
    .A2(net190),
    .B1(_06261_),
    .B2(net259),
    .X(_06262_));
 sky130_fd_sc_hd__and2_1 _13201_ (.A(net274),
    .B(_06262_),
    .X(_00118_));
 sky130_fd_sc_hd__nand2_1 _13202_ (.A(_06000_),
    .B(_06071_),
    .Y(_06263_));
 sky130_fd_sc_hd__xnor2_1 _13203_ (.A(_06070_),
    .B(_06263_),
    .Y(_06264_));
 sky130_fd_sc_hd__mux2_1 _13204_ (.A0(\div_shifter[52] ),
    .A1(_06264_),
    .S(net1),
    .X(_06266_));
 sky130_fd_sc_hd__a22o_1 _13205_ (.A1(net563),
    .A2(net190),
    .B1(_06266_),
    .B2(net259),
    .X(_06267_));
 sky130_fd_sc_hd__and2_1 _13206_ (.A(net274),
    .B(net564),
    .X(_00119_));
 sky130_fd_sc_hd__xnor2_1 _13207_ (.A(_06072_),
    .B(_06074_),
    .Y(_06268_));
 sky130_fd_sc_hd__mux2_1 _13208_ (.A0(\div_shifter[53] ),
    .A1(_06268_),
    .S(net1),
    .X(_06269_));
 sky130_fd_sc_hd__a22o_1 _13209_ (.A1(net561),
    .A2(net189),
    .B1(_06269_),
    .B2(net259),
    .X(_06270_));
 sky130_fd_sc_hd__and2_1 _13210_ (.A(net274),
    .B(net562),
    .X(_00120_));
 sky130_fd_sc_hd__nand2_1 _13211_ (.A(_05997_),
    .B(_06077_),
    .Y(_06271_));
 sky130_fd_sc_hd__xnor2_1 _13212_ (.A(_06076_),
    .B(_06271_),
    .Y(_06272_));
 sky130_fd_sc_hd__mux2_1 _13213_ (.A0(\div_shifter[54] ),
    .A1(_06272_),
    .S(net1),
    .X(_06273_));
 sky130_fd_sc_hd__a22o_1 _13214_ (.A1(net549),
    .A2(net190),
    .B1(_06273_),
    .B2(net259),
    .X(_06275_));
 sky130_fd_sc_hd__and2_1 _13215_ (.A(net276),
    .B(net550),
    .X(_00121_));
 sky130_fd_sc_hd__xnor2_1 _13216_ (.A(_06078_),
    .B(_06080_),
    .Y(_06276_));
 sky130_fd_sc_hd__mux2_1 _13217_ (.A0(net549),
    .A1(_06276_),
    .S(net1),
    .X(_06277_));
 sky130_fd_sc_hd__a22o_1 _13218_ (.A1(net573),
    .A2(net190),
    .B1(_06277_),
    .B2(net259),
    .X(_06278_));
 sky130_fd_sc_hd__and2_1 _13219_ (.A(net276),
    .B(_06278_),
    .X(_00122_));
 sky130_fd_sc_hd__nand2_1 _13220_ (.A(_05995_),
    .B(_06082_),
    .Y(_06279_));
 sky130_fd_sc_hd__xnor2_1 _13221_ (.A(_06081_),
    .B(_06279_),
    .Y(_06280_));
 sky130_fd_sc_hd__mux2_1 _13222_ (.A0(\div_shifter[56] ),
    .A1(_06280_),
    .S(net2),
    .X(_06281_));
 sky130_fd_sc_hd__a22o_1 _13223_ (.A1(net571),
    .A2(net190),
    .B1(_06281_),
    .B2(net259),
    .X(_06282_));
 sky130_fd_sc_hd__and2_1 _13224_ (.A(net276),
    .B(net572),
    .X(_00123_));
 sky130_fd_sc_hd__xnor2_1 _13225_ (.A(_05994_),
    .B(_06083_),
    .Y(_06284_));
 sky130_fd_sc_hd__mux2_1 _13226_ (.A0(net571),
    .A1(_06284_),
    .S(net1),
    .X(_06285_));
 sky130_fd_sc_hd__a22o_1 _13227_ (.A1(net579),
    .A2(net191),
    .B1(_06285_),
    .B2(net260),
    .X(_06286_));
 sky130_fd_sc_hd__and2_1 _13228_ (.A(net276),
    .B(_06286_),
    .X(_00124_));
 sky130_fd_sc_hd__nand2_1 _13229_ (.A(_05991_),
    .B(_06085_),
    .Y(_06287_));
 sky130_fd_sc_hd__xnor2_1 _13230_ (.A(_06084_),
    .B(_06287_),
    .Y(_06288_));
 sky130_fd_sc_hd__mux2_1 _13231_ (.A0(\div_shifter[58] ),
    .A1(_06288_),
    .S(net1),
    .X(_06289_));
 sky130_fd_sc_hd__a22o_1 _13232_ (.A1(net577),
    .A2(net191),
    .B1(_06289_),
    .B2(net260),
    .X(_06290_));
 sky130_fd_sc_hd__and2_1 _13233_ (.A(net282),
    .B(net578),
    .X(_00125_));
 sky130_fd_sc_hd__xnor2_1 _13234_ (.A(_06087_),
    .B(_06089_),
    .Y(_06292_));
 sky130_fd_sc_hd__mux2_1 _13235_ (.A0(net577),
    .A1(_06292_),
    .S(_06096_),
    .X(_06293_));
 sky130_fd_sc_hd__a22o_1 _13236_ (.A1(net582),
    .A2(net191),
    .B1(_06293_),
    .B2(net260),
    .X(_06294_));
 sky130_fd_sc_hd__and2_1 _13237_ (.A(net282),
    .B(_06294_),
    .X(_00126_));
 sky130_fd_sc_hd__nand2_1 _13238_ (.A(_05989_),
    .B(_06091_),
    .Y(_06295_));
 sky130_fd_sc_hd__xnor2_1 _13239_ (.A(_06090_),
    .B(_06295_),
    .Y(_06296_));
 sky130_fd_sc_hd__mux2_1 _13240_ (.A0(\div_shifter[60] ),
    .A1(_06296_),
    .S(net1),
    .X(_06297_));
 sky130_fd_sc_hd__a22o_1 _13241_ (.A1(net553),
    .A2(net191),
    .B1(_06297_),
    .B2(net260),
    .X(_06298_));
 sky130_fd_sc_hd__and2_1 _13242_ (.A(net282),
    .B(net554),
    .X(_00127_));
 sky130_fd_sc_hd__xnor2_1 _13243_ (.A(_05988_),
    .B(_06092_),
    .Y(_06299_));
 sky130_fd_sc_hd__mux2_1 _13244_ (.A0(\div_shifter[61] ),
    .A1(_06299_),
    .S(net1),
    .X(_06301_));
 sky130_fd_sc_hd__a22o_1 _13245_ (.A1(net545),
    .A2(net191),
    .B1(_06301_),
    .B2(net260),
    .X(_06302_));
 sky130_fd_sc_hd__and2_1 _13246_ (.A(net282),
    .B(net546),
    .X(_00128_));
 sky130_fd_sc_hd__nand2b_1 _13247_ (.A_N(_06094_),
    .B(_06095_),
    .Y(_06303_));
 sky130_fd_sc_hd__a32o_1 _13248_ (.A1(net592),
    .A2(net260),
    .A3(_06303_),
    .B1(net191),
    .B2(net470),
    .X(_06304_));
 sky130_fd_sc_hd__and2_1 _13249_ (.A(net276),
    .B(net471),
    .X(_00129_));
 sky130_fd_sc_hd__nand2_1 _13250_ (.A(net435),
    .B(net186),
    .Y(_06305_));
 sky130_fd_sc_hd__o211a_1 _13251_ (.A1(net435),
    .A2(net256),
    .B1(net280),
    .C1(net436),
    .X(_00130_));
 sky130_fd_sc_hd__a22o_1 _13252_ (.A1(net462),
    .A2(net187),
    .B1(_05937_),
    .B2(net255),
    .X(_06306_));
 sky130_fd_sc_hd__o211a_1 _13253_ (.A1(net462),
    .A2(net435),
    .B1(net280),
    .C1(_06306_),
    .X(_00131_));
 sky130_fd_sc_hd__a22o_1 _13254_ (.A1(net422),
    .A2(net187),
    .B1(_05938_),
    .B2(net255),
    .X(_06308_));
 sky130_fd_sc_hd__a21o_1 _13255_ (.A1(net462),
    .A2(net435),
    .B1(net422),
    .X(_06309_));
 sky130_fd_sc_hd__and3_1 _13256_ (.A(net281),
    .B(_06308_),
    .C(net601),
    .X(_00132_));
 sky130_fd_sc_hd__a22o_1 _13257_ (.A1(net361),
    .A2(net188),
    .B1(_05940_),
    .B2(net256),
    .X(_06310_));
 sky130_fd_sc_hd__a31o_1 _13258_ (.A1(net422),
    .A2(\div_counter[1] ),
    .A3(\div_counter[0] ),
    .B1(net361),
    .X(_06311_));
 sky130_fd_sc_hd__and3_1 _13259_ (.A(net281),
    .B(_06310_),
    .C(net423),
    .X(_00133_));
 sky130_fd_sc_hd__a22o_1 _13260_ (.A1(net298),
    .A2(_06465_),
    .B1(_05941_),
    .B2(net256),
    .X(_06312_));
 sky130_fd_sc_hd__o211a_1 _13261_ (.A1(net298),
    .A2(net594),
    .B1(_06312_),
    .C1(net281),
    .X(_00134_));
 sky130_fd_sc_hd__o21a_1 _13262_ (.A1(net455),
    .A2(_05942_),
    .B1(net283),
    .X(_00135_));
 sky130_fd_sc_hd__dfxtp_1 _13263_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net364),
    .Q(busy_l));
 sky130_fd_sc_hd__dfxtp_1 _13264_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00001_),
    .Q(divi1_sign));
 sky130_fd_sc_hd__dfxtp_1 _13265_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net307),
    .Q(\divi2_l[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13266_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00003_),
    .Q(\divi2_l[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13267_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00004_),
    .Q(\divi2_l[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13268_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00005_),
    .Q(\divi2_l[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13269_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00006_),
    .Q(\divi2_l[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13270_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00007_),
    .Q(\divi2_l[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13271_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00008_),
    .Q(\divi2_l[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13272_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00009_),
    .Q(\divi2_l[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13273_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00010_),
    .Q(\divi2_l[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13274_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00011_),
    .Q(\divi2_l[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13275_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00012_),
    .Q(\divi2_l[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13276_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00013_),
    .Q(\divi2_l[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13277_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00014_),
    .Q(\divi2_l[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13278_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00015_),
    .Q(\divi2_l[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13279_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00016_),
    .Q(\divi2_l[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13280_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00017_),
    .Q(\divi2_l[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13281_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00018_),
    .Q(\divi2_l[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13282_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00019_),
    .Q(\divi2_l[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13283_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00020_),
    .Q(\divi2_l[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13284_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00021_),
    .Q(\divi2_l[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13285_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00022_),
    .Q(\divi2_l[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13286_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00023_),
    .Q(\divi2_l[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13287_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00024_),
    .Q(\divi2_l[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13288_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00025_),
    .Q(\divi2_l[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13289_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00026_),
    .Q(\divi2_l[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13290_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00027_),
    .Q(\divi2_l[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13291_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00028_),
    .Q(\divi2_l[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13292_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00029_),
    .Q(\divi2_l[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13293_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00030_),
    .Q(\divi2_l[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13294_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00031_),
    .Q(\divi2_l[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13295_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00032_),
    .Q(\divi2_l[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13296_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00033_),
    .Q(\divi2_l[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13297_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00034_),
    .Q(\div_res[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13298_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00035_),
    .Q(\div_res[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13299_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00036_),
    .Q(\div_res[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13300_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net518),
    .Q(\div_res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13301_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00038_),
    .Q(\div_res[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13302_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00039_),
    .Q(\div_res[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13303_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00040_),
    .Q(\div_res[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13304_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00041_),
    .Q(\div_res[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13305_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00042_),
    .Q(\div_res[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13306_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net505),
    .Q(\div_res[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13307_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00044_),
    .Q(\div_res[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13308_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net482),
    .Q(\div_res[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13309_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00046_),
    .Q(\div_res[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13310_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net466),
    .Q(\div_res[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13311_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net490),
    .Q(\div_res[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13312_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net479),
    .Q(\div_res[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13313_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00050_),
    .Q(\div_res[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13314_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net474),
    .Q(\div_res[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13315_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00052_),
    .Q(\div_res[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13316_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00053_),
    .Q(\div_res[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13317_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net469),
    .Q(\div_res[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13318_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net485),
    .Q(\div_res[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13319_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00056_),
    .Q(\div_res[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13320_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net498),
    .Q(\div_res[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13321_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00058_),
    .Q(\div_res[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13322_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net459),
    .Q(\div_res[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13323_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net526),
    .Q(\div_res[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13324_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net521),
    .Q(\div_res[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13325_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00062_),
    .Q(\div_res[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13326_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00063_),
    .Q(\div_res[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13327_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net529),
    .Q(\div_res[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13328_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(net434),
    .Q(\div_res[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13329_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00066_),
    .Q(\div_shifter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13330_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00067_),
    .Q(\div_shifter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13331_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00068_),
    .Q(\div_shifter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13332_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net336),
    .Q(\div_shifter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13333_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00070_),
    .Q(\div_shifter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13334_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net297),
    .Q(\div_shifter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13335_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00072_),
    .Q(\div_shifter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13336_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net444),
    .Q(\div_shifter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13337_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00074_),
    .Q(\div_shifter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13338_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00075_),
    .Q(\div_shifter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13339_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00076_),
    .Q(\div_shifter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13340_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00077_),
    .Q(\div_shifter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13341_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net379),
    .Q(\div_shifter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13342_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net427),
    .Q(\div_shifter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13343_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00080_),
    .Q(\div_shifter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13344_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00081_),
    .Q(\div_shifter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13345_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net376),
    .Q(\div_shifter[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13346_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net397),
    .Q(\div_shifter[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13347_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00084_),
    .Q(\div_shifter[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13348_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net410),
    .Q(\div_shifter[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13349_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net400),
    .Q(\div_shifter[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13350_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net386),
    .Q(\div_shifter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13351_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00088_),
    .Q(\div_shifter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13352_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net405),
    .Q(\div_shifter[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13353_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net369),
    .Q(\div_shifter[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13354_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00091_),
    .Q(\div_shifter[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13355_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net310),
    .Q(\div_shifter[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13356_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net413),
    .Q(\div_shifter[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13357_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00094_),
    .Q(\div_shifter[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13358_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00095_),
    .Q(\div_shifter[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13359_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net303),
    .Q(\div_shifter[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13360_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net312),
    .Q(\div_shifter[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13361_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00098_),
    .Q(\div_shifter[32] ));
 sky130_fd_sc_hd__dfxtp_1 _13362_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00099_),
    .Q(\div_shifter[33] ));
 sky130_fd_sc_hd__dfxtp_1 _13363_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00100_),
    .Q(\div_shifter[34] ));
 sky130_fd_sc_hd__dfxtp_1 _13364_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00101_),
    .Q(\div_shifter[35] ));
 sky130_fd_sc_hd__dfxtp_1 _13365_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00102_),
    .Q(\div_shifter[36] ));
 sky130_fd_sc_hd__dfxtp_1 _13366_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00103_),
    .Q(\div_shifter[37] ));
 sky130_fd_sc_hd__dfxtp_1 _13367_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00104_),
    .Q(\div_shifter[38] ));
 sky130_fd_sc_hd__dfxtp_1 _13368_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00105_),
    .Q(\div_shifter[39] ));
 sky130_fd_sc_hd__dfxtp_1 _13369_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00106_),
    .Q(\div_shifter[40] ));
 sky130_fd_sc_hd__dfxtp_1 _13370_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00107_),
    .Q(\div_shifter[41] ));
 sky130_fd_sc_hd__dfxtp_1 _13371_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00108_),
    .Q(\div_shifter[42] ));
 sky130_fd_sc_hd__dfxtp_1 _13372_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00109_),
    .Q(\div_shifter[43] ));
 sky130_fd_sc_hd__dfxtp_1 _13373_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00110_),
    .Q(\div_shifter[44] ));
 sky130_fd_sc_hd__dfxtp_1 _13374_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00111_),
    .Q(\div_shifter[45] ));
 sky130_fd_sc_hd__dfxtp_1 _13375_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00112_),
    .Q(\div_shifter[46] ));
 sky130_fd_sc_hd__dfxtp_1 _13376_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00113_),
    .Q(\div_shifter[47] ));
 sky130_fd_sc_hd__dfxtp_1 _13377_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00114_),
    .Q(\div_shifter[48] ));
 sky130_fd_sc_hd__dfxtp_1 _13378_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00115_),
    .Q(\div_shifter[49] ));
 sky130_fd_sc_hd__dfxtp_1 _13379_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00116_),
    .Q(\div_shifter[50] ));
 sky130_fd_sc_hd__dfxtp_1 _13380_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00117_),
    .Q(\div_shifter[51] ));
 sky130_fd_sc_hd__dfxtp_1 _13381_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00118_),
    .Q(\div_shifter[52] ));
 sky130_fd_sc_hd__dfxtp_1 _13382_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00119_),
    .Q(\div_shifter[53] ));
 sky130_fd_sc_hd__dfxtp_1 _13383_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00120_),
    .Q(\div_shifter[54] ));
 sky130_fd_sc_hd__dfxtp_1 _13384_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00121_),
    .Q(\div_shifter[55] ));
 sky130_fd_sc_hd__dfxtp_1 _13385_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00122_),
    .Q(\div_shifter[56] ));
 sky130_fd_sc_hd__dfxtp_1 _13386_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00123_),
    .Q(\div_shifter[57] ));
 sky130_fd_sc_hd__dfxtp_1 _13387_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00124_),
    .Q(\div_shifter[58] ));
 sky130_fd_sc_hd__dfxtp_1 _13388_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00125_),
    .Q(\div_shifter[59] ));
 sky130_fd_sc_hd__dfxtp_1 _13389_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00126_),
    .Q(\div_shifter[60] ));
 sky130_fd_sc_hd__dfxtp_1 _13390_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00127_),
    .Q(\div_shifter[61] ));
 sky130_fd_sc_hd__dfxtp_1 _13391_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00128_),
    .Q(\div_shifter[62] ));
 sky130_fd_sc_hd__dfxtp_1 _13392_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00129_),
    .Q(\div_shifter[63] ));
 sky130_fd_sc_hd__dfxtp_1 _13393_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net437),
    .Q(\div_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13394_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net463),
    .Q(\div_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13395_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net602),
    .Q(\div_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13396_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net424),
    .Q(\div_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13397_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net299),
    .Q(\div_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13398_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net456),
    .Q(div_complete));
 sky130_fd_sc_hd__buf_12 _13399_ (.A(instruction[11]),
    .X(loadstore_dest[0]));
 sky130_fd_sc_hd__buf_12 _13400_ (.A(instruction[12]),
    .X(loadstore_dest[1]));
 sky130_fd_sc_hd__buf_12 _13401_ (.A(instruction[13]),
    .X(loadstore_dest[2]));
 sky130_fd_sc_hd__buf_12 _13402_ (.A(instruction[14]),
    .X(loadstore_dest[3]));
 sky130_fd_sc_hd__buf_12 _13403_ (.A(instruction[15]),
    .X(loadstore_dest[4]));
 sky130_fd_sc_hd__buf_12 _13404_ (.A(instruction[16]),
    .X(loadstore_dest[5]));
 sky130_fd_sc_hd__buf_12 _13405_ (.A(instruction[5]),
    .X(loadstore_size[0]));
 sky130_fd_sc_hd__buf_12 _13406_ (.A(instruction[6]),
    .X(loadstore_size[1]));
 sky130_fd_sc_hd__buf_12 _13407_ (.A(instruction[8]),
    .X(pred_idx[0]));
 sky130_fd_sc_hd__buf_12 _13408_ (.A(instruction[9]),
    .X(pred_idx[1]));
 sky130_fd_sc_hd__buf_12 _13409_ (.A(instruction[10]),
    .X(pred_idx[2]));
 sky130_fd_sc_hd__buf_12 _13410_ (.A(instruction[4]),
    .X(sign_extend));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__buf_6 fanout1 (.A(net2),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_8 fanout10 (.A(net11),
    .X(net10));
 sky130_fd_sc_hd__buf_8 fanout100 (.A(_00180_),
    .X(net100));
 sky130_fd_sc_hd__buf_4 fanout101 (.A(_00180_),
    .X(net101));
 sky130_fd_sc_hd__buf_6 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__buf_8 fanout105 (.A(_00391_),
    .X(net105));
 sky130_fd_sc_hd__buf_6 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_8 fanout107 (.A(_00390_),
    .X(net107));
 sky130_fd_sc_hd__buf_8 fanout108 (.A(_00375_),
    .X(net108));
 sky130_fd_sc_hd__buf_6 fanout109 (.A(_00329_),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_8 fanout11 (.A(_01968_),
    .X(net11));
 sky130_fd_sc_hd__buf_4 fanout110 (.A(_00329_),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_8 fanout111 (.A(_00325_),
    .X(net111));
 sky130_fd_sc_hd__buf_4 fanout112 (.A(_00325_),
    .X(net112));
 sky130_fd_sc_hd__buf_6 fanout114 (.A(_00313_),
    .X(net114));
 sky130_fd_sc_hd__buf_8 fanout115 (.A(_00309_),
    .X(net115));
 sky130_fd_sc_hd__buf_8 fanout117 (.A(_00290_),
    .X(net117));
 sky130_fd_sc_hd__buf_8 fanout119 (.A(_00286_),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_8 fanout12 (.A(net13),
    .X(net12));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(_00286_),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_16 fanout121 (.A(net123),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_16 fanout122 (.A(net123),
    .X(net122));
 sky130_fd_sc_hd__buf_12 fanout123 (.A(_00279_),
    .X(net123));
 sky130_fd_sc_hd__buf_12 fanout124 (.A(_00276_),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_16 fanout125 (.A(_00275_),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_8 fanout126 (.A(_00275_),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_8 fanout127 (.A(_00227_),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_4 fanout128 (.A(_00227_),
    .X(net128));
 sky130_fd_sc_hd__buf_6 fanout129 (.A(_00212_),
    .X(net129));
 sky130_fd_sc_hd__buf_4 fanout13 (.A(_01952_),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_4 fanout130 (.A(_00212_),
    .X(net130));
 sky130_fd_sc_hd__buf_6 fanout131 (.A(_00190_),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_8 fanout132 (.A(_00190_),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_8 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_8 fanout134 (.A(_00184_),
    .X(net134));
 sky130_fd_sc_hd__buf_12 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__buf_12 fanout136 (.A(_00341_),
    .X(net136));
 sky130_fd_sc_hd__buf_12 fanout137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__buf_12 fanout138 (.A(_00338_),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_8 fanout14 (.A(_00699_),
    .X(net14));
 sky130_fd_sc_hd__buf_6 fanout140 (.A(_00264_),
    .X(net140));
 sky130_fd_sc_hd__buf_6 fanout141 (.A(_00257_),
    .X(net141));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(_00257_),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_8 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__buf_4 fanout144 (.A(_00241_),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_8 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__buf_8 fanout146 (.A(_00166_),
    .X(net146));
 sky130_fd_sc_hd__buf_6 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__buf_8 fanout148 (.A(_00160_),
    .X(net148));
 sky130_fd_sc_hd__buf_8 fanout149 (.A(_06564_),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_8 fanout15 (.A(net16),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout150 (.A(_06564_),
    .X(net150));
 sky130_fd_sc_hd__buf_6 fanout151 (.A(_06558_),
    .X(net151));
 sky130_fd_sc_hd__buf_4 fanout152 (.A(_06558_),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_8 fanout153 (.A(_06542_),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_8 fanout154 (.A(_06542_),
    .X(net154));
 sky130_fd_sc_hd__buf_6 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__buf_8 fanout156 (.A(_06538_),
    .X(net156));
 sky130_fd_sc_hd__buf_4 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__buf_4 fanout159 (.A(net160),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_8 fanout16 (.A(_00688_),
    .X(net16));
 sky130_fd_sc_hd__buf_4 fanout160 (.A(_06490_),
    .X(net160));
 sky130_fd_sc_hd__buf_4 fanout161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 fanout162 (.A(net167),
    .X(net162));
 sky130_fd_sc_hd__buf_4 fanout163 (.A(net167),
    .X(net163));
 sky130_fd_sc_hd__buf_4 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__buf_4 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__buf_4 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__buf_4 fanout167 (.A(_06489_),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_8 fanout168 (.A(_05945_),
    .X(net168));
 sky130_fd_sc_hd__buf_2 fanout169 (.A(_05945_),
    .X(net169));
 sky130_fd_sc_hd__buf_6 fanout17 (.A(_00409_),
    .X(net17));
 sky130_fd_sc_hd__buf_4 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__buf_2 fanout171 (.A(_05945_),
    .X(net171));
 sky130_fd_sc_hd__buf_4 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_4 fanout173 (.A(_05944_),
    .X(net173));
 sky130_fd_sc_hd__buf_4 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__buf_2 fanout175 (.A(_05944_),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_8 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_8 fanout177 (.A(_02245_),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_8 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_8 fanout179 (.A(_02244_),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_8 fanout18 (.A(_02079_),
    .X(net18));
 sky130_fd_sc_hd__buf_12 fanout180 (.A(net182),
    .X(net180));
 sky130_fd_sc_hd__buf_12 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__buf_8 fanout182 (.A(_00178_),
    .X(net182));
 sky130_fd_sc_hd__buf_6 fanout183 (.A(_06496_),
    .X(net183));
 sky130_fd_sc_hd__buf_8 fanout184 (.A(_06495_),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(_06466_),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_4 fanout186 (.A(_06466_),
    .X(net186));
 sky130_fd_sc_hd__buf_4 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_8 fanout188 (.A(_06465_),
    .X(net188));
 sky130_fd_sc_hd__buf_4 fanout189 (.A(net191),
    .X(net189));
 sky130_fd_sc_hd__buf_6 fanout19 (.A(net21),
    .X(net19));
 sky130_fd_sc_hd__buf_4 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__buf_4 fanout191 (.A(_06465_),
    .X(net191));
 sky130_fd_sc_hd__buf_4 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__buf_4 fanout193 (.A(_02331_),
    .X(net193));
 sky130_fd_sc_hd__buf_4 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__buf_4 fanout195 (.A(_02329_),
    .X(net195));
 sky130_fd_sc_hd__buf_4 fanout196 (.A(_02326_),
    .X(net196));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(_02320_),
    .X(net197));
 sky130_fd_sc_hd__buf_4 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 fanout199 (.A(_02316_),
    .X(net199));
 sky130_fd_sc_hd__buf_6 fanout2 (.A(_06096_),
    .X(net2));
 sky130_fd_sc_hd__buf_4 fanout20 (.A(net21),
    .X(net20));
 sky130_fd_sc_hd__buf_4 fanout200 (.A(_02241_),
    .X(net200));
 sky130_fd_sc_hd__buf_12 fanout201 (.A(net203),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_16 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__buf_6 fanout203 (.A(_00155_),
    .X(net203));
 sky130_fd_sc_hd__buf_12 fanout204 (.A(_06534_),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_16 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__buf_6 fanout206 (.A(_06534_),
    .X(net206));
 sky130_fd_sc_hd__buf_12 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__buf_12 fanout208 (.A(_06531_),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_8 fanout209 (.A(_06488_),
    .X(net209));
 sky130_fd_sc_hd__buf_12 fanout21 (.A(_02079_),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_8 fanout210 (.A(_06475_),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_8 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_4 fanout212 (.A(net213),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(net214),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_8 fanout214 (.A(_06365_),
    .X(net214));
 sky130_fd_sc_hd__buf_6 fanout215 (.A(net216),
    .X(net215));
 sky130_fd_sc_hd__buf_8 fanout216 (.A(_06364_),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_8 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_8 fanout218 (.A(_06360_),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(net220),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_16 fanout22 (.A(_02078_),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(_06353_),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(net223),
    .X(net222));
 sky130_fd_sc_hd__buf_2 fanout223 (.A(_06347_),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_8 fanout224 (.A(_06346_),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_8 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_4 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_4 fanout228 (.A(_06340_),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_8 fanout229 (.A(_06331_),
    .X(net229));
 sky130_fd_sc_hd__buf_6 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__buf_4 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 fanout231 (.A(_04893_),
    .X(net231));
 sky130_fd_sc_hd__buf_4 fanout232 (.A(net234),
    .X(net232));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net234),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 fanout234 (.A(_02514_),
    .X(net234));
 sky130_fd_sc_hd__buf_4 fanout235 (.A(_02514_),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_8 fanout236 (.A(_02318_),
    .X(net236));
 sky130_fd_sc_hd__buf_6 fanout237 (.A(_06520_),
    .X(net237));
 sky130_fd_sc_hd__buf_12 fanout238 (.A(_06494_),
    .X(net238));
 sky130_fd_sc_hd__buf_8 fanout239 (.A(_06494_),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_8 fanout24 (.A(_00453_),
    .X(net24));
 sky130_fd_sc_hd__buf_4 fanout241 (.A(_06487_),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_8 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_4 fanout243 (.A(net244),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_4 fanout244 (.A(net247),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_8 fanout245 (.A(net246),
    .X(net245));
 sky130_fd_sc_hd__buf_6 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__buf_6 fanout247 (.A(_06458_),
    .X(net247));
 sky130_fd_sc_hd__buf_12 fanout248 (.A(_06457_),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_8 fanout249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__buf_6 fanout25 (.A(_00327_),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_8 fanout250 (.A(_06330_),
    .X(net250));
 sky130_fd_sc_hd__buf_8 fanout251 (.A(net252),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_8 fanout252 (.A(_04871_),
    .X(net252));
 sky130_fd_sc_hd__buf_4 fanout253 (.A(_04465_),
    .X(net253));
 sky130_fd_sc_hd__buf_4 fanout254 (.A(_04465_),
    .X(net254));
 sky130_fd_sc_hd__buf_4 fanout255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_4 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_8 fanout257 (.A(net486),
    .X(net257));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(net260),
    .X(net258));
 sky130_fd_sc_hd__buf_4 fanout259 (.A(net260),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_8 fanout26 (.A(_00327_),
    .X(net26));
 sky130_fd_sc_hd__buf_4 fanout260 (.A(net486),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_8 fanout261 (.A(net262),
    .X(net261));
 sky130_fd_sc_hd__buf_4 fanout262 (.A(_06491_),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_8 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_8 fanout264 (.A(_04795_),
    .X(net264));
 sky130_fd_sc_hd__buf_12 fanout265 (.A(_04795_),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_8 fanout266 (.A(_04795_),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_8 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_8 fanout268 (.A(net269),
    .X(net268));
 sky130_fd_sc_hd__buf_4 fanout269 (.A(_04784_),
    .X(net269));
 sky130_fd_sc_hd__buf_6 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_8 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_4 fanout271 (.A(_04773_),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_8 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__buf_4 fanout273 (.A(_04585_),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__buf_2 fanout275 (.A(net277),
    .X(net275));
 sky130_fd_sc_hd__buf_4 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__buf_2 fanout277 (.A(net278),
    .X(net277));
 sky130_fd_sc_hd__buf_4 fanout278 (.A(_04553_),
    .X(net278));
 sky130_fd_sc_hd__buf_4 fanout279 (.A(net283),
    .X(net279));
 sky130_fd_sc_hd__buf_8 fanout28 (.A(_00323_),
    .X(net28));
 sky130_fd_sc_hd__buf_4 fanout280 (.A(net281),
    .X(net280));
 sky130_fd_sc_hd__buf_4 fanout281 (.A(net283),
    .X(net281));
 sky130_fd_sc_hd__buf_4 fanout282 (.A(net283),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 fanout283 (.A(_04553_),
    .X(net283));
 sky130_fd_sc_hd__buf_6 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__buf_4 fanout285 (.A(net286),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_8 fanout286 (.A(_04542_),
    .X(net286));
 sky130_fd_sc_hd__buf_6 fanout287 (.A(_04509_),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_8 fanout288 (.A(_04509_),
    .X(net288));
 sky130_fd_sc_hd__buf_12 fanout289 (.A(reg1_val[1]),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_8 fanout29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__buf_6 fanout290 (.A(reg1_val[15]),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_8 fanout291 (.A(reg1_val[14]),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_8 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__buf_4 fanout293 (.A(reg1_val[0]),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_8 fanout294 (.A(net295),
    .X(net294));
 sky130_fd_sc_hd__buf_8 fanout295 (.A(instruction[7]),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_8 fanout30 (.A(_00310_),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_8 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_8 fanout32 (.A(_00305_),
    .X(net32));
 sky130_fd_sc_hd__buf_8 fanout33 (.A(_00293_),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 fanout34 (.A(_00293_),
    .X(net34));
 sky130_fd_sc_hd__buf_8 fanout35 (.A(_00284_),
    .X(net35));
 sky130_fd_sc_hd__buf_4 fanout36 (.A(_00284_),
    .X(net36));
 sky130_fd_sc_hd__buf_6 fanout37 (.A(_00266_),
    .X(net37));
 sky130_fd_sc_hd__buf_4 fanout38 (.A(_00266_),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_8 fanout39 (.A(_00262_),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_8 fanout40 (.A(_00262_),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_8 fanout41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__buf_6 fanout42 (.A(_00251_),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_8 fanout43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__buf_6 fanout44 (.A(_00249_),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_8 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_6 fanout46 (.A(_00229_),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_8 fanout47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_8 fanout48 (.A(_00223_),
    .X(net48));
 sky130_fd_sc_hd__buf_12 fanout49 (.A(net50),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_8 fanout5 (.A(net6),
    .X(net5));
 sky130_fd_sc_hd__buf_12 fanout50 (.A(_00217_),
    .X(net50));
 sky130_fd_sc_hd__buf_8 fanout51 (.A(_00171_),
    .X(net51));
 sky130_fd_sc_hd__buf_4 fanout52 (.A(_00171_),
    .X(net52));
 sky130_fd_sc_hd__buf_6 fanout53 (.A(_00164_),
    .X(net53));
 sky130_fd_sc_hd__buf_4 fanout54 (.A(_00164_),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_8 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_8 fanout56 (.A(_00142_),
    .X(net56));
 sky130_fd_sc_hd__buf_8 fanout57 (.A(_06562_),
    .X(net57));
 sky130_fd_sc_hd__buf_4 fanout58 (.A(_06562_),
    .X(net58));
 sky130_fd_sc_hd__buf_8 fanout59 (.A(_06560_),
    .X(net59));
 sky130_fd_sc_hd__buf_4 fanout6 (.A(_02081_),
    .X(net6));
 sky130_fd_sc_hd__buf_4 fanout60 (.A(_06560_),
    .X(net60));
 sky130_fd_sc_hd__buf_6 fanout61 (.A(_06546_),
    .X(net61));
 sky130_fd_sc_hd__buf_4 fanout62 (.A(_06546_),
    .X(net62));
 sky130_fd_sc_hd__buf_6 fanout63 (.A(_06541_),
    .X(net63));
 sky130_fd_sc_hd__buf_4 fanout64 (.A(_06541_),
    .X(net64));
 sky130_fd_sc_hd__buf_6 fanout65 (.A(_06524_),
    .X(net65));
 sky130_fd_sc_hd__buf_4 fanout66 (.A(_06524_),
    .X(net66));
 sky130_fd_sc_hd__buf_6 fanout67 (.A(net68),
    .X(net67));
 sky130_fd_sc_hd__buf_8 fanout68 (.A(_06518_),
    .X(net68));
 sky130_fd_sc_hd__buf_8 fanout69 (.A(net71),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_8 fanout7 (.A(net8),
    .X(net7));
 sky130_fd_sc_hd__buf_4 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_6 fanout71 (.A(_00679_),
    .X(net71));
 sky130_fd_sc_hd__buf_8 fanout72 (.A(net73),
    .X(net72));
 sky130_fd_sc_hd__buf_6 fanout73 (.A(_00365_),
    .X(net73));
 sky130_fd_sc_hd__buf_6 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__buf_8 fanout75 (.A(_00363_),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_8 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__buf_6 fanout77 (.A(_00362_),
    .X(net77));
 sky130_fd_sc_hd__buf_6 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__buf_8 fanout79 (.A(_00360_),
    .X(net79));
 sky130_fd_sc_hd__buf_6 fanout8 (.A(_02067_),
    .X(net8));
 sky130_fd_sc_hd__buf_6 fanout80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_8 fanout81 (.A(_00353_),
    .X(net81));
 sky130_fd_sc_hd__buf_8 fanout82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__buf_8 fanout83 (.A(_00350_),
    .X(net83));
 sky130_fd_sc_hd__buf_6 fanout84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__buf_6 fanout85 (.A(_00349_),
    .X(net85));
 sky130_fd_sc_hd__buf_8 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_8 fanout87 (.A(_00347_),
    .X(net87));
 sky130_fd_sc_hd__buf_12 fanout88 (.A(_00301_),
    .X(net88));
 sky130_fd_sc_hd__buf_12 fanout89 (.A(_00301_),
    .X(net89));
 sky130_fd_sc_hd__buf_8 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__buf_8 fanout91 (.A(_00245_),
    .X(net91));
 sky130_fd_sc_hd__buf_8 fanout92 (.A(net94),
    .X(net92));
 sky130_fd_sc_hd__buf_8 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_16 fanout94 (.A(_00238_),
    .X(net94));
 sky130_fd_sc_hd__buf_8 fanout95 (.A(_00208_),
    .X(net95));
 sky130_fd_sc_hd__buf_4 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_16 fanout97 (.A(_00208_),
    .X(net97));
 sky130_fd_sc_hd__buf_6 fanout98 (.A(_00188_),
    .X(net98));
 sky130_fd_sc_hd__buf_4 fanout99 (.A(_00188_),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\div_shifter[5] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_05946_),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\div_shifter[17] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_06156_),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_00083_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\div_shifter[20] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_06160_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_00086_),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\divi2_l[13] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_05963_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\div_shifter[23] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_06164_),
    .X(net404));
 sky130_fd_sc_hd__buf_1 hold11 (.A(\divi2_l[0] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(_00089_),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\divi2_l[4] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_05952_),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\div_shifter[19] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_06159_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_00085_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(net438),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_06168_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_00093_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\div_shifter[0] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_00002_),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_06136_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\divi2_l[18] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(_05969_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\div_shifter[22] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(_06162_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\div_shifter[1] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(_06137_),
    .X(net421));
 sky130_fd_sc_hd__buf_1 hold127 (.A(net495),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(_06311_),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_00133_),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net370),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\div_shifter[13] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(_06152_),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_00079_),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\div_shifter[18] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_06158_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(net447),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(_06154_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\div_res[31] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_06135_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_00065_),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_06167_),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 hold140 (.A(net600),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_06305_),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_00130_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\div_shifter[27] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(_06170_),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\div_shifter[9] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_06148_),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\div_shifter[7] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(_06144_),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_00073_),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_00092_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net453),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_06147_),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\div_shifter[14] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_06153_),
    .X(net448));
 sky130_fd_sc_hd__buf_1 hold154 (.A(\divi2_l[1] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(_05948_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\div_shifter[6] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(_06143_),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\div_shifter[8] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(_06146_),
    .X(net454));
 sky130_fd_sc_hd__buf_1 hold16 (.A(net597),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(div_complete),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(_00135_),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(net501),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_06128_),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(_00059_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\div_shifter[2] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(_06138_),
    .X(net461));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold167 (.A(\div_counter[1] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(_00131_),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net493),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_00097_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_06113_),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(_00047_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\div_res[19] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_06122_),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(_00054_),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\div_shifter[63] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_06304_),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\div_res[17] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_06118_),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(_00051_),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\divi2_l[6] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\div_res[18] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_06120_),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\div_res[15] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_06116_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(_00049_),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\div_res[11] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(_06111_),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_00045_),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\div_res[21] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(_06123_),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_05954_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_00055_),
    .X(net485));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold191 (.A(busy_l),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_06119_),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\div_res[14] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(_06114_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_00048_),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\div_res[5] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(_06104_),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\div_res[12] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_06112_),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_00071_),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\divi2_l[15] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\div_counter[2] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\div_res[23] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_06125_),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(_00057_),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\div_res[16] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(_06117_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\div_res[24] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(_06126_),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\div_res[9] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_06108_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_05965_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(_00043_),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\div_res[6] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_06105_),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\div_res[10] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_06110_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\div_res[7] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(_06106_),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\div_res[8] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(_06107_),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\div_res[22] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\divi2_l[10] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(_06124_),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\div_res[3] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(_06101_),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_00037_),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\div_res[27] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_06130_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_00061_),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\div_res[28] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(_06131_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\div_res[26] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(_05959_),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_06129_),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(_00060_),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\div_res[30] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(_06134_),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_00064_),
    .X(net529));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold235 (.A(\div_shifter[33] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_06180_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\div_res[2] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_06100_),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\div_res[4] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\divi2_l[23] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_06102_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\div_res[29] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_06132_),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\div_res[1] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_06099_),
    .X(net539));
 sky130_fd_sc_hd__buf_1 hold245 (.A(\div_shifter[32] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\div_shifter[49] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(_06250_),
    .X(net542));
 sky130_fd_sc_hd__buf_1 hold248 (.A(\div_shifter[37] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(_06196_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_05975_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\div_shifter[62] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(_06302_),
    .X(net546));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold252 (.A(\div_shifter[40] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(_06209_),
    .X(net548));
 sky130_fd_sc_hd__buf_1 hold254 (.A(\div_shifter[55] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(_06275_),
    .X(net550));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold256 (.A(\div_shifter[35] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(_06189_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\div_shifter[61] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(_06298_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\divi2_l[30] ),
    .X(net321));
 sky130_fd_sc_hd__buf_1 hold260 (.A(\div_shifter[38] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_06200_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\div_shifter[51] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(_06259_),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\div_shifter[50] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(_06254_),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\div_shifter[54] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(_06270_),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\div_shifter[53] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_06267_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_05983_),
    .X(net322));
 sky130_fd_sc_hd__buf_1 hold270 (.A(\div_shifter[45] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(_06232_),
    .X(net566));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold272 (.A(\div_shifter[46] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(_06236_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\div_shifter[52] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\div_shifter[47] ),
    .X(net570));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold276 (.A(\div_shifter[57] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(_06282_),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\div_shifter[56] ),
    .X(net573));
 sky130_fd_sc_hd__buf_1 hold279 (.A(\div_shifter[42] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\divi2_l[29] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_06218_),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\div_shifter[39] ),
    .X(net576));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold282 (.A(\div_shifter[59] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(_06290_),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\div_shifter[58] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\div_shifter[44] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_06227_),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\div_shifter[60] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\div_shifter[43] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(_06223_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(_05982_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\div_shifter[36] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(_06192_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\div_shifter[48] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\div_res[0] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\div_shifter[41] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\div_shifter[34] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\div_shifter[30] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\div_shifter[62] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\div_counter[1] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(_05939_),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\div_counter[4] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\divi2_l[8] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\div_res[4] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\div_res[1] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\div_shifter[31] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(_06174_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(_06177_),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\div_counter[0] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(_06309_),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(_00132_),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_05957_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\divi2_l[9] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_05958_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\divi2_l[21] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(_05972_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\divi2_l[16] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(_05966_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\div_shifter[3] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_04444_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_00134_),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_06140_),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_00069_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\div_shifter[4] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_04433_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\divi2_l[26] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_05978_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\divi2_l[7] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(_05955_),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\divi2_l[31] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(_05984_),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\div_shifter[29] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\divi2_l[14] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_05964_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\divi2_l[20] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(_05971_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\divi2_l[5] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(_05953_),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\div_shifter[28] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_04422_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\divi2_l[28] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(_05981_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_04411_),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\divi2_l[27] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_05979_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\divi2_l[22] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_05973_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\divi2_l[25] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_05977_),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\div_counter[3] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_05939_),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(_05941_),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_00000_),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(_06172_),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\divi2_l[2] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_05949_),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\div_shifter[24] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_06165_),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_00090_),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\div_shifter[25] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(_06166_),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\divi2_l[24] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_05976_),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\div_shifter[15] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_00096_),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_06155_),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_00082_),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\div_shifter[11] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(_06150_),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_00078_),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\divi2_l[11] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_05960_),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\divi2_l[17] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(_05967_),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\div_shifter[21] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(divi1_sign),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_06161_),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_00087_),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\divi2_l[3] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_05951_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\divi2_l[12] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_05961_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\divi2_l[19] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(_05970_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\div_shifter[10] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_06149_),
    .X(net394));
 sky130_fd_sc_hd__buf_4 max_cap102 (.A(_00179_),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 max_cap103 (.A(_05773_),
    .X(net103));
 sky130_fd_sc_hd__buf_4 max_cap113 (.A(_00314_),
    .X(net113));
 sky130_fd_sc_hd__clkbuf_8 max_cap116 (.A(_00291_),
    .X(net116));
 sky130_fd_sc_hd__buf_4 max_cap118 (.A(_00287_),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 max_cap139 (.A(_00312_),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_8 max_cap225 (.A(_06341_),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_8 max_cap240 (.A(_06493_),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 max_cap3 (.A(_03745_),
    .X(net3));
 sky130_fd_sc_hd__buf_1 max_cap4 (.A(_03091_),
    .X(net4));
 sky130_fd_sc_hd__buf_4 max_cap9 (.A(_02066_),
    .X(net9));
endmodule

