magic
tech sky130B
magscale 1 2
timestamp 1717695836
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 934 2128 59510 57928
<< metal2 >>
rect 938 59200 994 60000
rect 2594 59200 2650 60000
rect 4250 59200 4306 60000
rect 5906 59200 5962 60000
rect 7562 59200 7618 60000
rect 9218 59200 9274 60000
rect 10874 59200 10930 60000
rect 12530 59200 12586 60000
rect 14186 59200 14242 60000
rect 15842 59200 15898 60000
rect 17498 59200 17554 60000
rect 19154 59200 19210 60000
rect 20810 59200 20866 60000
rect 22466 59200 22522 60000
rect 24122 59200 24178 60000
rect 25778 59200 25834 60000
rect 27434 59200 27490 60000
rect 29090 59200 29146 60000
rect 30746 59200 30802 60000
rect 32402 59200 32458 60000
rect 34058 59200 34114 60000
rect 35714 59200 35770 60000
rect 37370 59200 37426 60000
rect 39026 59200 39082 60000
rect 40682 59200 40738 60000
rect 42338 59200 42394 60000
rect 43994 59200 44050 60000
rect 45650 59200 45706 60000
rect 47306 59200 47362 60000
rect 48962 59200 49018 60000
rect 50618 59200 50674 60000
rect 52274 59200 52330 60000
rect 53930 59200 53986 60000
rect 55586 59200 55642 60000
rect 57242 59200 57298 60000
rect 58898 59200 58954 60000
rect 938 0 994 800
rect 2594 0 2650 800
rect 4250 0 4306 800
rect 5906 0 5962 800
rect 7562 0 7618 800
rect 9218 0 9274 800
rect 10874 0 10930 800
rect 12530 0 12586 800
rect 14186 0 14242 800
rect 15842 0 15898 800
rect 17498 0 17554 800
rect 19154 0 19210 800
rect 20810 0 20866 800
rect 22466 0 22522 800
rect 24122 0 24178 800
rect 25778 0 25834 800
rect 27434 0 27490 800
rect 29090 0 29146 800
rect 30746 0 30802 800
rect 32402 0 32458 800
rect 34058 0 34114 800
rect 35714 0 35770 800
rect 37370 0 37426 800
rect 39026 0 39082 800
rect 40682 0 40738 800
rect 42338 0 42394 800
rect 43994 0 44050 800
rect 45650 0 45706 800
rect 47306 0 47362 800
rect 48962 0 49018 800
rect 50618 0 50674 800
rect 52274 0 52330 800
rect 53930 0 53986 800
rect 55586 0 55642 800
rect 57242 0 57298 800
rect 58898 0 58954 800
<< obsm2 >>
rect 1050 59144 2538 59200
rect 2706 59144 4194 59200
rect 4362 59144 5850 59200
rect 6018 59144 7506 59200
rect 7674 59144 9162 59200
rect 9330 59144 10818 59200
rect 10986 59144 12474 59200
rect 12642 59144 14130 59200
rect 14298 59144 15786 59200
rect 15954 59144 17442 59200
rect 17610 59144 19098 59200
rect 19266 59144 20754 59200
rect 20922 59144 22410 59200
rect 22578 59144 24066 59200
rect 24234 59144 25722 59200
rect 25890 59144 27378 59200
rect 27546 59144 29034 59200
rect 29202 59144 30690 59200
rect 30858 59144 32346 59200
rect 32514 59144 34002 59200
rect 34170 59144 35658 59200
rect 35826 59144 37314 59200
rect 37482 59144 38970 59200
rect 39138 59144 40626 59200
rect 40794 59144 42282 59200
rect 42450 59144 43938 59200
rect 44106 59144 45594 59200
rect 45762 59144 47250 59200
rect 47418 59144 48906 59200
rect 49074 59144 50562 59200
rect 50730 59144 52218 59200
rect 52386 59144 53874 59200
rect 54042 59144 55530 59200
rect 55698 59144 57186 59200
rect 57354 59144 58842 59200
rect 59010 59144 59504 59200
rect 938 856 59504 59144
rect 1050 734 2538 856
rect 2706 734 4194 856
rect 4362 734 5850 856
rect 6018 734 7506 856
rect 7674 734 9162 856
rect 9330 734 10818 856
rect 10986 734 12474 856
rect 12642 734 14130 856
rect 14298 734 15786 856
rect 15954 734 17442 856
rect 17610 734 19098 856
rect 19266 734 20754 856
rect 20922 734 22410 856
rect 22578 734 24066 856
rect 24234 734 25722 856
rect 25890 734 27378 856
rect 27546 734 29034 856
rect 29202 734 30690 856
rect 30858 734 32346 856
rect 32514 734 34002 856
rect 34170 734 35658 856
rect 35826 734 37314 856
rect 37482 734 38970 856
rect 39138 734 40626 856
rect 40794 734 42282 856
rect 42450 734 43938 856
rect 44106 734 45594 856
rect 45762 734 47250 856
rect 47418 734 48906 856
rect 49074 734 50562 856
rect 50730 734 52218 856
rect 52386 734 53874 856
rect 54042 734 55530 856
rect 55698 734 57186 856
rect 57354 734 58842 856
rect 59010 734 59504 856
<< metal3 >>
rect 59200 58488 60000 58608
rect 59200 56856 60000 56976
rect 0 55224 800 55344
rect 59200 55224 60000 55344
rect 59200 53592 60000 53712
rect 59200 51960 60000 52080
rect 59200 50328 60000 50448
rect 59200 48696 60000 48816
rect 59200 47064 60000 47184
rect 0 46792 800 46912
rect 59200 45432 60000 45552
rect 59200 43800 60000 43920
rect 59200 42168 60000 42288
rect 59200 40536 60000 40656
rect 59200 38904 60000 39024
rect 0 38360 800 38480
rect 59200 37272 60000 37392
rect 59200 35640 60000 35760
rect 59200 34008 60000 34128
rect 59200 32376 60000 32496
rect 59200 30744 60000 30864
rect 0 29928 800 30048
rect 59200 29112 60000 29232
rect 59200 27480 60000 27600
rect 59200 25848 60000 25968
rect 59200 24216 60000 24336
rect 59200 22584 60000 22704
rect 0 21496 800 21616
rect 59200 20952 60000 21072
rect 59200 19320 60000 19440
rect 59200 17688 60000 17808
rect 59200 16056 60000 16176
rect 59200 14424 60000 14544
rect 0 13064 800 13184
rect 59200 12792 60000 12912
rect 59200 11160 60000 11280
rect 59200 9528 60000 9648
rect 59200 7896 60000 8016
rect 59200 6264 60000 6384
rect 0 4632 800 4752
rect 59200 4632 60000 4752
rect 59200 3000 60000 3120
rect 59200 1368 60000 1488
<< obsm3 >>
rect 798 58408 59120 58581
rect 798 57056 59327 58408
rect 798 56776 59120 57056
rect 798 55424 59327 56776
rect 880 55144 59120 55424
rect 798 53792 59327 55144
rect 798 53512 59120 53792
rect 798 52160 59327 53512
rect 798 51880 59120 52160
rect 798 50528 59327 51880
rect 798 50248 59120 50528
rect 798 48896 59327 50248
rect 798 48616 59120 48896
rect 798 47264 59327 48616
rect 798 46992 59120 47264
rect 880 46984 59120 46992
rect 880 46712 59327 46984
rect 798 45632 59327 46712
rect 798 45352 59120 45632
rect 798 44000 59327 45352
rect 798 43720 59120 44000
rect 798 42368 59327 43720
rect 798 42088 59120 42368
rect 798 40736 59327 42088
rect 798 40456 59120 40736
rect 798 39104 59327 40456
rect 798 38824 59120 39104
rect 798 38560 59327 38824
rect 880 38280 59327 38560
rect 798 37472 59327 38280
rect 798 37192 59120 37472
rect 798 35840 59327 37192
rect 798 35560 59120 35840
rect 798 34208 59327 35560
rect 798 33928 59120 34208
rect 798 32576 59327 33928
rect 798 32296 59120 32576
rect 798 30944 59327 32296
rect 798 30664 59120 30944
rect 798 30128 59327 30664
rect 880 29848 59327 30128
rect 798 29312 59327 29848
rect 798 29032 59120 29312
rect 798 27680 59327 29032
rect 798 27400 59120 27680
rect 798 26048 59327 27400
rect 798 25768 59120 26048
rect 798 24416 59327 25768
rect 798 24136 59120 24416
rect 798 22784 59327 24136
rect 798 22504 59120 22784
rect 798 21696 59327 22504
rect 880 21416 59327 21696
rect 798 21152 59327 21416
rect 798 20872 59120 21152
rect 798 19520 59327 20872
rect 798 19240 59120 19520
rect 798 17888 59327 19240
rect 798 17608 59120 17888
rect 798 16256 59327 17608
rect 798 15976 59120 16256
rect 798 14624 59327 15976
rect 798 14344 59120 14624
rect 798 13264 59327 14344
rect 880 12992 59327 13264
rect 880 12984 59120 12992
rect 798 12712 59120 12984
rect 798 11360 59327 12712
rect 798 11080 59120 11360
rect 798 9728 59327 11080
rect 798 9448 59120 9728
rect 798 8096 59327 9448
rect 798 7816 59120 8096
rect 798 6464 59327 7816
rect 798 6184 59120 6464
rect 798 4832 59327 6184
rect 880 4552 59120 4832
rect 798 3200 59327 4552
rect 798 2920 59120 3200
rect 798 1568 59327 2920
rect 798 1395 59120 1568
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< obsm4 >>
rect 8339 3843 19488 56677
rect 19968 3843 34848 56677
rect 35328 3843 50208 56677
rect 50688 3843 57901 56677
<< labels >>
rlabel metal3 s 0 21496 800 21616 6 custom_settings[0]
port 1 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 custom_settings[1]
port 2 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 custom_settings[2]
port 3 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 custom_settings[3]
port 4 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 custom_settings[4]
port 5 nsew signal input
rlabel metal2 s 938 59200 994 60000 6 io_in[0]
port 6 nsew signal input
rlabel metal2 s 17498 59200 17554 60000 6 io_in[10]
port 7 nsew signal input
rlabel metal2 s 19154 59200 19210 60000 6 io_in[11]
port 8 nsew signal input
rlabel metal2 s 20810 59200 20866 60000 6 io_in[12]
port 9 nsew signal input
rlabel metal2 s 22466 59200 22522 60000 6 io_in[13]
port 10 nsew signal input
rlabel metal2 s 24122 59200 24178 60000 6 io_in[14]
port 11 nsew signal input
rlabel metal2 s 25778 59200 25834 60000 6 io_in[15]
port 12 nsew signal input
rlabel metal2 s 27434 59200 27490 60000 6 io_in[16]
port 13 nsew signal input
rlabel metal2 s 29090 59200 29146 60000 6 io_in[17]
port 14 nsew signal input
rlabel metal2 s 30746 59200 30802 60000 6 io_in[18]
port 15 nsew signal input
rlabel metal2 s 32402 59200 32458 60000 6 io_in[19]
port 16 nsew signal input
rlabel metal2 s 2594 59200 2650 60000 6 io_in[1]
port 17 nsew signal input
rlabel metal2 s 34058 59200 34114 60000 6 io_in[20]
port 18 nsew signal input
rlabel metal2 s 35714 59200 35770 60000 6 io_in[21]
port 19 nsew signal input
rlabel metal2 s 37370 59200 37426 60000 6 io_in[22]
port 20 nsew signal input
rlabel metal2 s 39026 59200 39082 60000 6 io_in[23]
port 21 nsew signal input
rlabel metal2 s 40682 59200 40738 60000 6 io_in[24]
port 22 nsew signal input
rlabel metal2 s 42338 59200 42394 60000 6 io_in[25]
port 23 nsew signal input
rlabel metal2 s 43994 59200 44050 60000 6 io_in[26]
port 24 nsew signal input
rlabel metal2 s 45650 59200 45706 60000 6 io_in[27]
port 25 nsew signal input
rlabel metal2 s 47306 59200 47362 60000 6 io_in[28]
port 26 nsew signal input
rlabel metal2 s 48962 59200 49018 60000 6 io_in[29]
port 27 nsew signal input
rlabel metal2 s 4250 59200 4306 60000 6 io_in[2]
port 28 nsew signal input
rlabel metal2 s 50618 59200 50674 60000 6 io_in[30]
port 29 nsew signal input
rlabel metal2 s 52274 59200 52330 60000 6 io_in[31]
port 30 nsew signal input
rlabel metal2 s 53930 59200 53986 60000 6 io_in[32]
port 31 nsew signal input
rlabel metal2 s 55586 59200 55642 60000 6 io_in[33]
port 32 nsew signal input
rlabel metal2 s 57242 59200 57298 60000 6 io_in[34]
port 33 nsew signal input
rlabel metal2 s 58898 59200 58954 60000 6 io_in[35]
port 34 nsew signal input
rlabel metal2 s 5906 59200 5962 60000 6 io_in[3]
port 35 nsew signal input
rlabel metal2 s 7562 59200 7618 60000 6 io_in[4]
port 36 nsew signal input
rlabel metal2 s 9218 59200 9274 60000 6 io_in[5]
port 37 nsew signal input
rlabel metal2 s 10874 59200 10930 60000 6 io_in[6]
port 38 nsew signal input
rlabel metal2 s 12530 59200 12586 60000 6 io_in[7]
port 39 nsew signal input
rlabel metal2 s 14186 59200 14242 60000 6 io_in[8]
port 40 nsew signal input
rlabel metal2 s 15842 59200 15898 60000 6 io_in[9]
port 41 nsew signal input
rlabel metal2 s 938 0 994 800 6 io_oeb[0]
port 42 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 io_oeb[10]
port 43 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 io_oeb[11]
port 44 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 io_oeb[12]
port 45 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 io_oeb[13]
port 46 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 io_oeb[14]
port 47 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 io_oeb[15]
port 48 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 io_oeb[16]
port 49 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 io_oeb[17]
port 50 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 io_oeb[18]
port 51 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 io_oeb[19]
port 52 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 io_oeb[1]
port 53 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 io_oeb[20]
port 54 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 io_oeb[21]
port 55 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 io_oeb[22]
port 56 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 io_oeb[23]
port 57 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 io_oeb[24]
port 58 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 io_oeb[25]
port 59 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 io_oeb[26]
port 60 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 io_oeb[27]
port 61 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 io_oeb[28]
port 62 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 io_oeb[29]
port 63 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 io_oeb[2]
port 64 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 io_oeb[30]
port 65 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 io_oeb[31]
port 66 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 io_oeb[32]
port 67 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 io_oeb[33]
port 68 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 io_oeb[34]
port 69 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 io_oeb[35]
port 70 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 io_oeb[3]
port 71 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 io_oeb[4]
port 72 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 io_oeb[5]
port 73 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 io_oeb[6]
port 74 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 io_oeb[7]
port 75 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 io_oeb[8]
port 76 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 io_oeb[9]
port 77 nsew signal output
rlabel metal3 s 59200 1368 60000 1488 6 io_out[0]
port 78 nsew signal output
rlabel metal3 s 59200 17688 60000 17808 6 io_out[10]
port 79 nsew signal output
rlabel metal3 s 59200 19320 60000 19440 6 io_out[11]
port 80 nsew signal output
rlabel metal3 s 59200 20952 60000 21072 6 io_out[12]
port 81 nsew signal output
rlabel metal3 s 59200 22584 60000 22704 6 io_out[13]
port 82 nsew signal output
rlabel metal3 s 59200 24216 60000 24336 6 io_out[14]
port 83 nsew signal output
rlabel metal3 s 59200 25848 60000 25968 6 io_out[15]
port 84 nsew signal output
rlabel metal3 s 59200 27480 60000 27600 6 io_out[16]
port 85 nsew signal output
rlabel metal3 s 59200 29112 60000 29232 6 io_out[17]
port 86 nsew signal output
rlabel metal3 s 59200 30744 60000 30864 6 io_out[18]
port 87 nsew signal output
rlabel metal3 s 59200 32376 60000 32496 6 io_out[19]
port 88 nsew signal output
rlabel metal3 s 59200 3000 60000 3120 6 io_out[1]
port 89 nsew signal output
rlabel metal3 s 59200 34008 60000 34128 6 io_out[20]
port 90 nsew signal output
rlabel metal3 s 59200 35640 60000 35760 6 io_out[21]
port 91 nsew signal output
rlabel metal3 s 59200 37272 60000 37392 6 io_out[22]
port 92 nsew signal output
rlabel metal3 s 59200 38904 60000 39024 6 io_out[23]
port 93 nsew signal output
rlabel metal3 s 59200 40536 60000 40656 6 io_out[24]
port 94 nsew signal output
rlabel metal3 s 59200 42168 60000 42288 6 io_out[25]
port 95 nsew signal output
rlabel metal3 s 59200 43800 60000 43920 6 io_out[26]
port 96 nsew signal output
rlabel metal3 s 59200 45432 60000 45552 6 io_out[27]
port 97 nsew signal output
rlabel metal3 s 59200 47064 60000 47184 6 io_out[28]
port 98 nsew signal output
rlabel metal3 s 59200 48696 60000 48816 6 io_out[29]
port 99 nsew signal output
rlabel metal3 s 59200 4632 60000 4752 6 io_out[2]
port 100 nsew signal output
rlabel metal3 s 59200 50328 60000 50448 6 io_out[30]
port 101 nsew signal output
rlabel metal3 s 59200 51960 60000 52080 6 io_out[31]
port 102 nsew signal output
rlabel metal3 s 59200 53592 60000 53712 6 io_out[32]
port 103 nsew signal output
rlabel metal3 s 59200 55224 60000 55344 6 io_out[33]
port 104 nsew signal output
rlabel metal3 s 59200 56856 60000 56976 6 io_out[34]
port 105 nsew signal output
rlabel metal3 s 59200 58488 60000 58608 6 io_out[35]
port 106 nsew signal output
rlabel metal3 s 59200 6264 60000 6384 6 io_out[3]
port 107 nsew signal output
rlabel metal3 s 59200 7896 60000 8016 6 io_out[4]
port 108 nsew signal output
rlabel metal3 s 59200 9528 60000 9648 6 io_out[5]
port 109 nsew signal output
rlabel metal3 s 59200 11160 60000 11280 6 io_out[6]
port 110 nsew signal output
rlabel metal3 s 59200 12792 60000 12912 6 io_out[7]
port 111 nsew signal output
rlabel metal3 s 59200 14424 60000 14544 6 io_out[8]
port 112 nsew signal output
rlabel metal3 s 59200 16056 60000 16176 6 io_out[9]
port 113 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 rst_n
port 114 nsew signal input
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 115 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 116 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 116 nsew ground bidirectional
rlabel metal3 s 0 4632 800 4752 6 wb_clk_i
port 117 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16034142
string GDS_FILE /home/tholin/Desktop/ci2406-rej-pommedeterrible-tholin/openlane/Z80/runs/24_06_06_19_30/results/signoff/ci2406_z80.magic.gds
string GDS_START 1324990
<< end >>

