* NGSPICE file created from ci2406_z80.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_4 abstract view
.subckt sky130_fd_sc_hd__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_4 abstract view
.subckt sky130_fd_sc_hd__and2b_4 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_2 abstract view
.subckt sky130_fd_sc_hd__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

.subckt ci2406_z80 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15]
+ io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23]
+ io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31]
+ io_in[32] io_in[33] io_in[34] io_in[35] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[3]
+ io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10]
+ io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18]
+ io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25]
+ io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32]
+ io_out[33] io_out[34] io_out[35] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] rst_n vccd1 vssd1 wb_clk_i
XFILLER_0_94_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3676__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3155_ _3777_/B _4412_/A _3129_/X _3137_/A _3180_/B vssd1 vssd1 vccd1 vccd1 _3155_/X
+ sky130_fd_sc_hd__o32a_1
X_3086_ _3086_/A _3177_/A _3086_/C vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__or3_2
XFILLER_0_27_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5196__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3988_ _3988_/A _3988_/B _3988_/C vssd1 vssd1 vccd1 vccd1 _3988_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5727_ hold452/X _5714_/Y _5726_/X _5767_/A vssd1 vssd1 vccd1 vccd1 _5727_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5658_ _5658_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5659_/B sky130_fd_sc_hd__or2_1
XANTENNA__5705__S _5705_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4609_ _4609_/A _4609_/B vssd1 vssd1 vccd1 vccd1 _4611_/C sky130_fd_sc_hd__nand2_1
X_5589_ _5590_/A _5590_/B vssd1 vssd1 vccd1 vccd1 _5604_/A sky130_fd_sc_hd__nor2_1
Xhold340 _4989_/X vssd1 vssd1 vccd1 vccd1 _6091_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 _5497_/X vssd1 vssd1 vccd1 vccd1 _6187_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold351 _6081_/Q vssd1 vssd1 vccd1 vccd1 hold351/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold395 _5697_/X vssd1 vssd1 vccd1 vccd1 _6202_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 _6119_/Q vssd1 vssd1 vccd1 vccd1 _2980_/A sky130_fd_sc_hd__buf_1
Xhold373 _6117_/Q vssd1 vssd1 vccd1 vccd1 _2979_/A sky130_fd_sc_hd__buf_1
XANTENNA__6209__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4459__A1 _4391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4698__A1 _4990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3362__C _4043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5111__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5350__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4474__B _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4960_ _6240_/Q _5008_/B vssd1 vssd1 vccd1 vccd1 _4960_/X sky130_fd_sc_hd__and2_1
X_3911_ _3911_/A _4007_/S vssd1 vssd1 vccd1 vccd1 _3944_/A sky130_fd_sc_hd__or2_1
X_4891_ _6061_/Q _5595_/S _5607_/B1 _4890_/X vssd1 vssd1 vccd1 vccd1 _4891_/X sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_48_wb_clk_i_A _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3842_ _3239_/X _3646_/X _6117_/Q vssd1 vssd1 vccd1 vccd1 _3842_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_46_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3818__B _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3773_ _3773_/A _3773_/B vssd1 vssd1 vccd1 vccd1 _5387_/A sky130_fd_sc_hd__xnor2_2
X_5512_ _2984_/Y _5507_/Y _5508_/X vssd1 vssd1 vccd1 vccd1 _5514_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3537__C _4726_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5443_ _5317_/A _5343_/X _5352_/Y _6176_/Q vssd1 vssd1 vccd1 vccd1 _5443_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_14_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5374_ _5374_/A _5374_/B vssd1 vssd1 vccd1 vccd1 _5376_/A sky130_fd_sc_hd__xor2_1
X_4325_ _3930_/X hold147/X _4327_/S vssd1 vssd1 vccd1 vccd1 _4325_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout138 _6165_/Q vssd1 vssd1 vccd1 vccd1 _4714_/S sky130_fd_sc_hd__clkbuf_4
Xfanout127 _3426_/A vssd1 vssd1 vccd1 vccd1 _3777_/A sky130_fd_sc_hd__buf_4
Xfanout116 _3498_/A vssd1 vssd1 vccd1 vccd1 _3446_/A sky130_fd_sc_hd__buf_6
Xfanout105 _5424_/B vssd1 vssd1 vccd1 vccd1 _3457_/A sky130_fd_sc_hd__clkbuf_8
X_4256_ _4254_/X _4255_/X _4256_/S vssd1 vssd1 vccd1 vccd1 _4256_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout149 _4725_/B vssd1 vssd1 vccd1 vccd1 _3302_/A sky130_fd_sc_hd__buf_4
X_4187_ _4250_/A _4187_/B vssd1 vssd1 vccd1 vccd1 _4195_/B sky130_fd_sc_hd__xnor2_1
X_3207_ _4460_/A _4415_/A vssd1 vssd1 vccd1 vccd1 _3207_/X sky130_fd_sc_hd__or2_1
X_3138_ _3511_/C _4117_/C vssd1 vssd1 vccd1 vccd1 _3545_/A sky130_fd_sc_hd__and2_4
XFILLER_0_96_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3069_ _4726_/C _4614_/B _4728_/C vssd1 vssd1 vccd1 vccd1 _3177_/A sky130_fd_sc_hd__or3_1
XFILLER_0_9_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3744__A _5209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold170 _4275_/X vssd1 vssd1 vccd1 vccd1 _5937_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3463__B _4759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold181 _6166_/Q vssd1 vssd1 vccd1 vccd1 _3539_/B sky130_fd_sc_hd__buf_2
Xhold192 _6045_/Q vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4575__A _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3407__A2 _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4080__A2 _4750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4907__A2 _4761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4460__D _5341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4383__A3 _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5868__A0 _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4110_ hold94/X _3789_/X _4115_/S vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__mux2_1
X_5090_ _4451_/C _4392_/A _4385_/B _3439_/Y vssd1 vssd1 vccd1 vccd1 _5090_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5096__B2 _3488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4041_ _4070_/B _4446_/B _4412_/A vssd1 vssd1 vccd1 vccd1 _4750_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__4843__A1 _6158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4843__B2 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5992_ _6149_/CLK hold97/X vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_4_wb_clk_i_A _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4943_ _4990_/A _4943_/B vssd1 vssd1 vccd1 vccd1 _4943_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4874_ _5606_/S _4873_/X _4866_/X vssd1 vssd1 vccd1 vccd1 _4874_/X sky130_fd_sc_hd__a21o_1
X_3825_ _5033_/A _5387_/B _5403_/B _3648_/A vssd1 vssd1 vccd1 vccd1 _3825_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_6_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3756_ _4250_/A _3757_/B vssd1 vssd1 vccd1 vccd1 _3756_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5426_ _5426_/A _5426_/B vssd1 vssd1 vccd1 vccd1 _5426_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3687_ _3687_/A _3687_/B vssd1 vssd1 vccd1 vccd1 _3687_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3283__B _5093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5357_ _5484_/S vssd1 vssd1 vccd1 vccd1 _5794_/B sky130_fd_sc_hd__clkinv_4
X_4308_ _4242_/X hold254/X _4309_/S vssd1 vssd1 vccd1 vccd1 _5971_/D sky130_fd_sc_hd__mux2_1
X_5288_ _5245_/A hold482/X _5245_/Y _5287_/X vssd1 vssd1 vccd1 vccd1 _5288_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4509__S1 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4239_ _4239_/A _4239_/B vssd1 vssd1 vccd1 vccd1 _4239_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4395__A _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4598__A0 _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4334__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3193__B _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5173__S1 _5116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4684__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4590_ _4699_/A _4591_/B vssd1 vssd1 vccd1 vccd1 _4590_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3610_ _3616_/B _3607_/X _3609_/Y _3968_/A vssd1 vssd1 vccd1 vccd1 _3610_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3541_ _3545_/A _3540_/X _5502_/A vssd1 vssd1 vccd1 vccd1 _3541_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_51_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3472_ _4077_/A _3370_/B _3471_/Y _4460_/A vssd1 vssd1 vccd1 vccd1 _3472_/X sky130_fd_sc_hd__o2bb2a_1
X_5211_ _4260_/X _5185_/S _5210_/X vssd1 vssd1 vccd1 vccd1 _5211_/X sky130_fd_sc_hd__a21o_1
X_6191_ _6256_/CLK _6191_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6191_/Q sky130_fd_sc_hd__dfrtp_1
X_5142_ _6014_/Q _5200_/A2 _5200_/B1 _5947_/Q _4256_/S vssd1 vssd1 vccd1 vccd1 _5144_/B
+ sky130_fd_sc_hd__o221a_1
X_5073_ hold5/X _4233_/Y _5073_/S vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__mux2_1
XANTENNA__4816__A1 _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4024_ _5046_/A _3921_/A _3827_/B _6172_/Q _4023_/X vssd1 vssd1 vccd1 vccd1 _5394_/B
+ sky130_fd_sc_hd__a221o_2
XANTENNA__4943__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5975_ _6129_/CLK hold57/X fanout170/X vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__5241__A1 _5107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4926_ _4925_/X _6155_/Q _4926_/S vssd1 vssd1 vccd1 vccd1 _4926_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4857_ _6209_/Q _4768_/Y _4769_/Y _4850_/B _4815_/B vssd1 vssd1 vccd1 vccd1 _4857_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3278__B _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3808_ _6138_/Q _3808_/B _3808_/C vssd1 vssd1 vccd1 vccd1 _3809_/B sky130_fd_sc_hd__nor3_1
XANTENNA__4752__B1 _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4788_ hold382/X _4787_/X _4927_/S vssd1 vssd1 vccd1 vccd1 _4788_/X sky130_fd_sc_hd__mux2_1
X_3739_ hold94/A hold74/A _3739_/S vssd1 vssd1 vccd1 vccd1 _3739_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5409_ _5408_/A _5408_/B _5408_/Y _3648_/Y vssd1 vssd1 vccd1 vccd1 _5409_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_2_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4329__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5623__S _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5471__A1 _5484_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5223__A1 _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5760_ hold464/X _5741_/Y _5759_/X _5767_/A vssd1 vssd1 vccd1 vccd1 _5760_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2972_ _5997_/Q vssd1 vssd1 vccd1 vccd1 _2972_/Y sky130_fd_sc_hd__inv_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ _5691_/A _5691_/B vssd1 vssd1 vccd1 vccd1 _5691_/X sky130_fd_sc_hd__or2_1
XANTENNA__4982__A0 _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4711_ _5944_/Q _5935_/Q _5927_/Q _6035_/Q _6112_/Q _5936_/Q vssd1 vssd1 vccd1 vccd1
+ _4711_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_44_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4642_ _4699_/A _4643_/B vssd1 vssd1 vccd1 vccd1 _4676_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4573_ _4572_/X _4571_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4865_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3524_ _3328_/Y _3523_/Y _5566_/S vssd1 vssd1 vccd1 vccd1 _3524_/X sky130_fd_sc_hd__o21a_1
X_6243_ _6243_/CLK _6243_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6243_/Q sky130_fd_sc_hd__dfstp_2
X_3455_ _4415_/A _3210_/C _4070_/B _3454_/Y _4618_/B vssd1 vssd1 vccd1 vccd1 _3455_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__5533__S _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6174_ _6178_/CLK _6174_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6174_/Q sky130_fd_sc_hd__dfstp_4
X_3386_ _4124_/B _5296_/S _5875_/B vssd1 vssd1 vccd1 vccd1 _3386_/X sky130_fd_sc_hd__and3_1
X_5125_ _6172_/Q _5104_/Y _5108_/Y _6236_/Q _5124_/X vssd1 vssd1 vccd1 vccd1 _5125_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5056_ _4223_/B _4239_/B _4251_/Y _5055_/X _5051_/X vssd1 vssd1 vccd1 vccd1 _5056_/X
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5462__A1 _6177_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4007_ _5046_/A _5407_/A _4007_/S vssd1 vssd1 vccd1 vccd1 _4008_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5214__B2 _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5765__A2 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5958_ _6151_/CLK _5958_/D vssd1 vssd1 vccd1 vccd1 _5958_/Q sky130_fd_sc_hd__dfxtp_1
X_4909_ _4908_/X _6154_/Q _4926_/S vssd1 vssd1 vccd1 vccd1 _4909_/X sky130_fd_sc_hd__mux2_1
X_5889_ hold633/X _5875_/X _5876_/Y _5888_/X vssd1 vssd1 vccd1 vccd1 _5889_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_90_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5205__A1 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4639__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5756__A2 _5771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3216__B1 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_14_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6030_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5508__A2 _5507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_5 _4448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3777_/A _4735_/A _3643_/A vssd1 vssd1 vccd1 vccd1 _3921_/A sky130_fd_sc_hd__and3_2
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _3507_/C _4417_/A vssd1 vssd1 vccd1 vccd1 _3171_/X sky130_fd_sc_hd__or2_1
XFILLER_0_83_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4247__A2 _3588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3455__B1 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5812_ _2989_/A _5811_/X _5832_/S vssd1 vssd1 vccd1 vccd1 _5812_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4955__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5743_ _4119_/A _4895_/B _4610_/X _5762_/C vssd1 vssd1 vccd1 vccd1 _5743_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5747__A2 _5771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2955_ _3302_/A vssd1 vssd1 vccd1 vccd1 _3498_/A sky130_fd_sc_hd__inv_2
X_5674_ _6067_/Q _5702_/A2 _5702_/B1 _5673_/X vssd1 vssd1 vccd1 vccd1 _5674_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4707__B1 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4625_ _6021_/Q _5966_/Q _6013_/Q _5946_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4625_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold511 _4694_/X vssd1 vssd1 vccd1 vccd1 _6067_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4556_ hold104/X hold147/X hold102/X _5962_/Q _5076_/A0 _4272_/B vssd1 vssd1 vccd1
+ vccd1 _4556_/X sky130_fd_sc_hd__mux4_1
Xhold500 _5320_/X vssd1 vssd1 vccd1 vccd1 _6163_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold544 _6197_/Q vssd1 vssd1 vccd1 vccd1 _5626_/A sky130_fd_sc_hd__clkbuf_2
Xhold522 _6136_/Q vssd1 vssd1 vccd1 vccd1 hold522/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold533 _4455_/X vssd1 vssd1 vccd1 vccd1 _6049_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3507_ _4398_/A _5502_/A _3507_/C _3507_/D vssd1 vssd1 vccd1 vccd1 _3508_/C sky130_fd_sc_hd__or4_2
Xhold555 _5772_/X vssd1 vssd1 vccd1 vccd1 _6219_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 _5757_/X vssd1 vssd1 vccd1 vccd1 _6216_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold577 _5466_/X vssd1 vssd1 vccd1 vccd1 _6177_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold588 _5918_/Q vssd1 vssd1 vccd1 vccd1 hold588/X sky130_fd_sc_hd__clkbuf_2
X_4487_ _5338_/C _5338_/D _4487_/C vssd1 vssd1 vccd1 vccd1 _4761_/A sky130_fd_sc_hd__nor3_2
X_6226_ _6243_/CLK _6226_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6226_/Q sky130_fd_sc_hd__dfstp_1
Xhold599 _6239_/Q vssd1 vssd1 vccd1 vccd1 _2989_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5132__B1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3438_ _4390_/A _2964_/Y _4043_/C vssd1 vssd1 vccd1 vccd1 _4054_/C sky130_fd_sc_hd__a21oi_2
XANTENNA__5683__A1 _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6157_ _6235_/CLK _6157_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6157_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ hold33/X _3353_/X _3372_/A vssd1 vssd1 vccd1 vccd1 _5978_/D sky130_fd_sc_hd__a21o_1
X_5108_ _5108_/A _5121_/A vssd1 vssd1 vccd1 vccd1 _5108_/Y sky130_fd_sc_hd__nor2_2
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6088_ _6227_/CLK _6088_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6088_/Q sky130_fd_sc_hd__dfrtp_2
X_5039_ _5039_/A _5039_/B vssd1 vssd1 vccd1 vccd1 _5039_/X sky130_fd_sc_hd__or2_1
XANTENNA__5199__B1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4946__A0 _6199_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5738__A2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4850__B _4850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4342__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput42 _6248_/Q vssd1 vssd1 vccd1 vccd1 io_out[28] sky130_fd_sc_hd__buf_12
Xoutput31 _6088_/Q vssd1 vssd1 vccd1 vccd1 io_out[18] sky130_fd_sc_hd__buf_12
Xoutput20 _6299_/X vssd1 vssd1 vccd1 vccd1 io_oeb[30] sky130_fd_sc_hd__buf_12
XFILLER_0_31_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4229__A2 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3437__B1 _5424_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_38_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5729__A2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3835__S1 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4410_ _5773_/A _4410_/B vssd1 vssd1 vccd1 vccd1 _4410_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5872__A _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5390_ _6173_/Q _5390_/B vssd1 vssd1 vccd1 vccd1 _5390_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_22_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4341_ hold108/X _3836_/X _4345_/S vssd1 vssd1 vccd1 vccd1 _4341_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4488__A _5875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4272_ _5296_/S _4272_/B vssd1 vssd1 vccd1 vccd1 _4272_/X sky130_fd_sc_hd__or2_1
X_6011_ _6152_/CLK _6011_/D vssd1 vssd1 vccd1 vccd1 _6011_/Q sky130_fd_sc_hd__dfxtp_1
X_3223_ _3715_/B _3135_/B _4417_/A _3131_/B _3221_/X vssd1 vssd1 vccd1 vccd1 _3223_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4000__B _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3676__B1 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3154_ _3154_/A _3154_/B _3154_/C _3153_/X vssd1 vssd1 vccd1 vccd1 _3158_/C sky130_fd_sc_hd__or4b_1
X_3085_ _4615_/B _4727_/B _3085_/C _4729_/A vssd1 vssd1 vccd1 vccd1 _3086_/C sky130_fd_sc_hd__or4_1
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout155_A _5164_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3987_ _6003_/Q _3724_/S _3986_/X _3616_/B vssd1 vssd1 vccd1 vccd1 _3988_/C sky130_fd_sc_hd__a211o_1
X_5726_ _3832_/Y _5715_/B _5715_/Y _5725_/X vssd1 vssd1 vccd1 vccd1 _5726_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_45_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3286__B _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5657_ _5658_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5659_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5353__B1 _5343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4608_ _4609_/A _4609_/B vssd1 vssd1 vccd1 vccd1 _4631_/B sky130_fd_sc_hd__or2_1
X_5588_ _6160_/Q _5507_/Y _5508_/X vssd1 vssd1 vccd1 vccd1 _5590_/B sky130_fd_sc_hd__o21ai_1
X_4539_ hold60/A _5910_/Q _5896_/Q _6008_/Q _5076_/A0 _4272_/B vssd1 vssd1 vccd1 vccd1
+ _4539_/X sky130_fd_sc_hd__mux4_1
XANTENNA__4398__A _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold341 _6079_/Q vssd1 vssd1 vccd1 vccd1 hold341/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _4835_/X vssd1 vssd1 vccd1 vccd1 _6081_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold330 _6084_/Q vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 _6088_/Q vssd1 vssd1 vccd1 vccd1 hold396/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _5205_/X vssd1 vssd1 vccd1 vccd1 _6119_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold374 _5177_/X vssd1 vssd1 vccd1 vccd1 _6117_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold363 _6113_/Q vssd1 vssd1 vccd1 vccd1 hold363/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6209_ _6211_/CLK _6209_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6209_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__3667__B1 _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout68_A _4926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5344__B1 _5343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3416__S _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3362__D _3503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5662__A4 _6199_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4622__A2 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3910_ _6139_/Q _6140_/Q _3910_/C vssd1 vssd1 vccd1 vccd1 _4007_/S sky130_fd_sc_hd__and3_1
X_4890_ _6061_/Q _4889_/X _5606_/S vssd1 vssd1 vccd1 vccd1 _4890_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3830__A0 _4522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3841_ _6117_/Q _3655_/B _3238_/Y vssd1 vssd1 vccd1 vccd1 _3841_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3818__C _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3772_ _6136_/Q _6137_/Q vssd1 vssd1 vccd1 vccd1 _3773_/B sky130_fd_sc_hd__xor2_1
XANTENNA__4386__B2 _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4386__A1 _5502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3387__A _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5511_ _5762_/A _5629_/B vssd1 vssd1 vccd1 vccd1 _5511_/X sky130_fd_sc_hd__or2_2
XANTENNA__6194__RESET_B fanout184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4710__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5442_ _5440_/X _5441_/X _5773_/A hold404/X vssd1 vssd1 vccd1 vccd1 _6175_/D sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6123__RESET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5373_ _5373_/A _5373_/B vssd1 vssd1 vccd1 vccd1 _5377_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__5107__A _5107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4324_ _3880_/X hold96/X _4327_/S vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__mux2_1
Xfanout128 _3050_/C vssd1 vssd1 vccd1 vccd1 _3426_/A sky130_fd_sc_hd__buf_4
Xfanout117 _5360_/A vssd1 vssd1 vccd1 vccd1 _4124_/A sky130_fd_sc_hd__clkbuf_8
Xfanout106 _3207_/X vssd1 vssd1 vccd1 vccd1 _5424_/B sky130_fd_sc_hd__clkbuf_8
X_4255_ hold250/X hold214/X _4255_/S vssd1 vssd1 vccd1 vccd1 _4255_/X sky130_fd_sc_hd__mux2_1
Xfanout139 hold654/X vssd1 vssd1 vccd1 vccd1 _5046_/A sky130_fd_sc_hd__buf_4
XANTENNA__3649__A0 _6113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4186_ _4186_/A _4186_/B vssd1 vssd1 vccd1 vccd1 _4187_/B sky130_fd_sc_hd__or2_2
X_3206_ _4460_/A _4415_/A vssd1 vssd1 vccd1 vccd1 _5838_/A sky130_fd_sc_hd__nor2_4
XFILLER_0_38_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3137_ _3137_/A _3182_/B vssd1 vssd1 vccd1 vccd1 _4460_/C sky130_fd_sc_hd__nor2_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3068_ _3434_/B _4116_/B vssd1 vssd1 vccd1 vccd1 _4728_/C sky130_fd_sc_hd__or2_2
XANTENNA__3389__D_N _3517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3585__C1 _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5709_ _5834_/D _5740_/B vssd1 vssd1 vccd1 vccd1 _5715_/B sky130_fd_sc_hd__or2_4
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold160 _4267_/X vssd1 vssd1 vccd1 vccd1 _5931_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 _6024_/Q vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold484_A _6114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold182 _5324_/X vssd1 vssd1 vccd1 vccd1 _6167_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 _4452_/X vssd1 vssd1 vccd1 vccd1 _6045_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold651_A _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5801__A1 _3707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3407__A3 _5093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5868__A1 _6116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4485__B _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4040_ _4615_/B _4040_/B vssd1 vssd1 vccd1 vccd1 _4416_/B sky130_fd_sc_hd__or2_1
XANTENNA__4843__A2 _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5991_ _6149_/CLK _5991_/D vssd1 vssd1 vccd1 vccd1 _5991_/Q sky130_fd_sc_hd__dfxtp_1
X_4942_ hold396/X _4941_/Y _5020_/S vssd1 vssd1 vccd1 vccd1 _4942_/X sky130_fd_sc_hd__mux2_1
X_4873_ _4870_/Y _4871_/X _4872_/X _4767_/X _6194_/Q vssd1 vssd1 vccd1 vccd1 _4873_/X
+ sky130_fd_sc_hd__o32a_1
XANTENNA__4006__A _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3824_ _3920_/A _5396_/B vssd1 vssd1 vccd1 vccd1 _3824_/X sky130_fd_sc_hd__and2_1
XFILLER_0_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3755_ _3757_/B vssd1 vssd1 vccd1 vccd1 _3755_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_6_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5308__A0 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3686_ _3687_/A _3687_/B vssd1 vssd1 vccd1 vccd1 _3686_/X sky130_fd_sc_hd__or2_1
XANTENNA__5859__B2 _5245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5425_ _5475_/S _5423_/Y _5426_/B _5414_/Y vssd1 vssd1 vccd1 vccd1 _5425_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_30_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5356_ _5356_/A _6165_/Q _5489_/C _5838_/A vssd1 vssd1 vccd1 vccd1 _5484_/S sky130_fd_sc_hd__and4_4
X_4307_ _4226_/X hold253/X _4309_/S vssd1 vssd1 vccd1 vccd1 _5970_/D sky130_fd_sc_hd__mux2_1
X_5287_ _5248_/Y _5284_/X _5286_/X vssd1 vssd1 vccd1 vccd1 _5287_/X sky130_fd_sc_hd__a21o_1
X_4238_ _4238_/A _4238_/B vssd1 vssd1 vccd1 vccd1 _4239_/B sky130_fd_sc_hd__or2_1
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4169_ _5922_/Q _3588_/X _3603_/X _6014_/Q vssd1 vssd1 vccd1 vccd1 _4169_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_69_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4350__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3193__C _3193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5181__S _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_39_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6256_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5786__A0 _6176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4589__A1 _4879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4133__S0 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4525__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4684__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5002__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3540_ _3540_/A _3540_/B vssd1 vssd1 vccd1 vccd1 _3540_/X sky130_fd_sc_hd__or2_1
XFILLER_0_24_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5210_ _5116_/A _4033_/X _5105_/B _5209_/X vssd1 vssd1 vccd1 vccd1 _5210_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5880__A input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3471_ _4737_/A _4398_/B _5838_/B _3469_/Y _3470_/Y vssd1 vssd1 vccd1 vccd1 _3471_/Y
+ sky130_fd_sc_hd__a311oi_1
XANTENNA__4513__A1 _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5710__B1 _5875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6190_ _6190_/CLK _6190_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6190_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5141_ _6206_/Q _5106_/Y _5122_/Y _2992_/A vssd1 vssd1 vccd1 vccd1 _5150_/A sky130_fd_sc_hd__a22o_1
XANTENNA__3721__C1 _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5072_ hold31/X _4219_/B _5772_/S vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__mux2_1
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4023_ _3654_/S _6141_/Q _3052_/A _4022_/X vssd1 vssd1 vccd1 vccd1 _4023_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4943__B _4943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5777__A0 _6239_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5120__A _5120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5974_ _6129_/CLK hold43/X fanout170/X vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dfrtp_1
X_4925_ _5694_/A _4924_/X _4911_/Y vssd1 vssd1 vccd1 vccd1 _4925_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4856_ _4856_/A _4856_/B vssd1 vssd1 vccd1 vccd1 _4856_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3278__C _3434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4201__B1 _3615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3807_ _6071_/Q _3809_/A vssd1 vssd1 vccd1 vccd1 _3807_/X sky130_fd_sc_hd__or2_1
XANTENNA__4752__A1 _5245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3555__A2 _5424_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4787_ _4786_/X _6054_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _4787_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3738_ hold191/X _3737_/X _4035_/S vssd1 vssd1 vccd1 vccd1 _5893_/D sky130_fd_sc_hd__mux2_1
X_3669_ hold116/X _3668_/X _4035_/S vssd1 vssd1 vccd1 vccd1 _3669_/X sky130_fd_sc_hd__mux2_1
X_5408_ _5408_/A _5408_/B vssd1 vssd1 vccd1 vccd1 _5408_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5339_ _5507_/A wire93/X vssd1 vssd1 vccd1 vccd1 _5457_/A sky130_fd_sc_hd__and2_4
XANTENNA__3712__C1 _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4345__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3469__B _4759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold614_A _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4743__A1 _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3929__S0 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3932__B _6119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output31_A _6088_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5208__C1 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2971_ _5958_/Q vssd1 vssd1 vccd1 vccd1 _2971_/Y sky130_fd_sc_hd__inv_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5690_ _5690_/A _5690_/B vssd1 vssd1 vccd1 vccd1 _5691_/B sky130_fd_sc_hd__and2_1
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4710_ hold423/X _4709_/X _5073_/S vssd1 vssd1 vccd1 vccd1 _4710_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_84_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5875__A _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4641_ _6214_/Q _4928_/B _4714_/S vssd1 vssd1 vccd1 vccd1 _4643_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4734__A1 _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4572_ hold161/X _5994_/Q _6002_/Q _5963_/Q _5076_/A0 _4272_/B vssd1 vssd1 vccd1
+ vccd1 _4572_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_12_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3523_ _3523_/A _3523_/B vssd1 vssd1 vccd1 vccd1 _3523_/Y sky130_fd_sc_hd__nor2_1
X_6242_ _6242_/CLK _6242_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6242_/Q sky130_fd_sc_hd__dfstp_2
X_3454_ _4077_/A _5424_/C vssd1 vssd1 vccd1 vccd1 _3454_/Y sky130_fd_sc_hd__nor2_1
X_6173_ _6247_/CLK _6173_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6173_/Q sky130_fd_sc_hd__dfstp_4
X_3385_ _4460_/A _4486_/B vssd1 vssd1 vccd1 vccd1 _3388_/B sky130_fd_sc_hd__and2_1
X_5124_ _5109_/Y _5115_/X _5117_/X _5106_/Y _6204_/Q vssd1 vssd1 vccd1 vccd1 _5124_/X
+ sky130_fd_sc_hd__a32o_1
X_5055_ _5055_/A _5055_/B _5055_/C _5055_/D vssd1 vssd1 vccd1 vccd1 _5055_/X sky130_fd_sc_hd__and4_1
XFILLER_0_79_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4006_ _5046_/A _6141_/Q vssd1 vssd1 vccd1 vccd1 _5407_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3473__A1 hold588/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5765__A3 _4990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5957_ _6151_/CLK _5957_/D vssd1 vssd1 vccd1 vccd1 _5957_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4422__B1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4973__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4908_ _5694_/A _4907_/X _4895_/Y vssd1 vssd1 vccd1 vccd1 _4908_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5888_ input7/X _5890_/B vssd1 vssd1 vccd1 vccd1 _5888_/X sky130_fd_sc_hd__and2_1
X_4839_ _6057_/Q _6058_/Q _4839_/C vssd1 vssd1 vccd1 vccd1 _4854_/B sky130_fd_sc_hd__and3_1
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout98_A _4765_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3161__B1 _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5679__B _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__6060__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4639__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4964__A1 _4104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4803__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4104__A _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_6 _5136_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3507_/C _4417_/A vssd1 vssd1 vccd1 vccd1 _3709_/B sky130_fd_sc_hd__nor2_2
Xci2406_z80_210 vssd1 vssd1 vccd1 vccd1 ci2406_z80_210/HI io_out[33] sky130_fd_sc_hd__conb_1
XANTENNA__3455__A1 _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5811_ _5810_/X _3832_/Y _5831_/S vssd1 vssd1 vccd1 vccd1 _5811_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4404__B1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4713__S _5914_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5742_ _5764_/B _5771_/S vssd1 vssd1 vccd1 vccd1 _5742_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2954_ _4398_/B vssd1 vssd1 vccd1 vccd1 _5360_/A sky130_fd_sc_hd__inv_2
XFILLER_0_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5673_ hold380/X _6201_/Q _5701_/S vssd1 vssd1 vccd1 vccd1 _5673_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4624_ hold62/A hold78/A _5921_/Q _6029_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4624_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold501 _6066_/Q vssd1 vssd1 vccd1 vccd1 hold501/X sky130_fd_sc_hd__dlygate4sd3_1
X_4555_ hold216/X hold98/A _5897_/Q _6009_/Q _5076_/A0 _4272_/B vssd1 vssd1 vccd1
+ vccd1 _4555_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold545 _5635_/X vssd1 vssd1 vccd1 vccd1 _6197_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout100_A _5341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 _5263_/X vssd1 vssd1 vccd1 vccd1 _6136_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 _6061_/Q vssd1 vssd1 vccd1 vccd1 hold534/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_3506_ _5319_/A _3517_/C _3506_/C vssd1 vssd1 vccd1 vccd1 _3506_/X sky130_fd_sc_hd__and3b_1
Xhold512 _6189_/Q vssd1 vssd1 vccd1 vccd1 hold512/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5544__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 _6174_/Q vssd1 vssd1 vccd1 vccd1 hold567/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold578 _6204_/Q vssd1 vssd1 vccd1 vccd1 hold578/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold556 _6165_/Q vssd1 vssd1 vccd1 vccd1 hold556/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4486_ _4486_/A _4486_/B _5424_/C _4486_/D vssd1 vssd1 vccd1 vccd1 _4487_/C sky130_fd_sc_hd__or4_1
X_6225_ _6243_/CLK _6225_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6225_/Q sky130_fd_sc_hd__dfstp_1
Xhold589 _3474_/Y vssd1 vssd1 vccd1 vccd1 _5956_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3437_ _5362_/B _3713_/A _5424_/C vssd1 vssd1 vccd1 vccd1 _3437_/Y sky130_fd_sc_hd__a21oi_1
X_6156_ _6238_/CLK _6156_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6156_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _4765_/A _3368_/B _3368_/C vssd1 vssd1 vccd1 vccd1 _3372_/A sky130_fd_sc_hd__and3_1
XANTENNA__4891__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5107_ _5107_/A _5107_/B vssd1 vssd1 vccd1 vccd1 _5121_/A sky130_fd_sc_hd__nand2_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5435__A2 _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6087_ _6251_/CLK _6087_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6087_/Q sky130_fd_sc_hd__dfrtp_2
X_3299_ _5838_/B _4618_/C vssd1 vssd1 vccd1 vccd1 _4737_/B sky130_fd_sc_hd__nand2_2
X_5038_ _5502_/A _6178_/Q _3920_/A vssd1 vssd1 vccd1 vccd1 _5039_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput43 _6249_/Q vssd1 vssd1 vccd1 vccd1 io_out[29] sky130_fd_sc_hd__buf_12
Xoutput32 _6089_/Q vssd1 vssd1 vccd1 vccd1 io_out[19] sky130_fd_sc_hd__buf_12
Xoutput21 _6299_/A vssd1 vssd1 vccd1 vccd1 io_oeb[31] sky130_fd_sc_hd__buf_12
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5674__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3702__S _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4634__B1 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4340_ hold219/X _3789_/X _4345_/S vssd1 vssd1 vccd1 vccd1 _6006_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_22_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4271_ hold153/X _4261_/X _4271_/S vssd1 vssd1 vccd1 vccd1 _4271_/X sky130_fd_sc_hd__mux2_1
X_3222_ _4765_/A _6127_/Q _4124_/A vssd1 vssd1 vccd1 vccd1 _3246_/A sky130_fd_sc_hd__o21ai_4
X_6010_ _6010_/CLK _6010_/D vssd1 vssd1 vccd1 vccd1 _6010_/Q sky130_fd_sc_hd__dfxtp_1
X_3153_ _6130_/Q _4725_/B _3121_/X _3123_/X _3137_/A vssd1 vssd1 vccd1 vccd1 _3153_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3084_ _4038_/B _3063_/X _3083_/Y _4486_/B vssd1 vssd1 vccd1 vccd1 _4729_/A sky130_fd_sc_hd__a31o_1
XANTENNA__4009__A _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout148_A _3302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3986_ _3573_/C _3986_/A2 _3584_/X _3585_/X _5964_/Q vssd1 vssd1 vccd1 vccd1 _3986_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5725_ _4119_/A _4821_/B _4531_/Y _5762_/C vssd1 vssd1 vccd1 vccd1 _5725_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_45_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3567__B _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5656_ _5647_/A _5655_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _5656_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5353__A1 _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4607_ _4592_/B _4594_/B _4590_/X vssd1 vssd1 vccd1 vccd1 _4609_/B sky130_fd_sc_hd__a21oi_1
Xhold320 _5020_/X vssd1 vssd1 vccd1 vccd1 _6093_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5274__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5587_ hold421/X _5586_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _5587_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4538_ _4589_/S _4538_/B vssd1 vssd1 vccd1 vccd1 _4543_/B sky130_fd_sc_hd__nand2_1
Xhold353 _6252_/Q vssd1 vssd1 vccd1 vccd1 hold353/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold342 _4804_/X vssd1 vssd1 vccd1 vccd1 _6079_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold331 _4878_/X vssd1 vssd1 vccd1 vccd1 _6084_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold386 _6251_/Q vssd1 vssd1 vccd1 vccd1 hold386/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 _6250_/Q vssd1 vssd1 vccd1 vccd1 hold375/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold364 _5128_/X vssd1 vssd1 vccd1 vccd1 _6113_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4539__S0 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4469_ _4468_/X _4467_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4779_/B sky130_fd_sc_hd__mux2_4
Xhold397 _4942_/X vssd1 vssd1 vccd1 vccd1 _6088_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6208_ _6208_/CLK _6208_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6208_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_99_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6139_ _6175_/CLK _6139_/D vssd1 vssd1 vccd1 vccd1 _6139_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3419__A1 _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4711__S0 _6112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4353__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5344__A1 _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5184__S _5185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4855__B1 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3840_ _6139_/Q _3840_/B vssd1 vssd1 vccd1 vccd1 _5386_/A sky130_fd_sc_hd__xor2_2
X_3771_ _6173_/Q _2975_/Y _3912_/B vssd1 vssd1 vccd1 vccd1 _3773_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_73_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3387__B _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5510_ _4474_/A _5506_/X _5508_/X _5509_/Y _5875_/B vssd1 vssd1 vccd1 vccd1 _5629_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_89_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5441_ _3832_/A _5326_/X _5773_/A vssd1 vssd1 vccd1 vccd1 _5441_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3607__S _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5372_ _5372_/A _5372_/B vssd1 vssd1 vccd1 vccd1 _5378_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4323_ _3836_/X hold197/X _4327_/S vssd1 vssd1 vccd1 vccd1 _4323_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout129 _3050_/C vssd1 vssd1 vccd1 vccd1 _5868_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout107 _5838_/A vssd1 vssd1 vccd1 vccd1 _4618_/B sky130_fd_sc_hd__clkbuf_8
Xfanout118 _2950_/Y vssd1 vssd1 vccd1 vccd1 _4398_/A sky130_fd_sc_hd__buf_4
X_4254_ hold153/X hold110/X _4255_/S vssd1 vssd1 vccd1 vccd1 _4254_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3649__A1 _6117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4846__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4185_ _5948_/Q _3605_/X _3615_/X hold173/X _4184_/X vssd1 vssd1 vccd1 vccd1 _4186_/B
+ sky130_fd_sc_hd__a221o_1
X_3205_ _6129_/Q _3205_/B vssd1 vssd1 vccd1 vccd1 _3234_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3136_ _4726_/D wire93/A vssd1 vssd1 vccd1 vccd1 _3477_/A sky130_fd_sc_hd__or2_1
X_3067_ _3182_/B _3507_/D vssd1 vssd1 vccd1 vccd1 _4116_/B sky130_fd_sc_hd__nor2_2
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3821__A1 _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5269__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5708_ _5790_/C _5790_/D _5834_/C _5327_/B vssd1 vssd1 vccd1 vccd1 _5740_/B sky130_fd_sc_hd__or4b_1
X_3969_ _3988_/A _3963_/X _3968_/X vssd1 vssd1 vccd1 vccd1 _3970_/B sky130_fd_sc_hd__a21o_2
X_5639_ _5660_/A _5640_/B vssd1 vssd1 vccd1 vccd1 _5639_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_13_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold150 _4312_/X vssd1 vssd1 vccd1 vccd1 _5981_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 _5986_/Q vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 _6033_/Q vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 _4360_/X vssd1 vssd1 vccd1 vccd1 _6024_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 _5999_/Q vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout80_A _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3760__B _6115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4348__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5179__S _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4811__S _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3670__B _3671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5878__A input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5990_ _6006_/CLK hold89/X vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__dfxtp_1
X_4941_ _5704_/S _4939_/X _4940_/Y vssd1 vssd1 vccd1 vccd1 _4941_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_91_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4872_ _6160_/Q _5008_/B _4868_/X _4999_/A1 vssd1 vssd1 vccd1 vccd1 _4872_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_59_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3823_ _6137_/Q _6139_/Q _5868_/S vssd1 vssd1 vccd1 vccd1 _5396_/B sky130_fd_sc_hd__mux2_1
XANTENNA__5556__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4006__B _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6110_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3754_ _3988_/A _3753_/X _3750_/Y _3748_/Y vssd1 vssd1 vccd1 vccd1 _3757_/B sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3685_ _3636_/A _3636_/B _3628_/B vssd1 vssd1 vccd1 vccd1 _3687_/B sky130_fd_sc_hd__a21o_1
XANTENNA__5859__A2 _5836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5118__A _5120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4022__A _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3319__B1 _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5424_ _5424_/A _5424_/B _5424_/C vssd1 vssd1 vccd1 vccd1 _5426_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5355_ _5341_/A _5354_/Y _5352_/Y _6173_/Q vssd1 vssd1 vccd1 vccd1 _5355_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4306_ _4211_/X hold234/X _4309_/S vssd1 vssd1 vccd1 vccd1 _5969_/D sky130_fd_sc_hd__mux2_1
X_5286_ _6210_/Q _5251_/Y _5252_/Y _5767_/B _5285_/X vssd1 vssd1 vccd1 vccd1 _5286_/X
+ sky130_fd_sc_hd__a221o_1
X_4237_ _4236_/B _4237_/B vssd1 vssd1 vccd1 vccd1 _4238_/B sky130_fd_sc_hd__and2b_1
XANTENNA__5492__A0 _6238_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4168_ hold66/X _3611_/X _3613_/X hold54/X _4167_/X vssd1 vssd1 vccd1 vccd1 _4171_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5244__B1 _4409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4099_ _5078_/A _4099_/B _4099_/C vssd1 vssd1 vccd1 vccd1 _4099_/X sky130_fd_sc_hd__or3_1
XANTENNA__4047__A1 _4439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3119_ _3210_/A _3148_/B _3426_/A _3249_/A _4056_/B vssd1 vssd1 vccd1 vccd1 _3120_/B
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5547__A1 _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_hold594_A _6240_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4133__S1 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3946__A _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4541__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3470_ _3540_/A _4446_/A _3246_/A _3468_/X vssd1 vssd1 vccd1 vccd1 _3470_/Y sky130_fd_sc_hd__o31ai_1
XANTENNA__5171__C1 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5140_ _5164_/A1 hold484/X _5086_/Y _5139_/X vssd1 vssd1 vccd1 vccd1 _5140_/X sky130_fd_sc_hd__a22o_1
X_5071_ hold29/X _4203_/Y _5772_/S vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__mux2_1
X_4022_ _5868_/S _6135_/Q vssd1 vssd1 vccd1 vccd1 _4022_/X sky130_fd_sc_hd__and2_1
X_5973_ _6038_/CLK hold41/X fanout170/X vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4924_ _6063_/Q _5702_/A2 _5607_/B1 _4923_/X vssd1 vssd1 vccd1 vccd1 _4924_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5120__B _5185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4017__A _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3788__B1 _3671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4855_ _6059_/Q _4854_/B _4824_/B vssd1 vssd1 vccd1 vccd1 _4856_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3806_ _3808_/B _3808_/C _6138_/Q vssd1 vssd1 vccd1 vccd1 _3809_/A sky130_fd_sc_hd__o21a_1
X_4786_ _4119_/B _4785_/X _4757_/Y vssd1 vssd1 vccd1 vccd1 _4786_/X sky130_fd_sc_hd__a21bo_1
X_3737_ _4034_/S hold659/X _3735_/Y _3736_/X vssd1 vssd1 vccd1 vccd1 _3737_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3668_ _4034_/S _3595_/X _3666_/Y _3667_/Y vssd1 vssd1 vccd1 vccd1 _3668_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5407_ _5407_/A _5407_/B vssd1 vssd1 vccd1 vccd1 _5408_/B sky130_fd_sc_hd__xnor2_1
X_3599_ _3988_/A _3616_/B _3724_/S vssd1 vssd1 vccd1 vccd1 _3599_/X sky130_fd_sc_hd__and3_4
XFILLER_0_2_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3591__A _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5338_ _5338_/A _5338_/B _5338_/C _5338_/D vssd1 vssd1 vccd1 vccd1 _5338_/Y sky130_fd_sc_hd__nor4_1
XANTENNA__5465__A0 _3926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5269_ _3800_/B _4187_/B _5289_/S vssd1 vssd1 vccd1 vccd1 _5269_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_18_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4626__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5768__A1 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4440__A1 _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4361__S _4363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3929__S1 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4536__S _4598_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5759__A1 _3926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5208__B1 _3739_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3482__A2 _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2970_ _6074_/Q vssd1 vssd1 vccd1 vccd1 _3533_/S sky130_fd_sc_hd__inv_2
XANTENNA__4431__A1 _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5367__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5875__B _5875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4271__S _4271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4640_ _4639_/X _4638_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4928_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4571_ _6151_/Q _5912_/Q _5898_/Q _6010_/Q _5076_/A0 _4272_/B vssd1 vssd1 vccd1 vccd1
+ _4571_/X sky130_fd_sc_hd__mux4_1
X_3522_ _5317_/A _3520_/Y _5498_/C _3328_/B _5498_/A vssd1 vssd1 vccd1 vccd1 _3522_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6241_ _6242_/CLK _6241_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6241_/Q sky130_fd_sc_hd__dfstp_2
X_3453_ _4094_/B _3450_/X _3451_/X _3452_/X _4485_/B vssd1 vssd1 vccd1 vccd1 _3453_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6172_ _6247_/CLK _6172_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6172_/Q sky130_fd_sc_hd__dfstp_4
X_5123_ _2998_/Y _5129_/B _5121_/B vssd1 vssd1 vccd1 vccd1 _5123_/Y sky130_fd_sc_hd__o21ai_1
X_3384_ _5872_/A _5313_/S _3381_/Y _3405_/B vssd1 vssd1 vccd1 vccd1 _3384_/X sky130_fd_sc_hd__a211o_1
X_5054_ _5054_/A _5054_/B _5054_/C _5054_/D vssd1 vssd1 vccd1 vccd1 _5055_/D sky130_fd_sc_hd__and4_1
X_4005_ _4005_/A _4005_/B vssd1 vssd1 vccd1 vccd1 _4008_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout178_A fanout184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5956_ _6171_/CLK _5956_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _5956_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__4422__A1 _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4907_ _6062_/Q _4761_/X _5607_/B1 _4906_/X vssd1 vssd1 vccd1 vccd1 _4907_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_75_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5887_ _3643_/A _5875_/X _5876_/Y _5886_/X vssd1 vssd1 vccd1 vccd1 _6257_/D sky130_fd_sc_hd__o22a_1
X_4838_ _4836_/B _4837_/X _4963_/A vssd1 vssd1 vccd1 vccd1 _4838_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4769_ _4770_/A _4771_/C vssd1 vssd1 vccd1 vccd1 _4769_/Y sky130_fd_sc_hd__nor2_8
XANTENNA__4033__S0 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4356__S _4363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3464__A2 _5424_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3496__A _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3646__D _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4104__B _4104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_7 _5267_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5216__A _5216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_23_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6211_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4266__S _4271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_211 vssd1 vssd1 vccd1 vccd1 ci2406_z80_211/HI io_out[34] sky130_fd_sc_hd__conb_1
XANTENNA__4652__A1 _4507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3455__A2 _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_200 vssd1 vssd1 vccd1 vccd1 ci2406_z80_200/HI io_oeb[15] sky130_fd_sc_hd__conb_1
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5886__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6188__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5810_ hold398/X _5794_/Y _5809_/X _5794_/B vssd1 vssd1 vccd1 vccd1 _5810_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4404__A1 _5250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4955__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5741_ _5713_/A _5771_/S _5767_/A vssd1 vssd1 vccd1 vccd1 _5741_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2953_ _6259_/Q vssd1 vssd1 vccd1 vccd1 _3105_/A sky130_fd_sc_hd__inv_2
XFILLER_0_17_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5672_ _5658_/A _5671_/Y _5672_/S vssd1 vssd1 vccd1 vccd1 _5672_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4168__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4707__A2 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4623_ _5767_/A hold390/X _4621_/X _4622_/Y vssd1 vssd1 vccd1 vccd1 _4623_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold502 _4682_/X vssd1 vssd1 vccd1 vccd1 _6066_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4554_ _6159_/Q _4589_/S vssd1 vssd1 vccd1 vccd1 _4559_/B sky130_fd_sc_hd__nand2b_1
Xhold535 _4599_/X vssd1 vssd1 vccd1 vccd1 _6061_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3505_ _3715_/B _6164_/Q _3383_/B hold503/X vssd1 vssd1 vccd1 vccd1 _3505_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3391__A1 _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold524 _6053_/Q vssd1 vssd1 vccd1 vccd1 _2967_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold513 _5534_/X vssd1 vssd1 vccd1 vccd1 _6189_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6224_ _6243_/CLK _6224_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6224_/Q sky130_fd_sc_hd__dfstp_1
Xhold557 _6214_/Q vssd1 vssd1 vccd1 vccd1 hold557/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 _5429_/X vssd1 vssd1 vccd1 vccd1 _6174_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold579 _5718_/X vssd1 vssd1 vccd1 vccd1 _6204_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold546 _6058_/Q vssd1 vssd1 vccd1 vccd1 hold546/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4485_ _4485_/A _4485_/B vssd1 vssd1 vccd1 vccd1 _4486_/D sky130_fd_sc_hd__nand2_1
XANTENNA__5132__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3436_ _3446_/A _4618_/C vssd1 vssd1 vccd1 vccd1 _5424_/C sky130_fd_sc_hd__nand2_8
X_6155_ _6235_/CLK _6155_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6155_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5560__S _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3367_ hold244/X _3353_/X _3366_/X hold50/X vssd1 vssd1 vccd1 vccd1 _3402_/B sky130_fd_sc_hd__a22o_1
X_5106_ _5129_/A _5122_/B vssd1 vssd1 vccd1 vccd1 _5106_/Y sky130_fd_sc_hd__nor2_2
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6086_ _6086_/CLK _6086_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6086_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5037_ _5394_/A _5394_/B _5036_/X _5502_/A vssd1 vssd1 vccd1 vccd1 _5039_/A sky130_fd_sc_hd__o31a_1
X_3298_ _3298_/A _3540_/B vssd1 vssd1 vccd1 vccd1 _3298_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__5840__A0 _6113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5199__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5939_ _6110_/CLK hold67/X vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput33 _5875_/A vssd1 vssd1 vccd1 vccd1 io_out[1] sky130_fd_sc_hd__buf_12
Xoutput22 _2969_/Y vssd1 vssd1 vccd1 vccd1 io_out[0] sky130_fd_sc_hd__buf_12
XFILLER_0_31_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput44 _6153_/Q vssd1 vssd1 vccd1 vccd1 io_out[2] sky130_fd_sc_hd__buf_12
XANTENNA__3437__A2 _3713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4270_ hold80/X _4242_/X _4271_/S vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__mux2_1
X_3221_ _4765_/A _6127_/Q _4124_/A vssd1 vssd1 vccd1 vccd1 _3221_/X sky130_fd_sc_hd__o21a_2
XANTENNA__3676__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3152_ _4043_/A _3277_/A _3126_/X _3124_/Y vssd1 vssd1 vccd1 vccd1 _3158_/B sky130_fd_sc_hd__a31o_1
X_3083_ _3193_/A _3643_/B vssd1 vssd1 vccd1 vccd1 _3083_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_89_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4009__B _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3985_ _5987_/Q _3724_/S _3984_/X _3983_/S vssd1 vssd1 vccd1 vccd1 _3988_/B sky130_fd_sc_hd__a211o_1
X_5724_ hold470/X _5714_/Y _5723_/X _5767_/A vssd1 vssd1 vccd1 vccd1 _5724_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5655_ _5654_/X _5649_/Y _5670_/A vssd1 vssd1 vccd1 vccd1 _5655_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4606_ _4647_/A _4606_/B vssd1 vssd1 vccd1 vccd1 _4609_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5353__A2 _3193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5586_ _5579_/X _5585_/X _5670_/A vssd1 vssd1 vccd1 vccd1 _5586_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold310 _4820_/X vssd1 vssd1 vccd1 vccd1 _6080_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 _6186_/Q vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__buf_1
Xhold343 _6089_/Q vssd1 vssd1 vccd1 vccd1 hold343/X sky130_fd_sc_hd__dlygate4sd3_1
X_4537_ hold540/X _4536_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _4537_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold321 _5958_/Q vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 _5867_/X vssd1 vssd1 vccd1 vccd1 _6250_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 _5871_/X vssd1 vssd1 vccd1 vccd1 _6251_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 _6090_/Q vssd1 vssd1 vccd1 vccd1 hold365/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4539__S1 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4468_ _5980_/Q _5996_/Q _5988_/Q _5957_/Q _4272_/B _5076_/A0 vssd1 vssd1 vccd1 vccd1
+ _4468_/X sky130_fd_sc_hd__mux4_1
Xhold354 _5877_/X vssd1 vssd1 vccd1 vccd1 _6252_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 _6183_/Q vssd1 vssd1 vccd1 vccd1 hold398/X sky130_fd_sc_hd__dlygate4sd3_1
X_6207_ _6211_/CLK _6207_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6207_/Q sky130_fd_sc_hd__dfstp_2
X_3419_ _4038_/A _3172_/B _3237_/Y _3418_/X vssd1 vssd1 vccd1 vccd1 _3419_/X sky130_fd_sc_hd__a31o_1
X_6138_ _6175_/CLK _6138_/D vssd1 vssd1 vccd1 vccd1 _6138_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__4864__A1 _4863_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4399_ _4485_/B _4397_/X _4398_/X _5838_/A _4749_/A vssd1 vssd1 vccd1 vccd1 _4410_/B
+ sky130_fd_sc_hd__a32o_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ _6219_/CLK _6069_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6069_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__6039__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4711__S1 _5936_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4092__A2 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5041__A1 _6113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5344__A2 _3193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4552__A0 _6158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5280__A1 _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5280__B2 _6241_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3291__B1 _4116_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3770_ _2976_/Y _3647_/C _3764_/B _3769_/X vssd1 vssd1 vccd1 vccd1 _5375_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3387__C _5313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4791__B1 _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5440_ _3829_/Y _5363_/C _5439_/Y _5487_/S vssd1 vssd1 vccd1 vccd1 _5440_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5335__A2 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5371_ _3995_/B _3998_/Y _5370_/X vssd1 vssd1 vccd1 vccd1 _5371_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4322_ _3789_/X hold88/X _4327_/S vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__mux2_1
X_4253_ hold25/X _4253_/A2 _3671_/B vssd1 vssd1 vccd1 vccd1 _4253_/X sky130_fd_sc_hd__o21a_1
Xfanout119 _2950_/Y vssd1 vssd1 vccd1 vccd1 _3654_/S sky130_fd_sc_hd__buf_4
Xfanout108 _3894_/A vssd1 vssd1 vccd1 vccd1 _5024_/A sky130_fd_sc_hd__buf_4
XFILLER_0_10_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5099__A1 _3302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3204_ _3434_/B _3370_/B vssd1 vssd1 vccd1 vccd1 _3205_/B sky130_fd_sc_hd__nand2b_1
X_4184_ _5923_/Q _3588_/X _3603_/X _6015_/Q vssd1 vssd1 vccd1 vccd1 _4184_/X sky130_fd_sc_hd__a22o_1
X_3135_ _4398_/A _3135_/B _4417_/A _4051_/B vssd1 vssd1 vccd1 vccd1 wire93/A sky130_fd_sc_hd__nor4_1
XANTENNA__4059__C1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3066_ _4398_/A _3182_/A _3507_/C vssd1 vssd1 vccd1 vccd1 _3434_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_77_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3968_ _3968_/A _3968_/B _3968_/C vssd1 vssd1 vccd1 vccd1 _3968_/X sky130_fd_sc_hd__and3_1
X_5707_ _5698_/A _5706_/X _5707_/S vssd1 vssd1 vccd1 vccd1 _5707_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4782__B1 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3585__A1 _3513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3899_ _3899_/A _3899_/B vssd1 vssd1 vccd1 vccd1 _3900_/B sky130_fd_sc_hd__nand2_1
X_5638_ _5615_/X _5661_/A _5637_/X vssd1 vssd1 vccd1 vccd1 _5640_/B sky130_fd_sc_hd__a21o_1
X_5569_ _5569_/A _5569_/B vssd1 vssd1 vccd1 vccd1 _5569_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold151 _6020_/Q vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 _4296_/X vssd1 vssd1 vccd1 vccd1 _5960_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold162 _4317_/X vssd1 vssd1 vccd1 vccd1 _5986_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 _6031_/Q vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 _4370_/X vssd1 vssd1 vccd1 vccd1 _6033_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _4332_/X vssd1 vssd1 vccd1 vccd1 _5999_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5314__A _5314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold637_A _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4696__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5014__A1 _3270_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3488__B _3488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5014__B2 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3576__A1 _3513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4828__A1 _6157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4828__B2 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3500__B2 _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4940_ _6156_/Q _5704_/S vssd1 vssd1 vccd1 vccd1 _4940_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4871_ _6210_/Q _5009_/A2 _4769_/Y _4865_/B _4815_/B vssd1 vssd1 vccd1 vccd1 _4871_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3398__B _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3822_ _6116_/Q _6120_/Q _6070_/Q vssd1 vssd1 vccd1 vccd1 _5403_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3753_ _3751_/X _3752_/X _3983_/S vssd1 vssd1 vccd1 vccd1 _3753_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3618__S _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3684_ _3684_/A _3684_/B vssd1 vssd1 vccd1 vccd1 _3687_/A sky130_fd_sc_hd__and2_1
X_5423_ _5423_/A _5423_/B vssd1 vssd1 vccd1 vccd1 _5423_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__5118__B _5185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4022__B _6135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5354_ _5705_/S _5354_/B vssd1 vssd1 vccd1 vccd1 _5354_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4305_ _4193_/X hold248/X _4309_/S vssd1 vssd1 vccd1 vccd1 _4305_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5285_ _6160_/Q _5253_/Y _5254_/Y _6242_/Q vssd1 vssd1 vccd1 vccd1 _5285_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5134__A _5209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4236_ _4237_/B _4236_/B vssd1 vssd1 vccd1 vccd1 _4238_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4167_ _6022_/Q _3599_/X _3601_/X _5967_/Q vssd1 vssd1 vccd1 vccd1 _4167_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3118_ _3210_/A _3203_/B _3148_/C vssd1 vssd1 vccd1 vccd1 _4056_/B sky130_fd_sc_hd__or3_4
XFILLER_0_97_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5244__A1 _5250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4098_ _3221_/X _3442_/X _4084_/B _4097_/X vssd1 vssd1 vccd1 vccd1 _4099_/C sky130_fd_sc_hd__a211o_1
X_3049_ _3203_/A _4485_/A vssd1 vssd1 vccd1 vccd1 _3187_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3558__A1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_47_wb_clk_i_A _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4359__S _4363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6054__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5483__A1 _6179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5698__B _5698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4669__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5235__A1 _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4994__A0 _4990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_48_wb_clk_i _5978_/CLK vssd1 vssd1 vccd1 vccd1 _6144_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4746__B1 _4737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout90 _3536_/X vssd1 vssd1 vccd1 vccd1 _4034_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4777__B _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5710__A2 _6166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4269__S _4271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5070_ hold9/X _4187_/B _5073_/S vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__mux2_1
X_4021_ _6120_/Q _4021_/B vssd1 vssd1 vccd1 vccd1 _4021_/X sky130_fd_sc_hd__or2_1
XFILLER_0_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5972_ _6035_/CLK _5972_/D vssd1 vssd1 vccd1 vccd1 _5972_/Q sky130_fd_sc_hd__dfxtp_1
X_4923_ _6181_/Q _4922_/X _5701_/S vssd1 vssd1 vccd1 vccd1 _4923_/X sky130_fd_sc_hd__mux2_1
X_4854_ _6059_/Q _4854_/B vssd1 vssd1 vccd1 vccd1 _4856_/A sky130_fd_sc_hd__and2_1
XFILLER_0_7_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3805_ _5333_/B _3805_/B vssd1 vssd1 vccd1 vccd1 _3808_/C sky130_fd_sc_hd__nor2_1
X_4785_ _6054_/Q _5595_/S _5607_/B1 _4784_/X vssd1 vssd1 vccd1 vccd1 _4785_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_15_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3736_ hold11/X _4253_/A2 _3671_/B vssd1 vssd1 vccd1 vccd1 _3736_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3667_ _2999_/Y _3573_/B _4034_/S vssd1 vssd1 vccd1 vccd1 _3667_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5406_ _6139_/Q _6140_/Q vssd1 vssd1 vccd1 vccd1 _5407_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3598_ _5021_/B _3598_/B vssd1 vssd1 vccd1 vccd1 _4239_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_100_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5337_ _3650_/X _4005_/A _5334_/X _5025_/A _5336_/X vssd1 vssd1 vccd1 vccd1 _5337_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3591__B _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5268_ _5773_/A hold419/X _5245_/Y _5267_/X vssd1 vssd1 vccd1 vccd1 _5268_/X sky130_fd_sc_hd__a22o_1
X_4219_ _4219_/A _4219_/B vssd1 vssd1 vccd1 vccd1 _4220_/B sky130_fd_sc_hd__or2_1
X_5199_ _6018_/Q _5200_/A2 _5200_/B1 _5951_/Q _4256_/S vssd1 vssd1 vccd1 vccd1 _5201_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4208__A _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4440__A2 _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2951__A _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3951__A1 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_3_wb_clk_i_A _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5456__A1 _6177_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5502__A _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5759__A2 _5771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4552__S _4598_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4570_ _4589_/S _4570_/B vssd1 vssd1 vccd1 vccd1 _4575_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3395__C _6050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3521_ _4485_/B _4094_/B _4070_/B _4036_/B vssd1 vssd1 vccd1 vccd1 _5498_/C sky130_fd_sc_hd__and4_1
XFILLER_0_52_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6240_ _6243_/CLK _6240_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6240_/Q sky130_fd_sc_hd__dfstp_2
X_3452_ _3192_/B _3193_/X _3210_/C vssd1 vssd1 vccd1 vccd1 _3452_/X sky130_fd_sc_hd__a21o_1
X_6171_ _6171_/CLK _6171_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6171_/Q sky130_fd_sc_hd__dfrtp_1
X_3383_ _3383_/A _3383_/B vssd1 vssd1 vccd1 vccd1 _5313_/S sky130_fd_sc_hd__nand2_8
X_5122_ _5122_/A _5122_/B vssd1 vssd1 vccd1 vccd1 _5122_/Y sky130_fd_sc_hd__nor2_2
X_5053_ _5053_/A _5053_/B _5053_/C _5053_/D vssd1 vssd1 vccd1 vccd1 _5054_/D sky130_fd_sc_hd__and4_1
XANTENNA__3458__B1 _2960_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4004_ _5024_/A _5046_/A _6120_/Q _3848_/B _4003_/X vssd1 vssd1 vccd1 vccd1 _5372_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5558__S _5705_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5955_ _6171_/CLK _5955_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _5955_/Q sky130_fd_sc_hd__dfstp_1
X_4906_ _6180_/Q _4905_/X _5606_/S vssd1 vssd1 vccd1 vccd1 _4906_/X sky130_fd_sc_hd__mux2_1
X_5886_ input6/X _5890_/B vssd1 vssd1 vccd1 vccd1 _5886_/X sky130_fd_sc_hd__and2_1
XFILLER_0_90_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4837_ _6192_/Q _6058_/Q _5216_/A vssd1 vssd1 vccd1 vccd1 _4837_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4768_ _4771_/C _4770_/B _4770_/A vssd1 vssd1 vccd1 vccd1 _4768_/Y sky130_fd_sc_hd__nor3b_4
X_4699_ _4699_/A _4700_/B vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3719_ _3573_/C _3986_/A2 _3584_/X _3585_/X hold91/A vssd1 vssd1 vccd1 vccd1 _3719_/X
+ sky130_fd_sc_hd__o311a_1
XANTENNA__5135__B1 _5185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4033__S1 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4637__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__2946__A _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4372__S _4372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4104__C _5120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_8 _5506_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3017__A _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3152__A2 _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5429__A1 hold567/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xci2406_z80_212 vssd1 vssd1 vccd1 vccd1 ci2406_z80_212/HI io_out[35] sky130_fd_sc_hd__conb_1
XANTENNA__4652__A2 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3455__A3 _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_201 vssd1 vssd1 vccd1 vccd1 ci2406_z80_201/HI io_oeb[16] sky130_fd_sc_hd__conb_1
XFILLER_0_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4404__A2 _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5601__A1 _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5740_ _5740_/A _5740_/B vssd1 vssd1 vccd1 vccd1 _5771_/S sky130_fd_sc_hd__or2_4
X_2952_ _4061_/A vssd1 vssd1 vccd1 vccd1 _3694_/C sky130_fd_sc_hd__inv_6
XFILLER_0_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5671_ _5670_/A _5664_/Y _5670_/Y vssd1 vssd1 vccd1 vccd1 _5671_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4622_ _2984_/Y _4619_/X _5767_/A vssd1 vssd1 vccd1 vccd1 _4622_/Y sky130_fd_sc_hd__a21oi_1
X_4553_ hold546/X _4552_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _4553_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold525 _6199_/Q vssd1 vssd1 vccd1 vccd1 _5647_/A sky130_fd_sc_hd__buf_1
Xhold536 _6198_/Q vssd1 vssd1 vccd1 vccd1 _5636_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 _6232_/Q vssd1 vssd1 vccd1 vccd1 hold514/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5117__B1 _5105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3504_ _3504_/A _5566_/S _5216_/A vssd1 vssd1 vccd1 vccd1 _3517_/C sky130_fd_sc_hd__or3b_4
Xhold503 _6153_/Q vssd1 vssd1 vccd1 vccd1 hold503/X sky130_fd_sc_hd__dlygate4sd3_1
X_4484_ _4484_/A _4613_/A _4484_/C vssd1 vssd1 vccd1 vccd1 _5338_/D sky130_fd_sc_hd__or3_2
XFILLER_0_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5668__A1 _6158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6223_ _6251_/CLK _6223_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6223_/Q sky130_fd_sc_hd__dfstp_1
Xhold558 _5751_/X vssd1 vssd1 vccd1 vccd1 _6214_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold569 _6209_/Q vssd1 vssd1 vccd1 vccd1 hold569/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 _4553_/X vssd1 vssd1 vccd1 vccd1 _6058_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3435_ _4415_/A _4457_/B _3433_/X _4457_/A _3434_/X vssd1 vssd1 vccd1 vccd1 _5918_/D
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6154_ _6238_/CLK _6154_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6154_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3366_ _4474_/A _3368_/C vssd1 vssd1 vccd1 vccd1 _3366_/X sky130_fd_sc_hd__and2b_1
X_5105_ _5120_/A _5105_/B vssd1 vssd1 vccd1 vccd1 _5122_/B sky130_fd_sc_hd__or2_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ _6086_/CLK _6085_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6085_/Q sky130_fd_sc_hd__dfrtp_1
X_3297_ _4765_/A _4759_/B _4124_/A vssd1 vssd1 vccd1 vccd1 _3540_/B sky130_fd_sc_hd__o21ai_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5395_/A _5395_/B _5036_/C vssd1 vssd1 vccd1 vccd1 _5036_/X sky130_fd_sc_hd__or3_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5938_ _6030_/CLK hold63/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5869_ _6120_/Q _5868_/X _5869_/S vssd1 vssd1 vccd1 vccd1 _5869_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5317__A _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput34 _6090_/Q vssd1 vssd1 vccd1 vccd1 io_out[20] sky130_fd_sc_hd__buf_12
Xoutput23 _6080_/Q vssd1 vssd1 vccd1 vccd1 io_out[10] sky130_fd_sc_hd__buf_12
Xoutput45 _6250_/Q vssd1 vssd1 vccd1 vccd1 io_out[30] sky130_fd_sc_hd__buf_12
XANTENNA__4367__S _4372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5831__A1 _4030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4634__A2 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4095__B1 _3302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3842__B1 _6117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6204__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3300__A _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6250__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3970__A _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3220_ _4038_/A _3022_/B _3177_/Y vssd1 vssd1 vccd1 vccd1 _3220_/X sky130_fd_sc_hd__o21a_1
X_3151_ _3135_/B _4417_/B _4094_/B _3142_/Y vssd1 vssd1 vccd1 vccd1 _3154_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_89_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3082_ _4486_/A _3116_/A vssd1 vssd1 vccd1 vccd1 _3082_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4086__B1 _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3833__B1 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4389__A1 _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3984_ _3573_/C _3986_/A2 _3584_/X _3585_/X _5995_/Q vssd1 vssd1 vccd1 vccd1 _3984_/X
+ sky130_fd_sc_hd__o311a_1
X_5723_ _3785_/Y _5715_/B _5715_/Y _5722_/X vssd1 vssd1 vccd1 vccd1 _5723_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5654_ _5653_/X _5647_/A _5705_/S vssd1 vssd1 vccd1 vccd1 _5654_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4605_ _4699_/A _4605_/B vssd1 vssd1 vccd1 vccd1 _4606_/B sky130_fd_sc_hd__or2_1
XFILLER_0_72_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5353__A3 _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4010__B1 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5585_ _5592_/B _5585_/B vssd1 vssd1 vccd1 vccd1 _5585_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_53_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold311 _6086_/Q vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold300 _6036_/Q vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 _5496_/X vssd1 vssd1 vccd1 vccd1 _6186_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold344 _4958_/X vssd1 vssd1 vccd1 vccd1 _6089_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4536_ _6157_/Q _4535_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4536_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold322 _4294_/X vssd1 vssd1 vccd1 vccd1 _5958_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold366 _4975_/X vssd1 vssd1 vccd1 vccd1 _6090_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4976__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold355 _6247_/Q vssd1 vssd1 vccd1 vccd1 hold355/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 _5901_/Q vssd1 vssd1 vccd1 vccd1 hold377/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5902__RESET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4467_ hold84/A _5892_/Q hold86/A _6004_/Q _4272_/B _5076_/A0 vssd1 vssd1 vccd1 vccd1
+ _4467_/X sky130_fd_sc_hd__mux4_1
Xhold399 _5493_/X vssd1 vssd1 vccd1 vccd1 _6183_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold388 _6118_/Q vssd1 vssd1 vccd1 vccd1 hold388/X sky130_fd_sc_hd__buf_1
X_6206_ _6206_/CLK _6206_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6206_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_68_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3418_ _4094_/B _3192_/B _4036_/B _3417_/X vssd1 vssd1 vccd1 vccd1 _3418_/X sky130_fd_sc_hd__a31o_1
X_4398_ _4398_/A _4398_/B _4398_/C vssd1 vssd1 vccd1 vccd1 _4398_/X sky130_fd_sc_hd__or3_1
XANTENNA__5510__B1 _5875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6137_ _6175_/CLK _6137_/D vssd1 vssd1 vccd1 vccd1 _6137_/Q sky130_fd_sc_hd__dfxtp_4
X_3349_ _5566_/S _3503_/C vssd1 vssd1 vccd1 vccd1 _3349_/Y sky130_fd_sc_hd__nor2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ _6219_/CLK _6068_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6068_/Q sky130_fd_sc_hd__dfrtp_2
X_5019_ _5018_/X _6161_/Q _5704_/S vssd1 vssd1 vccd1 vccd1 _5019_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5344__A3 _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5501__B1 _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5804__A1 _6238_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5804__B2 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4825__S _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3014__B _3694_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4126__A _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5656__S _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4791__B2 _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3594__A2 _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5370_ _6142_/Q _5370_/B _3995_/B vssd1 vssd1 vccd1 vccd1 _5370_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_22_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4321_ _3737_/X hold90/X _4327_/S vssd1 vssd1 vccd1 vccd1 _5989_/D sky130_fd_sc_hd__mux2_1
X_4252_ _4239_/A _4251_/Y _4031_/Y vssd1 vssd1 vccd1 vccd1 _4252_/Y sky130_fd_sc_hd__o21bai_1
Xfanout109 _5875_/A vssd1 vssd1 vccd1 vccd1 _5296_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__4846__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3203_ _3203_/A _3203_/B _3203_/C _3203_/D vssd1 vssd1 vccd1 vccd1 _3370_/B sky130_fd_sc_hd__or4_4
X_4183_ _6023_/Q _3599_/X _3601_/X _5968_/Q _4182_/X vssd1 vssd1 vccd1 vccd1 _4186_/A
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3205__A _6129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3134_ _3426_/A _3150_/A _4117_/C vssd1 vssd1 vccd1 vccd1 _4726_/D sky130_fd_sc_hd__and3_4
XANTENNA__3806__B1 _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3065_ _3249_/B _3116_/A vssd1 vssd1 vccd1 vccd1 _4614_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4036__A _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4231__B1 _3615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3967_ _5898_/Q _3724_/S _3966_/X _3616_/B vssd1 vssd1 vccd1 vccd1 _3968_/C sky130_fd_sc_hd__a211o_1
X_5706_ _5699_/Y _5700_/X _5705_/X _5511_/X vssd1 vssd1 vccd1 vccd1 _5706_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5566__S _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4782__A1 _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3898_ _3898_/A _3898_/B vssd1 vssd1 vccd1 vccd1 _3900_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_45_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5637_ _6196_/Q _6197_/Q _5685_/B vssd1 vssd1 vccd1 vccd1 _5637_/X sky130_fd_sc_hd__o21a_1
X_5568_ _5569_/A _5569_/B vssd1 vssd1 vccd1 vccd1 _5584_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4534__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 _5924_/Q vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 _4356_/X vssd1 vssd1 vccd1 vccd1 _6020_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_37_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3742__C1 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4519_ _4517_/X _4518_/X _5872_/A vssd1 vssd1 vccd1 vccd1 _4519_/X sky130_fd_sc_hd__mux2_1
Xhold130 _6004_/Q vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 _4368_/X vssd1 vssd1 vccd1 vccd1 _6031_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 _5909_/Q vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _5998_/Q vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ _5609_/S _4761_/B _5498_/X _5872_/A vssd1 vssd1 vccd1 vccd1 _5499_/X sky130_fd_sc_hd__o31a_1
Xhold196 _6044_/Q vssd1 vssd1 vccd1 vccd1 _4129_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5314__B _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold365_A _6090_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout66_A _5711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4696__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold532_A _6047_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5330__A _5330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3785__A _3785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4773__A1 _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3724__S _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4828__A2 _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5789__A0 _6179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4870_ _6060_/Q _4856_/A _4869_/Y vssd1 vssd1 vccd1 vccd1 _4870_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3821_ _6173_/Q _3912_/C _3817_/Y _3820_/Y vssd1 vssd1 vccd1 vccd1 _5387_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_46_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4213__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4290__S _4291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3752_ _5998_/Q _5959_/Q _3982_/S vssd1 vssd1 vccd1 vccd1 _3752_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3683_ _6136_/Q _3683_/B _3683_/C vssd1 vssd1 vccd1 vccd1 _3684_/B sky130_fd_sc_hd__or3_1
X_5422_ _5422_/A _5422_/B vssd1 vssd1 vccd1 vccd1 _5423_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5353_ _5507_/A _3193_/C _4614_/B _5343_/X vssd1 vssd1 vccd1 vccd1 _5354_/B sky130_fd_sc_hd__a31oi_2
XFILLER_0_2_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5415__A _6157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4304_ _4180_/X hold100/X _4309_/S vssd1 vssd1 vccd1 vccd1 _4304_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_49_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5284_ _3970_/B _4233_/Y _5289_/S vssd1 vssd1 vccd1 vccd1 _5284_/X sky130_fd_sc_hd__mux2_1
X_4235_ _4207_/A _4207_/B _4222_/A _4220_/A _4206_/A vssd1 vssd1 vccd1 vccd1 _4237_/B
+ sky130_fd_sc_hd__o311a_1
X_4166_ hold209/X _4165_/X _4262_/S vssd1 vssd1 vccd1 vccd1 _4166_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3117_ _3643_/A _3081_/B _3192_/B _3052_/A _3116_/Y vssd1 vssd1 vccd1 vccd1 _3117_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5244__A2 _5250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3589__B _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4097_ _4485_/A _4750_/B _4094_/X _4096_/X _4416_/A vssd1 vssd1 vccd1 vccd1 _4097_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3048_ _3193_/C _3172_/B _4726_/B _3041_/Y _3411_/B vssd1 vssd1 vccd1 vccd1 _3057_/C
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4999_ _4999_/A1 _4994_/X _4998_/X _4824_/B vssd1 vssd1 vccd1 vccd1 _4999_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_80_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5180__A1 _3739_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5180__B2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold482_A _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4669__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout80 _5179_/S vssd1 vssd1 vccd1 vccd1 _5182_/S sky130_fd_sc_hd__clkbuf_8
Xfanout91 _3536_/X vssd1 vssd1 vccd1 vccd1 _4242_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__4746__B2 _5424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_17_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6033_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3721__A2 _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4020_ _6070_/Q _4021_/B vssd1 vssd1 vccd1 vccd1 _4020_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4285__S _4291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5971_ _6032_/CLK _5971_/D vssd1 vssd1 vccd1 vccd1 _5971_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_35_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4922_ _6197_/Q _4815_/B _4913_/X _4921_/X vssd1 vssd1 vccd1 vccd1 _4922_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3788__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4853_ _4850_/B _4852_/X _4963_/A vssd1 vssd1 vccd1 vccd1 _4853_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_51_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3804_ _5024_/A _6116_/Q vssd1 vssd1 vccd1 vccd1 _3808_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_7_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4784_ _6054_/Q _4783_/X _5606_/S vssd1 vssd1 vccd1 vccd1 _4784_/X sky130_fd_sc_hd__mux2_1
X_3735_ _5052_/A _3734_/X _3708_/X vssd1 vssd1 vccd1 vccd1 _3735_/Y sky130_fd_sc_hd__o21bai_1
XANTENNA__5844__S _5869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3960__A2 _3959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5162__A1 _6239_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5405_ _5405_/A _5405_/B vssd1 vssd1 vccd1 vccd1 _5408_/A sky130_fd_sc_hd__xnor2_1
X_3666_ _4223_/A _3620_/X _3665_/Y vssd1 vssd1 vccd1 vccd1 _3666_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3597_ _5021_/B _3598_/B vssd1 vssd1 vccd1 vccd1 _3597_/X sky130_fd_sc_hd__and2_2
XFILLER_0_100_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5336_ _6172_/Q _6073_/Q _3647_/B _3920_/A _5335_/X vssd1 vssd1 vccd1 vccd1 _5336_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_2_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5267_ _5248_/Y _5264_/X _5266_/X vssd1 vssd1 vccd1 vccd1 _5267_/X sky130_fd_sc_hd__a21o_1
X_4218_ _4219_/A _4219_/B vssd1 vssd1 vccd1 vccd1 _4220_/A sky130_fd_sc_hd__nand2_1
X_5198_ _5198_/A _5198_/B vssd1 vssd1 vccd1 vccd1 _5198_/X sky130_fd_sc_hd__or2_1
X_4149_ hold21/X _3539_/Y _3671_/B vssd1 vssd1 vccd1 vccd1 _4149_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_46_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3400__A1 _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4587__S0 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3164__B1 _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4664__B1 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5502__B _5502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5208__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4719__B2 _4474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3520_ _3405_/B _5314_/A _3503_/C vssd1 vssd1 vccd1 vccd1 _3520_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3451_ _3446_/A _4043_/C _3447_/X _3445_/X vssd1 vssd1 vccd1 vccd1 _3451_/X sky130_fd_sc_hd__a31o_1
X_3382_ _3382_/A _3383_/B vssd1 vssd1 vccd1 vccd1 _5875_/B sky130_fd_sc_hd__and2_4
X_6170_ _6170_/CLK _6170_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6170_/Q sky130_fd_sc_hd__dfrtp_1
X_5121_ _5121_/A _5121_/B vssd1 vssd1 vccd1 vccd1 _5121_/Y sky130_fd_sc_hd__nor2_2
X_5052_ _5052_/A _5052_/B _5052_/C _5052_/D vssd1 vssd1 vccd1 vccd1 _5053_/D sky130_fd_sc_hd__and4_1
XANTENNA__3458__A1 hold567/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4003_ _3848_/B _3997_/X _3998_/Y _4002_/X vssd1 vssd1 vccd1 vccd1 _4003_/X sky130_fd_sc_hd__a31o_1
X_5954_ _6171_/CLK _5954_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _5954_/Q sky130_fd_sc_hd__dfstp_1
X_4905_ _6196_/Q _4815_/B _4897_/X _4904_/X vssd1 vssd1 vccd1 vccd1 _4905_/X sky130_fd_sc_hd__a211o_1
X_5885_ _5356_/A _5875_/X _5876_/Y _5884_/X vssd1 vssd1 vccd1 vccd1 _6256_/D sky130_fd_sc_hd__o22a_1
XFILLER_0_47_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4836_ _4990_/A _4836_/B vssd1 vssd1 vccd1 vccd1 _4836_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5574__S _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4767_ _4771_/B _4770_/C vssd1 vssd1 vccd1 vccd1 _4767_/X sky130_fd_sc_hd__or2_2
X_4698_ _6218_/Q _4990_/B _4714_/S vssd1 vssd1 vccd1 vccd1 _4700_/B sky130_fd_sc_hd__mux2_1
X_3718_ _4234_/A vssd1 vssd1 vccd1 vccd1 _4250_/A sky130_fd_sc_hd__inv_4
XFILLER_0_31_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5135__A1 _5116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3649_ _6113_/Q _6117_/Q _6070_/Q vssd1 vssd1 vccd1 vccd1 _5404_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_101_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3697__B2 _6114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5319_ _5319_/A _5319_/B vssd1 vssd1 vccd1 vccd1 _5319_/X sky130_fd_sc_hd__or2_1
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
X_6299_ _6299_/A vssd1 vssd1 vccd1 vccd1 _6299_/X sky130_fd_sc_hd__buf_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3449__A1 _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4653__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5484__S _5484_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_9 _3498_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5126__A1 _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5429__A2 _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5513__A _6188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_202 vssd1 vssd1 vccd1 vccd1 ci2406_z80_202/HI io_oeb[17] sky130_fd_sc_hd__conb_1
XANTENNA__3033__A _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_213 vssd1 vssd1 vccd1 vccd1 io_oeb[32] ci2406_z80_213/LO sky130_fd_sc_hd__conb_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3968__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2951_ _3556_/A vssd1 vssd1 vccd1 vccd1 _4735_/A sky130_fd_sc_hd__inv_4
Xclkbuf_leaf_32_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6227_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5670_ _5670_/A _5670_/B vssd1 vssd1 vccd1 vccd1 _5670_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_84_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4621_ hold390/X _4612_/X _4619_/X _4611_/X vssd1 vssd1 vccd1 vccd1 _4621_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4168__A2 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4552_ _6158_/Q _4551_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4552_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold526 _5656_/X vssd1 vssd1 vccd1 vccd1 _6199_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 _5786_/X vssd1 vssd1 vccd1 vccd1 _6232_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5117__A1 _5209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold504 _3505_/X vssd1 vssd1 vccd1 vccd1 _3506_/C sky130_fd_sc_hd__dlygate4sd3_1
X_3503_ _4077_/A _6047_/Q _3503_/C _5218_/B vssd1 vssd1 vccd1 vccd1 _3504_/A sky130_fd_sc_hd__or4_1
X_4483_ _4483_/A _4483_/B _4613_/B vssd1 vssd1 vccd1 vccd1 _4484_/C sky130_fd_sc_hd__or3_1
X_6222_ _6242_/CLK _6222_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6222_/Q sky130_fd_sc_hd__dfstp_1
Xhold537 _5646_/X vssd1 vssd1 vccd1 vccd1 _6198_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 _6059_/Q vssd1 vssd1 vccd1 vccd1 hold559/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6126__RESET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3434_ _4124_/B _3434_/B _5875_/B _3434_/D vssd1 vssd1 vccd1 vccd1 _3434_/X sky130_fd_sc_hd__and4_1
Xhold548 _6055_/Q vssd1 vssd1 vccd1 vccd1 hold548/X sky130_fd_sc_hd__buf_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6153_ _6171_/CLK _6153_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6153_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_0_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3365_ hold44/X _3353_/X _3364_/Y vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__a21o_1
X_5104_ _5129_/A _5108_/A vssd1 vssd1 vccd1 vccd1 _5104_/Y sky130_fd_sc_hd__nor2_2
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3296_ _4451_/C _4759_/B _4124_/A vssd1 vssd1 vccd1 vccd1 _3296_/X sky130_fd_sc_hd__o21a_1
X_6084_ _6086_/CLK _6084_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6084_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5396_/A _5396_/B _5397_/A _5397_/B vssd1 vssd1 vccd1 vccd1 _5036_/C sky130_fd_sc_hd__or4_1
XANTENNA_fanout183_A fanout184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5937_ _6149_/CLK _5937_/D vssd1 vssd1 vccd1 vccd1 _5937_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5868_ _6138_/Q _6116_/Q _5868_/S vssd1 vssd1 vccd1 vccd1 _5868_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5799_ _6237_/Q _5791_/X _5798_/X _5764_/B vssd1 vssd1 vccd1 vccd1 _5799_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_63_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4819_ _4818_/X _6056_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _4819_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput24 _6081_/Q vssd1 vssd1 vccd1 vccd1 io_out[11] sky130_fd_sc_hd__buf_12
XFILLER_0_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput46 _6251_/Q vssd1 vssd1 vccd1 vccd1 io_out[31] sky130_fd_sc_hd__buf_12
Xoutput35 _6091_/Q vssd1 vssd1 vccd1 vccd1 io_out[21] sky130_fd_sc_hd__buf_12
XFILLER_0_31_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2957__A _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4619__B1 _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4095__A1 _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5347__B2 _3377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5347__A1 _6172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3150_ _3150_/A _4094_/B vssd1 vssd1 vccd1 vccd1 _3439_/B sky130_fd_sc_hd__nand2_2
X_3081_ _3135_/B _3081_/B _3178_/B vssd1 vssd1 vccd1 vccd1 _4486_/B sky130_fd_sc_hd__and3_2
XFILLER_0_89_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4293__S _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5722_ _4119_/A _4805_/B _4516_/Y _5762_/C vssd1 vssd1 vccd1 vccd1 _5722_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3983_ _3981_/X _3982_/X _3983_/S vssd1 vssd1 vccd1 vccd1 _3983_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5653_ _5652_/X _6157_/Q _5704_/S vssd1 vssd1 vccd1 vccd1 _5653_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5418__A _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4604_ _4699_/A _4605_/B vssd1 vssd1 vccd1 vccd1 _4647_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5584_ _5584_/A _5584_/B _5582_/Y vssd1 vssd1 vccd1 vccd1 _5585_/B sky130_fd_sc_hd__or3b_1
XANTENNA__4010__A1 _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4535_ _4533_/X _4534_/X _5872_/A vssd1 vssd1 vccd1 vccd1 _4535_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold301 _3430_/X vssd1 vssd1 vccd1 vccd1 _6036_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_27_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xhold334 _6248_/Q vssd1 vssd1 vccd1 vccd1 hold334/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 _6249_/Q vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5852__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold312 _4910_/X vssd1 vssd1 vccd1 vccd1 _6086_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold345 _6092_/Q vssd1 vssd1 vccd1 vccd1 hold345/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4976__B _4976_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold356 _5855_/X vssd1 vssd1 vccd1 vccd1 _6247_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold378 _3424_/X vssd1 vssd1 vccd1 vccd1 hold378/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 _5905_/Q vssd1 vssd1 vccd1 vccd1 hold367/X sky130_fd_sc_hd__dlygate4sd3_1
X_4466_ _4497_/S _4466_/B vssd1 vssd1 vccd1 vccd1 _4598_/S sky130_fd_sc_hd__nand2_4
Xhold389 _5192_/X vssd1 vssd1 vccd1 vccd1 _6118_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6210__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6205_ _6208_/CLK _6205_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6205_/Q sky130_fd_sc_hd__dfstp_2
X_4397_ _3426_/A _6127_/Q _5502_/C _4396_/X vssd1 vssd1 vccd1 vccd1 _4397_/X sky130_fd_sc_hd__a31o_1
X_3417_ _3105_/A _4070_/B _4085_/B _4439_/A _3276_/A vssd1 vssd1 vccd1 vccd1 _3417_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__5510__A1 _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6136_ _6175_/CLK _6136_/D vssd1 vssd1 vccd1 vccd1 _6136_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3348_ _3513_/A _3383_/B vssd1 vssd1 vccd1 vccd1 _3503_/C sky130_fd_sc_hd__nor2_4
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ _6219_/CLK _6067_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6067_/Q sky130_fd_sc_hd__dfrtp_4
X_3279_ _3484_/A _5502_/D _3279_/C vssd1 vssd1 vccd1 vccd1 _3281_/B sky130_fd_sc_hd__or3_1
X_5018_ _5694_/A _5017_/X _5007_/Y vssd1 vssd1 vccd1 vccd1 _5018_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__5299__S _5305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5577__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4931__S _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold408_A _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4378__S _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4068__A1 _5502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5017__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4791__A2 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5672__S _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4320_ _3668_/X hold189/X _4327_/S vssd1 vssd1 vccd1 vccd1 _4320_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4288__S _4291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4251_ _4251_/A _4251_/B vssd1 vssd1 vccd1 vccd1 _4251_/Y sky130_fd_sc_hd__xnor2_1
X_3202_ _3177_/Y _3200_/X _3201_/X _3164_/Y vssd1 vssd1 vccd1 vccd1 _3218_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_38_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4182_ hold82/A _3611_/X _3613_/X _5931_/Q vssd1 vssd1 vccd1 vccd1 _4182_/X sky130_fd_sc_hd__a22o_1
X_3133_ _5502_/D _4772_/B vssd1 vssd1 vccd1 vccd1 _3478_/A sky130_fd_sc_hd__or2_1
XANTENNA__4059__A1 _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3064_ _3203_/A _3148_/B _3148_/C vssd1 vssd1 vccd1 vccd1 _3116_/A sky130_fd_sc_hd__or3_4
XFILLER_0_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4036__B _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3966_ _3573_/C _3986_/A2 _3584_/X _3585_/X _6010_/Q vssd1 vssd1 vccd1 vccd1 _3966_/X
+ sky130_fd_sc_hd__o311a_1
X_5705_ _5704_/X _5698_/A _5705_/S vssd1 vssd1 vccd1 vccd1 _5705_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4782__A2 _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5636_ _5636_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5660_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3897_ _6140_/Q _3897_/B _3897_/C vssd1 vssd1 vccd1 vccd1 _3898_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_45_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5731__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5567_ _6158_/Q _5507_/Y _5508_/X vssd1 vssd1 vccd1 vccd1 _5569_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__5731__A1 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold153 _5935_/Q vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 _4212_/X vssd1 vssd1 vccd1 vccd1 _5924_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 _5910_/Q vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3742__B1 _3739_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5498_ _5498_/A _5498_/B _5498_/C vssd1 vssd1 vccd1 vccd1 _5498_/X sky130_fd_sc_hd__or3_2
Xhold131 _4338_/X vssd1 vssd1 vccd1 vccd1 _6004_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ hold542/X input3/X _4596_/S vssd1 vssd1 vccd1 vccd1 _4518_/X sky130_fd_sc_hd__mux2_1
Xhold175 _5933_/Q vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 _6022_/Q vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _4111_/X vssd1 vssd1 vccd1 vccd1 _5909_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4449_ _4124_/A _3488_/B _4429_/X _3426_/A vssd1 vssd1 vccd1 vccd1 _4449_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5495__A0 _6241_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold197 _5991_/Q vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4926__S _4926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6119_ _6119_/CLK _6119_/D vssd1 vssd1 vccd1 vccd1 _6119_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout59_A _5707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold525_A _6199_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4758__C1 _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4773__A2 _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5492__S _5497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5722__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5722__A1 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3740__S _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3820_ _3820_/A _3820_/B vssd1 vssd1 vccd1 vccd1 _3820_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3976__A _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3751_ _5982_/Q hold88/A _3982_/S vssd1 vssd1 vccd1 vccd1 _3751_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3972__B1 _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3682_ _5024_/A _3684_/A vssd1 vssd1 vccd1 vccd1 _3682_/Y sky130_fd_sc_hd__nand2_1
X_5421_ _6155_/Q _6154_/Q vssd1 vssd1 vccd1 vccd1 _5422_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__3915__S _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5352_ _5352_/A vssd1 vssd1 vccd1 vccd1 _5352_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5415__B _6156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4303_ _4165_/X hold238/X _4309_/S vssd1 vssd1 vccd1 vccd1 _5966_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_10_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5283_ _5773_/A hold406/X _5245_/Y _5282_/X vssd1 vssd1 vccd1 vccd1 _5283_/X sky130_fd_sc_hd__a22o_1
X_4234_ _4234_/A _4234_/B vssd1 vssd1 vccd1 vccd1 _4236_/B sky130_fd_sc_hd__xnor2_1
X_4165_ _4242_/S _4164_/X _4163_/X vssd1 vssd1 vccd1 vccd1 _4165_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3116_ _3116_/A _3116_/B vssd1 vssd1 vccd1 vccd1 _3116_/Y sky130_fd_sc_hd__nor2_1
X_4096_ _4061_/A _3477_/B _4095_/X _3543_/B _3082_/Y vssd1 vssd1 vccd1 vccd1 _4096_/X
+ sky130_fd_sc_hd__a32o_1
X_3047_ _3135_/B _3184_/A vssd1 vssd1 vccd1 vccd1 _4726_/B sky130_fd_sc_hd__and2_1
XANTENNA__4452__A1 _5164_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5792__A2_N _5352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4998_ _6160_/Q _4997_/Y _5013_/S vssd1 vssd1 vccd1 vccd1 _4998_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5401__B1 _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3949_ _3945_/Y _3948_/Y _6173_/Q vssd1 vssd1 vccd1 vccd1 _5384_/A sky130_fd_sc_hd__mux2_1
XANTENNA__5704__A1 _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5619_ _5694_/A _5618_/X _4895_/Y vssd1 vssd1 vccd1 vccd1 _5619_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__3191__A1 _3302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4656__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5341__A _5341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6063__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout81 _3593_/X vssd1 vssd1 vccd1 vccd1 _5179_/S sky130_fd_sc_hd__buf_6
Xfanout70 _3793_/D vssd1 vssd1 vccd1 vccd1 _3724_/S sky130_fd_sc_hd__buf_4
Xfanout92 _5007_/A vssd1 vssd1 vccd1 vccd1 _4990_/A sky130_fd_sc_hd__buf_4
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5156__C1 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3706__A0 _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5171__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4131__B1 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4566__S _4596_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5970_ _6033_/CLK _5970_/D vssd1 vssd1 vccd1 vccd1 _5970_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4434__A1 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4434__B2 _4043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4921_ _4824_/B _4919_/X _4920_/Y _4916_/X vssd1 vssd1 vccd1 vccd1 _4921_/X sky130_fd_sc_hd__a31o_1
XANTENNA__6177__SET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4852_ _6193_/Q _6059_/Q _5216_/A vssd1 vssd1 vccd1 vccd1 _4852_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3803_ _4223_/A _5052_/C vssd1 vssd1 vccd1 vccd1 _3803_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4783_ _6188_/Q _4767_/X _4780_/X _4782_/X vssd1 vssd1 vccd1 vccd1 _4783_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5823__A1_N _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3734_ _5249_/A _3733_/B _4223_/A vssd1 vssd1 vccd1 vccd1 _3734_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3665_ _4223_/A _3664_/X _3573_/B vssd1 vssd1 vccd1 vccd1 _3665_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5404_ _5404_/A _5404_/B vssd1 vssd1 vccd1 vccd1 _5405_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout109_A _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3596_ _4124_/B _3513_/A _3567_/Y vssd1 vssd1 vccd1 vccd1 _3598_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__5860__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5335_ _3654_/S _5046_/A _4022_/X vssd1 vssd1 vccd1 vccd1 _5335_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_2_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5266_ _6206_/Q _5251_/Y _5252_/Y _6214_/Q _5265_/X vssd1 vssd1 vccd1 vccd1 _5266_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4217_ _4217_/A _4217_/B vssd1 vssd1 vccd1 vccd1 _4219_/B sky130_fd_sc_hd__or2_2
XANTENNA__3476__A2 _5424_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5197_ _5898_/Q _3591_/A _3740_/S _6010_/Q _5179_/S vssd1 vssd1 vccd1 vccd1 _5198_/B
+ sky130_fd_sc_hd__o221a_1
X_4148_ _4223_/A _5054_/B _3665_/Y vssd1 vssd1 vccd1 vccd1 _4148_/Y sky130_fd_sc_hd__o21ai_1
X_4079_ _4439_/B _3193_/X _3448_/Y _4124_/B vssd1 vssd1 vccd1 vccd1 _4079_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_78_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3164__A1 _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4587__S1 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5861__A0 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6244__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5010__S _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4415__A _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4719__A2 _4612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3450_ _4726_/A _4618_/C _3443_/X _3449_/X vssd1 vssd1 vccd1 vccd1 _3450_/X sky130_fd_sc_hd__a211o_1
X_3381_ _4474_/A _4457_/A _5872_/A vssd1 vssd1 vccd1 vccd1 _3381_/Y sky130_fd_sc_hd__a21oi_1
X_5120_ _5120_/A _5185_/S vssd1 vssd1 vccd1 vccd1 _5121_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5051_ _5051_/A _5051_/B vssd1 vssd1 vccd1 vccd1 _5051_/X sky130_fd_sc_hd__or2_1
XANTENNA__4296__S _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5852__A0 _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4002_ _3639_/X _3999_/X _4001_/B _4001_/Y _5024_/B vssd1 vssd1 vccd1 vccd1 _4002_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3458__A2 _5424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3213__B _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4407__A1 _5502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5953_ _6123_/CLK _5953_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _5953_/Q sky130_fd_sc_hd__dfstp_1
X_4904_ _4999_/A1 _4899_/X _4903_/X _4824_/B vssd1 vssd1 vccd1 vccd1 _4904_/X sky130_fd_sc_hd__a22o_1
X_5884_ input5/X _5890_/B vssd1 vssd1 vccd1 vccd1 _5884_/X sky130_fd_sc_hd__and2_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4835_ hold351/X _4834_/X _4927_/S vssd1 vssd1 vccd1 vccd1 _4835_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4766_ _4771_/B _4770_/C vssd1 vssd1 vccd1 vccd1 _4766_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__3394__A1 _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3472__A2_N _3370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3717_ _4618_/B _3714_/X _3716_/X _3712_/Y vssd1 vssd1 vccd1 vccd1 _3717_/X sky130_fd_sc_hd__a31o_2
X_4697_ _4696_/X _4695_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4990_/B sky130_fd_sc_hd__mux2_2
X_3648_ _3648_/A vssd1 vssd1 vccd1 vccd1 _3648_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3579_ _3573_/X _3577_/X _3574_/Y vssd1 vssd1 vccd1 vccd1 _3579_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_101_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5318_ _6162_/Q _5320_/S _5317_/Y hold280/X vssd1 vssd1 vccd1 vccd1 _5318_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4894__A1 _4893_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
X_6298_ _6299_/A vssd1 vssd1 vccd1 vccd1 _6298_/X sky130_fd_sc_hd__buf_1
XANTENNA__5843__A0 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5249_ _5249_/A _5259_/B vssd1 vssd1 vccd1 vccd1 _5249_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_2_wb_clk_i _5978_/CLK vssd1 vssd1 vccd1 vccd1 _6006_/CLK sky130_fd_sc_hd__clkbuf_16
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3449__A2 _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4934__S _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xci2406_z80_203 vssd1 vssd1 vccd1 vccd1 ci2406_z80_203/HI io_oeb[18] sky130_fd_sc_hd__conb_1
Xci2406_z80_214 vssd1 vssd1 vccd1 vccd1 io_oeb[33] ci2406_z80_214/LO sky130_fd_sc_hd__conb_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2950_ _3050_/C vssd1 vssd1 vccd1 vccd1 _2950_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4620_ _4617_/X _4618_/X _4497_/S vssd1 vssd1 vccd1 vccd1 _4620_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_17_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4551_ _4549_/X _4550_/X _5872_/A vssd1 vssd1 vccd1 vccd1 _4551_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4482_ _6154_/Q _4481_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4482_/X sky130_fd_sc_hd__mux2_1
Xhold527 _6054_/Q vssd1 vssd1 vccd1 vccd1 hold527/X sky130_fd_sc_hd__buf_1
Xhold505 _3506_/X vssd1 vssd1 vccd1 vccd1 _6153_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold516 _6075_/Q vssd1 vssd1 vccd1 vccd1 _5225_/B sky130_fd_sc_hd__buf_1
X_3502_ _3502_/A _3502_/B vssd1 vssd1 vccd1 vccd1 _5218_/B sky130_fd_sc_hd__nor2_1
X_6221_ _6242_/CLK _6221_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6221_/Q sky130_fd_sc_hd__dfstp_1
Xhold538 _6213_/Q vssd1 vssd1 vccd1 vccd1 hold538/X sky130_fd_sc_hd__dlygate4sd3_1
X_3433_ _4474_/A _5875_/A _5341_/A vssd1 vssd1 vccd1 vccd1 _3433_/X sky130_fd_sc_hd__and3_1
Xhold549 _4506_/X vssd1 vssd1 vccd1 vccd1 _6055_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4876__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6152_ _6152_/CLK hold77/X vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__dfxtp_1
X_5103_ _5120_/A _5105_/B vssd1 vssd1 vccd1 vccd1 _5108_/A sky130_fd_sc_hd__nand2_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ _5566_/S _3364_/B vssd1 vssd1 vccd1 vccd1 _3364_/Y sky130_fd_sc_hd__nor2_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _6127_/Q hold50/A vssd1 vssd1 vccd1 vccd1 _4759_/B sky130_fd_sc_hd__and2b_2
X_6083_ _6086_/CLK _6083_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6083_/Q sky130_fd_sc_hd__dfrtp_1
X_5034_ _6135_/Q _5034_/B _5034_/C _5383_/B vssd1 vssd1 vccd1 vccd1 _5034_/X sky130_fd_sc_hd__or4b_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4039__B _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout176_A input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5936_ _6144_/CLK _5936_/D vssd1 vssd1 vccd1 vccd1 _5936_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__4800__A1 _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5867_ hold375/X _5836_/A _5866_/X _5245_/A vssd1 vssd1 vccd1 vccd1 _5867_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5798_ _6237_/Q _5352_/A _5457_/A hold492/X vssd1 vssd1 vccd1 vccd1 _5798_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__4564__A0 _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4451__A_N _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4818_ _4119_/B _4817_/X _4805_/Y vssd1 vssd1 vccd1 vccd1 _4818_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4749_ _4749_/A _4749_/B _4749_/C vssd1 vssd1 vccd1 vccd1 _4749_/X sky130_fd_sc_hd__or3_1
XFILLER_0_101_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput14 _6293_/X vssd1 vssd1 vccd1 vccd1 io_oeb[24] sky130_fd_sc_hd__buf_12
XFILLER_0_31_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput25 _6082_/Q vssd1 vssd1 vccd1 vccd1 io_out[12] sky130_fd_sc_hd__buf_12
Xoutput36 _6092_/Q vssd1 vssd1 vccd1 vccd1 io_out[22] sky130_fd_sc_hd__buf_12
Xoutput47 _5954_/Q vssd1 vssd1 vccd1 vccd1 io_out[3] sky130_fd_sc_hd__buf_12
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold388_A _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4619__A1 _4617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3134__A _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2973__A _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4095__A2 _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5495__S _5497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3309__A _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4858__B2 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4858__A1 _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3080_ _3131_/B _3079_/X _3077_/X vssd1 vssd1 vccd1 vccd1 _3085_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__5283__A1 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4086__A2 _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3833__A2 _3832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3982_ _5899_/Q _6011_/Q _3982_/S vssd1 vssd1 vccd1 vccd1 _3982_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5721_ hold506/X _5714_/Y _5720_/X _5023_/A vssd1 vssd1 vccd1 vccd1 _5721_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3210__C _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5652_ _5694_/A _5651_/X _4943_/Y vssd1 vssd1 vccd1 vccd1 _5652_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_72_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5418__B _6158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4603_ _6212_/Q _4895_/B _4714_/S vssd1 vssd1 vccd1 vccd1 _4605_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_72_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5583_ _5584_/A _5584_/B _5582_/Y vssd1 vssd1 vccd1 vccd1 _5592_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4534_ hold540/X input4/X _4596_/S vssd1 vssd1 vccd1 vccd1 _4534_/X sky130_fd_sc_hd__mux2_1
Xhold302 _6048_/Q vssd1 vssd1 vccd1 vccd1 _3252_/B sky130_fd_sc_hd__clkbuf_2
Xhold324 _5863_/X vssd1 vssd1 vccd1 vccd1 _6249_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 _5859_/X vssd1 vssd1 vccd1 vccd1 _6248_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold313 _6085_/Q vssd1 vssd1 vccd1 vccd1 hold313/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold346 _5006_/X vssd1 vssd1 vccd1 vccd1 _6092_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 _6087_/Q vssd1 vssd1 vccd1 vccd1 hold357/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4849__A1 _4848_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4465_ _4398_/B _4618_/B _4464_/Y _4463_/X _4460_/A vssd1 vssd1 vccd1 vccd1 _4466_/B
+ sky130_fd_sc_hd__a32o_2
Xhold368 _4106_/X vssd1 vssd1 vccd1 vccd1 _5905_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6204_ _6208_/CLK _6204_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6204_/Q sky130_fd_sc_hd__dfstp_2
Xhold379 _3425_/X vssd1 vssd1 vccd1 vccd1 _5901_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3416_ hold126/X _3415_/X _5875_/A vssd1 vssd1 vccd1 vccd1 _3416_/X sky130_fd_sc_hd__mux2_1
X_4396_ _3426_/A _3276_/A _4618_/C _4728_/B vssd1 vssd1 vccd1 vccd1 _4396_/X sky130_fd_sc_hd__a22o_1
X_6135_ _6175_/CLK _6135_/D vssd1 vssd1 vccd1 vccd1 _6135_/Q sky130_fd_sc_hd__dfxtp_4
X_3347_ _5566_/S vssd1 vssd1 vccd1 vccd1 _5317_/A sky130_fd_sc_hd__inv_6
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ _6219_/CLK _6066_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6066_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _6069_/Q _5702_/A2 _5607_/B1 _5016_/X vssd1 vssd1 vccd1 vccd1 _5017_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3889__A _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3278_ _4726_/C _4614_/B _3434_/B _4615_/B vssd1 vssd1 vccd1 vccd1 _3279_/C sky130_fd_sc_hd__or4_1
XFILLER_0_95_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5919_ _6190_/CLK hold93/X fanout172/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__4785__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5329__A2 _3496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2968__A _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5265__A1 _6156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5265__B2 _6238_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3815__A2 _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4240__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3738__S _4035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5254__A _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4569__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4250_ _4250_/A _4250_/B vssd1 vssd1 vccd1 vccd1 _4251_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4181_ hold143/X _4180_/X _4262_/S vssd1 vssd1 vccd1 vccd1 _4181_/X sky130_fd_sc_hd__mux2_1
X_3201_ _3715_/B _4398_/C _3249_/B _3249_/A _3022_/B vssd1 vssd1 vccd1 vccd1 _3201_/X
+ sky130_fd_sc_hd__o221a_1
X_3132_ _3694_/C _5502_/B vssd1 vssd1 vccd1 vccd1 _4772_/B sky130_fd_sc_hd__and2_1
X_3063_ _3210_/A _3203_/B _4485_/A vssd1 vssd1 vccd1 vccd1 _3063_/X sky130_fd_sc_hd__and3_1
XFILLER_0_77_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3965_ _6151_/Q _3724_/S _3964_/X _3983_/S vssd1 vssd1 vccd1 vccd1 _3968_/B sky130_fd_sc_hd__a211o_1
X_5704_ _5703_/X _6161_/Q _5704_/S vssd1 vssd1 vccd1 vccd1 _5704_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3896_ _3897_/B _3897_/C _6140_/Q vssd1 vssd1 vccd1 vccd1 _3898_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5635_ _5626_/A _5625_/Y _5634_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _5635_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold110 _5944_/Q vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5731__A2 _4850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5566_ _5565_/X hold431/X _5566_/S vssd1 vssd1 vccd1 vccd1 _5566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5497_ _6243_/Q hold361/X _5497_/S vssd1 vssd1 vccd1 vccd1 _5497_/X sky130_fd_sc_hd__mux2_1
Xhold143 _5922_/Q vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold121 _4112_/X vssd1 vssd1 vccd1 vccd1 _5910_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4517_ hold542/X _4612_/B _4516_/Y _4474_/X vssd1 vssd1 vccd1 vccd1 _4517_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_13_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold132 _6146_/Q vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 _4269_/X vssd1 vssd1 vccd1 vccd1 _5933_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold154 _4271_/X vssd1 vssd1 vccd1 vccd1 _5935_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 _6040_/Q vssd1 vssd1 vccd1 vccd1 _3527_/A sky130_fd_sc_hd__dlygate4sd3_1
X_4448_ _4737_/A _3469_/Y _4749_/C _4447_/X _4618_/B vssd1 vssd1 vccd1 vccd1 _4448_/X
+ sky130_fd_sc_hd__o311a_1
Xhold198 _4323_/X vssd1 vssd1 vccd1 vccd1 _5991_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _5962_/Q vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4379_ _4485_/A _3050_/C _3113_/B _4117_/B vssd1 vssd1 vccd1 vccd1 _4379_/X sky130_fd_sc_hd__a31o_1
X_6118_ _6178_/CLK _6118_/D vssd1 vssd1 vccd1 vccd1 _6118_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ _6123_/CLK _6049_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6049_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3412__A _5502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4942__S _5020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5339__A _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4930__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5486__A1 _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5238__A1 _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5013__S _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4852__S _5216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4213__A2 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5249__A _5249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3750_ _3616_/B _3749_/X _3968_/A vssd1 vssd1 vccd1 vccd1 _3750_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3681_ _3683_/B _3683_/C _6136_/Q vssd1 vssd1 vccd1 vccd1 _3684_/A sky130_fd_sc_hd__o21ai_1
X_5420_ _5474_/C _5420_/B vssd1 vssd1 vccd1 vccd1 _5422_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5351_ _5502_/A _5566_/S _5338_/Y _3921_/A vssd1 vssd1 vccd1 vccd1 _5352_/A sky130_fd_sc_hd__or4bb_4
XANTENNA__4299__S _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5282_ _5248_/Y _5279_/X _5281_/X vssd1 vssd1 vccd1 vccd1 _5282_/X sky130_fd_sc_hd__a21o_1
X_4302_ _4150_/X hold145/X _4309_/S vssd1 vssd1 vccd1 vccd1 _4302_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4233_ _4234_/B vssd1 vssd1 vccd1 vccd1 _4233_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3931__S _4035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4164_ hold238/X hold78/X hold201/X hold62/X _5182_/S _5200_/B1 vssd1 vssd1 vccd1
+ vccd1 _4164_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4095_ _4735_/A _4038_/A _3302_/A vssd1 vssd1 vccd1 vccd1 _4095_/X sky130_fd_sc_hd__a21o_1
X_3115_ _3777_/A _5356_/A _3643_/A vssd1 vssd1 vccd1 vccd1 _3116_/B sky130_fd_sc_hd__nand3_1
X_3046_ _4486_/A _4051_/B vssd1 vssd1 vccd1 vccd1 _3184_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_77_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4997_ _5012_/B _4997_/B vssd1 vssd1 vccd1 vccd1 _4997_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_58_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3948_ _4012_/B _3948_/B vssd1 vssd1 vccd1 vccd1 _3948_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_18_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3879_ hold96/X hold120/X hold205/X hold60/X _5182_/S _5200_/B1 vssd1 vssd1 vccd1
+ vccd1 _3879_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5618_ _6062_/Q _5702_/A2 _5702_/B1 _5617_/X vssd1 vssd1 vccd1 vccd1 _5618_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_5_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5549_ _6157_/Q _5507_/Y _5508_/X vssd1 vssd1 vccd1 vccd1 _5551_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3191__A2 _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout71_A _3795_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold635_A _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2981__A _6176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3954__A1 _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout82 _3739_/S vssd1 vssd1 vccd1 vccd1 _3740_/S sky130_fd_sc_hd__clkbuf_8
Xfanout71 _3795_/C vssd1 vssd1 vccd1 vccd1 _3983_/S sky130_fd_sc_hd__clkbuf_8
Xfanout60 _4763_/Y vssd1 vssd1 vccd1 vccd1 _5607_/B1 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3954__B2 _6119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5156__B1 _3739_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4903__A0 _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4131__A1 _3671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_26_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6178_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4434__A2 _3713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4920_ _4948_/C _4918_/Y _5013_/S vssd1 vssd1 vccd1 vccd1 _4920_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4582__S _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4851_ _6059_/Q _4764_/X _4763_/B vssd1 vssd1 vccd1 vccd1 _4851_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_51_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3802_ _3802_/A _3802_/B vssd1 vssd1 vccd1 vccd1 _5052_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4782_ _6154_/Q _5008_/B _4824_/B _4777_/X _4781_/X vssd1 vssd1 vccd1 vccd1 _4782_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3733_ _5249_/A _3733_/B vssd1 vssd1 vccd1 vccd1 _5052_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_82_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3664_ _3663_/X hold363/X _3958_/S vssd1 vssd1 vccd1 vccd1 _3664_/X sky130_fd_sc_hd__mux2_4
XANTENNA__5426__B _5426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5403_ _5403_/A _5403_/B vssd1 vssd1 vccd1 vccd1 _5405_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3227__A _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3595_ hold189/X hold217/X hold86/X hold84/X _3740_/S _5179_/S vssd1 vssd1 vccd1
+ vccd1 _3595_/X sky130_fd_sc_hd__mux4_1
X_5334_ _5332_/B _5333_/Y _5332_/Y vssd1 vssd1 vccd1 vccd1 _5334_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_11_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5265_ _6156_/Q _5253_/Y _5254_/Y _6238_/Q vssd1 vssd1 vccd1 vccd1 _5265_/X sky130_fd_sc_hd__a22o_1
X_4216_ _5950_/Q _3605_/X _3615_/X _6033_/Q _4215_/X vssd1 vssd1 vccd1 vccd1 _4217_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5196_ _6002_/Q _3591_/A _3740_/S _5963_/Q _4256_/S vssd1 vssd1 vccd1 vccd1 _5198_/A
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5870__A1 _4030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4147_ _4147_/A _4147_/B vssd1 vssd1 vccd1 vccd1 _5054_/B sky130_fd_sc_hd__or2_1
XANTENNA__4425__A2 _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5083__C1 _5220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4078_ _3446_/A _3496_/C _4045_/X vssd1 vssd1 vccd1 vccd1 _4416_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3029_ _3193_/A _4417_/A vssd1 vssd1 vccd1 vccd1 _3070_/A sky130_fd_sc_hd__or2_2
XFILLER_0_93_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4667__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2976__A _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5310__A0 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5352__A _5352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4664__A2 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3600__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3927__A1 _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5246__B _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3380_ _4486_/B _3392_/A vssd1 vssd1 vccd1 vccd1 _4457_/A sky130_fd_sc_hd__and2b_1
X_5050_ _5052_/D _5050_/B vssd1 vssd1 vccd1 vccd1 _5051_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_20_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5852__A1 _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4001_ _5024_/A _4001_/B vssd1 vssd1 vccd1 vccd1 _4001_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3312__C1 _6130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5952_ _6035_/CLK _5952_/D vssd1 vssd1 vccd1 vccd1 _5952_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4407__A2 _4391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4903_ _6154_/Q _4902_/Y _5013_/S vssd1 vssd1 vccd1 vccd1 _4903_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4812__C1 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_46_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5883_ _3050_/C _5875_/X _5876_/Y _5882_/X vssd1 vssd1 vccd1 vccd1 _5883_/X sky130_fd_sc_hd__o22a_1
X_4834_ _4833_/X _6057_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3379__C1 _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4765_ _4765_/A _6050_/Q _6036_/Q vssd1 vssd1 vccd1 vccd1 _4765_/Y sky130_fd_sc_hd__nand3_2
XANTENNA_fanout121_A _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3394__A2 _5093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3716_ _4737_/A _4043_/C _4124_/B vssd1 vssd1 vccd1 vccd1 _3716_/X sky130_fd_sc_hd__a21o_1
X_4696_ _6026_/Q _5971_/Q _6018_/Q _5951_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4696_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_70_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3647_ _6073_/Q _3647_/B _3647_/C vssd1 vssd1 vccd1 vccd1 _3648_/A sky130_fd_sc_hd__and3_2
XFILLER_0_11_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3578_ _3573_/X _3577_/X _3574_/Y vssd1 vssd1 vccd1 vccd1 _3968_/A sky130_fd_sc_hd__o21a_4
X_5317_ _5317_/A _5320_/S vssd1 vssd1 vccd1 vccd1 _5317_/Y sky130_fd_sc_hd__nor2_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
X_6297_ _6299_/A vssd1 vssd1 vccd1 vccd1 _6297_/X sky130_fd_sc_hd__buf_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5843__A1 _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5248_ _5250_/A _5250_/B _4409_/X vssd1 vssd1 vccd1 vccd1 _5248_/Y sky130_fd_sc_hd__a21oi_4
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
X_5179_ _6001_/Q _5897_/Q _5179_/S vssd1 vssd1 vccd1 vccd1 _5179_/X sky130_fd_sc_hd__mux2_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3420__A _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3793__C _3795_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xci2406_z80_204 vssd1 vssd1 vccd1 vccd1 ci2406_z80_204/HI io_oeb[19] sky130_fd_sc_hd__conb_1
Xci2406_z80_215 vssd1 vssd1 vccd1 vccd1 io_oeb[34] ci2406_z80_215/LO sky130_fd_sc_hd__conb_1
XFILLER_0_57_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4550_ hold546/X input5/X _4596_/S vssd1 vssd1 vccd1 vccd1 _4550_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold506 _6205_/Q vssd1 vssd1 vccd1 vccd1 hold506/X sky130_fd_sc_hd__buf_1
XFILLER_0_52_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4481_ _4473_/Y _4611_/A _4480_/X _5872_/A vssd1 vssd1 vccd1 vccd1 _4481_/X sky130_fd_sc_hd__a22o_1
Xhold517 _5225_/X vssd1 vssd1 vccd1 vccd1 hold517/X sky130_fd_sc_hd__dlygate4sd3_1
X_3501_ _4038_/A _4118_/A _6094_/Q _3334_/B _4762_/B vssd1 vssd1 vccd1 vccd1 _3502_/B
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_40_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6220_ _6243_/CLK _6220_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6220_/Q sky130_fd_sc_hd__dfstp_1
Xhold539 _5748_/X vssd1 vssd1 vccd1 vccd1 _6213_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold528 _4491_/X vssd1 vssd1 vccd1 vccd1 _6054_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3432_ hold92/X _4457_/B vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__and2_1
XFILLER_0_40_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _5216_/A _3363_/B _3363_/C _3370_/B vssd1 vssd1 vccd1 vccd1 _3364_/B sky130_fd_sc_hd__or4b_1
X_6151_ _6151_/CLK _6151_/D vssd1 vssd1 vccd1 vccd1 _6151_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_41_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6086_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5185_/S vssd1 vssd1 vccd1 vccd1 _5105_/B sky130_fd_sc_hd__inv_2
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _3294_/A _3294_/B _3294_/C vssd1 vssd1 vccd1 vccd1 _3294_/X sky130_fd_sc_hd__or3_1
X_6082_ _6086_/CLK _6082_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6082_/Q sky130_fd_sc_hd__dfrtp_1
X_5033_ _5033_/A _5387_/A _5387_/B vssd1 vssd1 vccd1 vccd1 _5034_/C sky130_fd_sc_hd__or3b_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_A _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5935_ _6111_/CLK _5935_/D vssd1 vssd1 vccd1 vccd1 _5935_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5866_ _3959_/Y _5834_/X _5837_/X _5865_/X vssd1 vssd1 vccd1 vccd1 _5866_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3894__B _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4817_ _4816_/X _6056_/Q _5595_/S vssd1 vssd1 vccd1 vccd1 _4817_/X sky130_fd_sc_hd__mux2_1
X_5797_ hold598/X _5796_/X _5832_/S vssd1 vssd1 vccd1 vccd1 _6236_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_16_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4748_ _5164_/A1 hold614/X _4927_/S _4747_/Y vssd1 vssd1 vccd1 vccd1 _4748_/X sky130_fd_sc_hd__a22o_1
X_4679_ hold501/X _5762_/A _4619_/X vssd1 vssd1 vccd1 vccd1 _4679_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_31_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput15 _6294_/X vssd1 vssd1 vccd1 vccd1 io_oeb[25] sky130_fd_sc_hd__buf_12
XFILLER_0_101_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput37 _6093_/Q vssd1 vssd1 vccd1 vccd1 io_out[23] sky130_fd_sc_hd__buf_12
Xoutput48 _5955_/Q vssd1 vssd1 vccd1 vccd1 io_out[4] sky130_fd_sc_hd__buf_12
Xoutput26 _6083_/Q vssd1 vssd1 vccd1 vccd1 io_out[13] sky130_fd_sc_hd__buf_12
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5816__A1 _3864_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5052__D _5052_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5504__B1 _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4858__A2 _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3981_ hold76/A hold58/A _3982_/S vssd1 vssd1 vccd1 vccd1 _3981_/X sky130_fd_sc_hd__mux2_1
X_5720_ _3707_/X _5715_/B _5715_/Y _5719_/X vssd1 vssd1 vccd1 vccd1 _5720_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3995__A _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5651_ _6065_/Q _5702_/A2 _5702_/B1 _5650_/X vssd1 vssd1 vccd1 vccd1 _5651_/X sky130_fd_sc_hd__a22o_1
X_4602_ _4601_/X _4600_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4895_/B sky130_fd_sc_hd__mux2_2
X_5582_ _5582_/A _5582_/B vssd1 vssd1 vccd1 vccd1 _5582_/Y sky130_fd_sc_hd__xnor2_1
X_4533_ _4531_/Y _4532_/X _4565_/S vssd1 vssd1 vccd1 vccd1 _4533_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold325 hold661/X vssd1 vssd1 vccd1 vccd1 _5790_/D sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5715__A _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold314 _4894_/X vssd1 vssd1 vccd1 vccd1 _6085_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold303 _5243_/X vssd1 vssd1 vccd1 vccd1 _6133_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6203_ _6203_/CLK _6203_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6203_/Q sky130_fd_sc_hd__dfrtp_2
Xhold358 _4927_/X vssd1 vssd1 vccd1 vccd1 _6087_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold336 _6244_/Q vssd1 vssd1 vccd1 vccd1 hold336/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4464_ _3302_/A _3554_/A _3439_/B vssd1 vssd1 vccd1 vccd1 _4464_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold369 _5917_/Q vssd1 vssd1 vccd1 vccd1 _3389_/B sky130_fd_sc_hd__dlygate4sd3_1
Xhold347 _6083_/Q vssd1 vssd1 vccd1 vccd1 hold347/X sky130_fd_sc_hd__dlygate4sd3_1
X_4395_ _5289_/S vssd1 vssd1 vccd1 vccd1 _5259_/B sky130_fd_sc_hd__inv_2
X_3415_ _5918_/Q _3210_/C _4070_/B _3413_/X _3414_/Y vssd1 vssd1 vccd1 vccd1 _3415_/X
+ sky130_fd_sc_hd__a311o_1
X_6134_ _6227_/CLK _6134_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6134_/Q sky130_fd_sc_hd__dfrtp_1
X_3346_ _6162_/Q _3343_/A _3340_/X _5319_/B vssd1 vssd1 vccd1 vccd1 _3346_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ _6219_/CLK _6065_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6065_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _6187_/Q _5015_/X _5701_/S vssd1 vssd1 vccd1 vccd1 _5016_/X sky130_fd_sc_hd__mux2_1
X_3277_ _3277_/A _4439_/A vssd1 vssd1 vccd1 vccd1 _4483_/B sky130_fd_sc_hd__or2_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4482__A0 _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5918_ _6038_/CLK _5918_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _5918_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5849_ _6115_/Q _5848_/X _5869_/S vssd1 vssd1 vccd1 vccd1 _5849_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3844__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5501__A3 _4043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__2984__A _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6057__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4068__A3 _4043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5360__A _5360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3815__A3 _6116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5017__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4528__A1 _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4180_ _4242_/S _4179_/X _4178_/X vssd1 vssd1 vccd1 vccd1 _4180_/X sky130_fd_sc_hd__a21o_2
X_3200_ _3200_/A _3200_/B _3200_/C vssd1 vssd1 vccd1 vccd1 _3200_/X sky130_fd_sc_hd__and3_1
X_3131_ _3249_/A _3131_/B vssd1 vssd1 vccd1 vccd1 _5502_/D sky130_fd_sc_hd__nor2_2
XFILLER_0_89_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3062_ _3507_/C _3507_/D vssd1 vssd1 vccd1 vccd1 _4726_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_89_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4216__B1 _3615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4614__A _5502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3964_ _3573_/C _3986_/A2 _3584_/X _3585_/X _5912_/Q vssd1 vssd1 vccd1 vccd1 _3964_/X
+ sky130_fd_sc_hd__o311a_1
X_5703_ _5694_/A _5702_/X _5007_/Y vssd1 vssd1 vccd1 vccd1 _5703_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_72_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3895_ _5024_/A _6118_/Q vssd1 vssd1 vccd1 vccd1 _3897_/C sky130_fd_sc_hd__and2_1
X_5634_ _5670_/A _5628_/Y _5629_/Y _5633_/X vssd1 vssd1 vccd1 vccd1 _5634_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5192__A1 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3727__C1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold100 _5967_/Q vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5565_ _5564_/X _6058_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _5565_/X sky130_fd_sc_hd__mux2_1
X_5496_ _6242_/Q hold332/X _5497_/S vssd1 vssd1 vccd1 vccd1 _5496_/X sky130_fd_sc_hd__mux2_1
Xhold111 _4282_/X vssd1 vssd1 vccd1 vccd1 _5944_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 _4181_/X vssd1 vssd1 vccd1 vccd1 _5922_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 _6026_/Q vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 _6028_/Q vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ _4516_/A _4516_/B vssd1 vssd1 vccd1 vccd1 _4516_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__3742__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold166 _5950_/Q vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 _5920_/Q vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold155 _5896_/Q vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
X_4447_ _3446_/A _3097_/Y _3264_/B _4444_/X _4445_/Y vssd1 vssd1 vccd1 vccd1 _4447_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold199 _6008_/Q vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 _4298_/X vssd1 vssd1 vccd1 vccd1 _5962_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6117_ _6119_/CLK _6117_/D vssd1 vssd1 vccd1 vccd1 _6117_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4378_ hold52/X _4377_/Y _4927_/S vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__mux2_1
X_3329_ _3715_/B _5498_/B vssd1 vssd1 vccd1 vccd1 _3329_/Y sky130_fd_sc_hd__nand2_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4455__B1 _5314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6048_ _6123_/CLK _6048_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6048_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4758__A1 _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5339__B wire93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5183__B2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3680_ _5333_/B _6114_/Q vssd1 vssd1 vccd1 vccd1 _3683_/C sky130_fd_sc_hd__and2b_1
XANTENNA__4921__A1 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5350_ hold649/X _5349_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _5350_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5281_ _6209_/Q _5251_/Y _5252_/Y _6217_/Q _5280_/X vssd1 vssd1 vccd1 vccd1 _5281_/X
+ sky130_fd_sc_hd__a221o_1
X_4301_ _4319_/B _4364_/B vssd1 vssd1 vccd1 vccd1 _4309_/S sky130_fd_sc_hd__or2_4
XFILLER_0_50_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4232_ _4232_/A _4232_/B vssd1 vssd1 vccd1 vccd1 _4234_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4163_ hold36/X _3539_/Y _3708_/X _4162_/Y _3671_/B vssd1 vssd1 vccd1 vccd1 _4163_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3513__A _3513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4094_ _3113_/B _4094_/B _4094_/C _4094_/D vssd1 vssd1 vccd1 vccd1 _4094_/X sky130_fd_sc_hd__and4b_1
X_3114_ _3777_/A _5356_/A _3193_/A vssd1 vssd1 vccd1 vccd1 _4021_/B sky130_fd_sc_hd__and3_2
XANTENNA__4988__A1 _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3232__B _5424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3045_ _4051_/B _3249_/B vssd1 vssd1 vccd1 vccd1 _3324_/A sky130_fd_sc_hd__or2_1
XANTENNA__3660__A1 _6135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4996_ _6067_/Q _4995_/C _6068_/Q vssd1 vssd1 vccd1 vccd1 _4997_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3947_ _4014_/A _4012_/A vssd1 vssd1 vccd1 vccd1 _3948_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3878_ hold13/X _4253_/A2 _3865_/Y _3877_/Y vssd1 vssd1 vccd1 vccd1 _3878_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5617_ _6180_/Q _6196_/Q _5701_/S vssd1 vssd1 vccd1 vccd1 _5617_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5165__B2 _6240_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5548_ _2992_/A _5547_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _5548_/X sky130_fd_sc_hd__mux2_1
X_5479_ _6179_/Q _5372_/B _5479_/S vssd1 vssd1 vccd1 vccd1 _5479_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold363_A _6113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4523__S0 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout64_A _4761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout61 _4763_/Y vssd1 vssd1 vccd1 vccd1 _5702_/B1 sky130_fd_sc_hd__buf_2
Xfanout83 _3739_/S vssd1 vssd1 vccd1 vccd1 _5200_/B1 sky130_fd_sc_hd__buf_4
Xfanout72 _3582_/Y vssd1 vssd1 vccd1 vccd1 _3616_/B sky130_fd_sc_hd__buf_4
XFILLER_0_91_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout94 _4412_/B vssd1 vssd1 vccd1 vccd1 _4070_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__5085__A _5107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5459__A2 _3377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4863__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5092__B1 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5631__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_36_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4850_ _4990_/A _4850_/B vssd1 vssd1 vccd1 vccd1 _4850_/Y sky130_fd_sc_hd__nand2_1
X_3801_ _3759_/A _5052_/B _3756_/Y vssd1 vssd1 vccd1 vccd1 _3802_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4781_ _6204_/Q _4768_/Y _4769_/Y _4779_/B _4815_/B vssd1 vssd1 vccd1 vccd1 _4781_/X
+ sky130_fd_sc_hd__a221o_1
X_3732_ _3730_/X _3732_/B vssd1 vssd1 vccd1 vccd1 _3733_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__5147__A1 _6174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5147__B2 _6156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3663_ _3533_/S _6154_/Q _3662_/X vssd1 vssd1 vccd1 vccd1 _3663_/X sky130_fd_sc_hd__a21o_1
X_5402_ _5480_/S _6174_/Q _5400_/Y _5401_/X vssd1 vssd1 vccd1 vccd1 _5402_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5333_ _6072_/Q _5333_/B vssd1 vssd1 vccd1 vccd1 _5333_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_23_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3594_ _5905_/Q _4034_/S _3592_/Y vssd1 vssd1 vccd1 vccd1 _3594_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_100_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5264_ _3755_/Y _4173_/B _5289_/S vssd1 vssd1 vccd1 vccd1 _5264_/X sky130_fd_sc_hd__mux2_1
X_4215_ _5925_/Q _3588_/X _3603_/X _6017_/Q vssd1 vssd1 vccd1 vccd1 _4215_/X sky130_fd_sc_hd__a22o_1
X_5195_ _6202_/Q _5119_/Y _5121_/Y _6160_/Q vssd1 vssd1 vccd1 vccd1 _5204_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4146_ _4145_/B _4146_/B vssd1 vssd1 vccd1 vccd1 _4147_/B sky130_fd_sc_hd__and2b_1
XANTENNA__5869__S _5869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4077_ _4077_/A _4415_/A vssd1 vssd1 vccd1 vccd1 _4077_/X sky130_fd_sc_hd__or2_2
X_3028_ _3203_/B _4485_/A _3210_/A vssd1 vssd1 vccd1 vccd1 _3249_/A sky130_fd_sc_hd__or3b_4
XANTENNA__4074__A _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4979_ _6201_/Q _6067_/Q _6038_/Q vssd1 vssd1 vccd1 vccd1 _4979_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3397__B1 _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5138__B2 _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5138__A1 _6197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4897__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3872__A1 _3795_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3600__B _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3927__A2 _3926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4000_ _5046_/A _6120_/Q vssd1 vssd1 vccd1 vccd1 _4001_/B sky130_fd_sc_hd__nand2_1
X_5951_ _6032_/CLK _5951_/D vssd1 vssd1 vccd1 vccd1 _5951_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4407__A3 _4043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4902_ _4918_/B _4902_/B vssd1 vssd1 vccd1 vccd1 _4902_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4812__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5882_ input4/X _5890_/B vssd1 vssd1 vccd1 vccd1 _5882_/X sky130_fd_sc_hd__and2_1
XANTENNA__5368__A1 _6174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4833_ _4119_/B _4832_/X _4821_/Y vssd1 vssd1 vccd1 vccd1 _4833_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4764_ _4765_/A _6050_/Q _6036_/Q vssd1 vssd1 vccd1 vccd1 _4764_/X sky130_fd_sc_hd__and3_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3715_ _3777_/A _3715_/B vssd1 vssd1 vccd1 vccd1 _3715_/Y sky130_fd_sc_hd__nor2_1
X_4695_ hold64/A hold80/A _5926_/Q _6034_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4695_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3238__A _3694_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3646_ _6072_/Q _6070_/Q _5024_/A _6073_/Q vssd1 vssd1 vccd1 vccd1 _3646_/X sky130_fd_sc_hd__and4b_4
XFILLER_0_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3672__S _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3577_ hold27/A _6052_/Q _3577_/S vssd1 vssd1 vccd1 vccd1 _3577_/X sky130_fd_sc_hd__mux2_1
X_6296_ _6299_/A vssd1 vssd1 vccd1 vccd1 _6296_/X sky130_fd_sc_hd__buf_1
X_5316_ _5314_/Y _5315_/X _3520_/Y vssd1 vssd1 vccd1 vccd1 _5320_/S sky130_fd_sc_hd__o21ai_4
XFILLER_0_11_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3551__B1 _5424_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5247_ _5250_/A _5250_/B vssd1 vssd1 vccd1 vccd1 _5254_/B sky130_fd_sc_hd__nand2_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5599__S _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5178_ _5962_/Q _6009_/Q _5179_/S vssd1 vssd1 vccd1 vccd1 _5178_/X sky130_fd_sc_hd__mux2_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4129_ _3527_/A _4129_/B vssd1 vssd1 vccd1 vccd1 _5834_/D sky130_fd_sc_hd__nand2b_1
XFILLER_0_97_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3701__A _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3420__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5359__A1 _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2987__A _6158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3611__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5302__S _5305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_205 vssd1 vssd1 vccd1 vccd1 ci2406_z80_205/HI io_oeb[20] sky130_fd_sc_hd__conb_1
Xci2406_z80_216 vssd1 vssd1 vccd1 vccd1 io_oeb[35] ci2406_z80_216/LO sky130_fd_sc_hd__conb_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5770__B2 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3500_ hold50/A _5902_/Q _5903_/Q _4765_/A _3499_/X vssd1 vssd1 vccd1 vccd1 _4762_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3058__A _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold507 _5721_/X vssd1 vssd1 vccd1 vccd1 _6205_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4480_ hold527/X input1/X _4596_/S vssd1 vssd1 vccd1 vccd1 _4480_/X sky130_fd_sc_hd__mux2_1
Xhold518 _5235_/X vssd1 vssd1 vccd1 vccd1 hold518/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4588__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold529 _6050_/Q vssd1 vssd1 vccd1 vccd1 _4478_/A sky130_fd_sc_hd__clkbuf_2
X_3431_ _3193_/C _5489_/D _3421_/Y _3429_/Y hold46/X vssd1 vssd1 vccd1 vccd1 hold47/A
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5522__A1 _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6150_ _6152_/CLK _6150_/D vssd1 vssd1 vccd1 vccd1 _6150_/Q sky130_fd_sc_hd__dfxtp_1
X_3362_ _4077_/A _6047_/Q _4043_/C _3503_/C vssd1 vssd1 vccd1 vccd1 _3363_/C sky130_fd_sc_hd__or4_1
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _3203_/B _5089_/X _5100_/Y _4077_/A vssd1 vssd1 vccd1 vccd1 _5185_/S sky130_fd_sc_hd__o2bb2a_4
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3293_ _3285_/Y _3286_/Y _3290_/X _3715_/B vssd1 vssd1 vccd1 vccd1 _3294_/C sky130_fd_sc_hd__a2bb2o_1
XANTENNA__4089__B2 _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6081_ _6086_/CLK _6081_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6081_/Q sky130_fd_sc_hd__dfrtp_1
X_5032_ _5386_/A _5032_/B vssd1 vssd1 vccd1 vccd1 _5034_/B sky130_fd_sc_hd__nand2_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3836__A1 _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_10_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6149_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3521__A _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3240__B _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5934_ _6032_/CLK hold81/X vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5865_ _6119_/Q _5864_/X _5869_/S vssd1 vssd1 vccd1 vccd1 _5865_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4816_ _5606_/S _4814_/X _4815_/Y _4806_/X vssd1 vssd1 vccd1 vccd1 _4816_/X sky130_fd_sc_hd__a31o_1
X_5796_ _5795_/X _3664_/X _5831_/S vssd1 vssd1 vccd1 vccd1 _5796_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5210__B1 _5105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4747_ _2957_/Y _4431_/X _4746_/X vssd1 vssd1 vccd1 vccd1 _4747_/Y sky130_fd_sc_hd__o21ai_1
X_4678_ hold501/X _4612_/B _4677_/X _4474_/X vssd1 vssd1 vccd1 vccd1 _4678_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3119__A3 _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3629_ _6135_/Q _3629_/B vssd1 vssd1 vccd1 vccd1 _3636_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_101_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput38 _6244_/Q vssd1 vssd1 vccd1 vccd1 io_out[24] sky130_fd_sc_hd__buf_12
Xoutput16 _6295_/X vssd1 vssd1 vccd1 vccd1 io_oeb[26] sky130_fd_sc_hd__buf_12
XANTENNA__3524__B1 _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput49 _5956_/Q vssd1 vssd1 vccd1 vccd1 io_out[5] sky130_fd_sc_hd__buf_12
Xoutput27 _6084_/Q vssd1 vssd1 vccd1 vccd1 io_out[14] sky130_fd_sc_hd__buf_12
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4527__A _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3150__B _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4252__A1 _4239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5752__A1 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5752__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3606__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3980_ hold271/X _3979_/X _4035_/S vssd1 vssd1 vccd1 vccd1 _3980_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5650_ _6183_/Q _6199_/Q _5701_/S vssd1 vssd1 vccd1 vccd1 _5650_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4601_ _6020_/Q _6012_/Q _5965_/Q _5945_/Q _4712_/S1 _4712_/S0 vssd1 vssd1 vccd1
+ vccd1 _4601_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5743__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5743__A1 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5581_ _5582_/A _5582_/B vssd1 vssd1 vccd1 vccd1 _5592_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_53_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4532_ _5868_/S hold540/X _4564_/S vssd1 vssd1 vccd1 vccd1 _4532_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5715__B _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold315 _6245_/Q vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4463_ _3303_/B _3396_/D _4462_/X _4398_/B vssd1 vssd1 vccd1 vccd1 _4463_/X sky130_fd_sc_hd__a22o_1
Xhold326 _5915_/Q vssd1 vssd1 vccd1 vccd1 _5330_/A sky130_fd_sc_hd__buf_1
Xhold304 _6096_/Q vssd1 vssd1 vccd1 vccd1 _2999_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6202_ _6203_/CLK _6202_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6202_/Q sky130_fd_sc_hd__dfrtp_2
Xhold337 _5842_/X vssd1 vssd1 vccd1 vccd1 _6244_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4111__S _4115_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3414_ _4445_/B _3554_/A _5424_/B vssd1 vssd1 vccd1 vccd1 _3414_/Y sky130_fd_sc_hd__a21oi_1
Xhold359 _6052_/Q vssd1 vssd1 vccd1 vccd1 _3272_/A sky130_fd_sc_hd__buf_1
XFILLER_0_40_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold348 _4864_/X vssd1 vssd1 vccd1 vccd1 _6083_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4394_ _3148_/B _2957_/Y _3457_/A _4393_/X _4388_/Y vssd1 vssd1 vccd1 vccd1 _5289_/S
+ sky130_fd_sc_hd__o221a_4
XFILLER_0_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3345_ hold280/X _3341_/Y _3344_/X _3343_/B _3343_/Y vssd1 vssd1 vccd1 vccd1 _5319_/B
+ sky130_fd_sc_hd__a221o_1
X_6133_ _6170_/CLK _6133_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6133_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ _6219_/CLK _6064_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6064_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3276_ _3276_/A _5502_/C _4094_/B _4439_/B vssd1 vssd1 vccd1 vccd1 _4424_/D sky130_fd_sc_hd__or4_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _6203_/Q _4766_/Y _5009_/X _5014_/X vssd1 vssd1 vccd1 vccd1 _5015_/X sky130_fd_sc_hd__a211o_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout181_A fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5917_ _6038_/CLK _5917_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _5917_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5848_ _6119_/Q _6137_/Q _5868_/S vssd1 vssd1 vccd1 vccd1 _5848_/X sky130_fd_sc_hd__mux2_1
X_5779_ _6241_/Q hold476/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5779_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5734__A1 _4116_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5734__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3426__A _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4170__B1 _3615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5360__B _5424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5725__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5725__A1 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3736__B1 _3671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3130_ _3012_/B _3079_/X _3203_/C vssd1 vssd1 vccd1 vccd1 _3140_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__4464__A1 _3302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3061_ _4486_/A _4406_/A vssd1 vssd1 vccd1 vccd1 _3507_/D sky130_fd_sc_hd__or2_2
XANTENNA__3071__A _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5110__C1 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4614__B _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3963_ _3961_/X _3962_/X _3983_/S vssd1 vssd1 vccd1 vccd1 _3963_/X sky130_fd_sc_hd__mux2_1
X_5702_ _6069_/Q _5702_/A2 _5702_/B1 _5701_/X vssd1 vssd1 vccd1 vccd1 _5702_/X sky130_fd_sc_hd__a22o_1
X_3894_ _3894_/A _6118_/Q vssd1 vssd1 vccd1 vccd1 _3897_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5633_ _5632_/X _6155_/Q _5704_/S vssd1 vssd1 vccd1 vccd1 _5633_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5716__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5716__A1 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5564_ _4119_/B _5563_/X _4836_/Y vssd1 vssd1 vccd1 vccd1 _5564_/X sky130_fd_sc_hd__a21bo_1
Xhold101 _4304_/X vssd1 vssd1 vccd1 vccd1 _5967_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5445__B _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4515_ _4501_/A _4500_/B _4498_/X vssd1 vssd1 vccd1 vccd1 _4516_/B sky130_fd_sc_hd__a21o_1
X_5495_ _6241_/Q hold380/X _5497_/S vssd1 vssd1 vccd1 vccd1 _5495_/X sky130_fd_sc_hd__mux2_1
Xhold134 _4362_/X vssd1 vssd1 vccd1 vccd1 _6026_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _4365_/X vssd1 vssd1 vccd1 vccd1 _6028_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 _6148_/Q vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__buf_1
XFILLER_0_41_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold167 _4289_/X vssd1 vssd1 vccd1 vccd1 _5950_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _5965_/Q vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 _3881_/X vssd1 vssd1 vccd1 vccd1 _5896_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ _4446_/A _4446_/B vssd1 vssd1 vccd1 vccd1 _4749_/C sky130_fd_sc_hd__nor2_1
Xhold178 _4151_/X vssd1 vssd1 vccd1 vccd1 _5920_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 _5988_/Q vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
X_4377_ _6095_/Q _4377_/B vssd1 vssd1 vccd1 vccd1 _4377_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_95_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6116_ _6119_/CLK _6116_/D vssd1 vssd1 vccd1 vccd1 _6116_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3328_ _3498_/A _3328_/B vssd1 vssd1 vccd1 vccd1 _3328_/Y sky130_fd_sc_hd__nor2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ _6227_/CLK _6047_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6047_/Q sky130_fd_sc_hd__dfrtp_4
X_3259_ _4124_/A _3540_/A vssd1 vssd1 vccd1 vccd1 _4044_/B sky130_fd_sc_hd__nor2_4
XANTENNA__3258__A2 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4455__A1 _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4077__A _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6190__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4805__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4758__A2 _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4016__S _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5168__C1 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3603__B _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_26_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__5310__S _5313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5159__C1 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3066__A _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4382__B1 _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5280_ _6159_/Q _5253_/Y _5254_/Y _6241_/Q vssd1 vssd1 vccd1 vccd1 _5280_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_49_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4300_ _4034_/X hold241/X _4300_/S vssd1 vssd1 vccd1 vccd1 _5964_/D sky130_fd_sc_hd__mux2_1
X_4231_ _5951_/Q _3605_/X _3615_/X _6034_/Q _4230_/X vssd1 vssd1 vccd1 vccd1 _4232_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4596__S _4596_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4162_ _4223_/A _5054_/C vssd1 vssd1 vccd1 vccd1 _4162_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3513__B _6170_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4437__A1 _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4093_ _3127_/B _4750_/A _4079_/X _4092_/X vssd1 vssd1 vccd1 vccd1 _4099_/B sky130_fd_sc_hd__a211o_1
X_3113_ _4485_/A _3113_/B vssd1 vssd1 vccd1 vccd1 _3192_/B sky130_fd_sc_hd__nand2_8
X_3044_ _4051_/B _3249_/B vssd1 vssd1 vccd1 vccd1 _3172_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4437__B2 _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4995_ _6067_/Q _6068_/Q _4995_/C vssd1 vssd1 vccd1 vccd1 _5012_/B sky130_fd_sc_hd__and3_1
XFILLER_0_81_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3946_ _6141_/Q _4009_/C vssd1 vssd1 vccd1 vccd1 _4012_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_18_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3877_ _4223_/A _5053_/A vssd1 vssd1 vccd1 vccd1 _3877_/Y sky130_fd_sc_hd__nor2_1
X_5616_ _5616_/A _5616_/B vssd1 vssd1 vccd1 vccd1 _5616_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5547_ _5670_/A _5552_/B _5540_/X _5546_/X vssd1 vssd1 vccd1 vccd1 _5547_/X sky130_fd_sc_hd__a31o_1
X_5478_ hold606/X _5477_/Y _5488_/S vssd1 vssd1 vccd1 vccd1 _6178_/D sky130_fd_sc_hd__mux2_1
X_4429_ _5338_/B _4429_/B _5338_/C vssd1 vssd1 vccd1 vccd1 _4429_/X sky130_fd_sc_hd__or3_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5625__B1 _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4523__S1 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout57_A _4766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout62 _5511_/X vssd1 vssd1 vccd1 vccd1 _5670_/A sky130_fd_sc_hd__clkbuf_8
Xfanout73 _4715_/A vssd1 vssd1 vccd1 vccd1 _4699_/A sky130_fd_sc_hd__buf_4
Xfanout84 _3739_/S vssd1 vssd1 vccd1 vccd1 _4255_/S sky130_fd_sc_hd__clkbuf_4
Xfanout95 _4056_/A vssd1 vssd1 vccd1 vccd1 _3210_/C sky130_fd_sc_hd__buf_4
XFILLER_0_101_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5156__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5085__B _5085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5864__A0 _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5305__S _5305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6041__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3642__A2 _6135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3800_ _4234_/A _3800_/B vssd1 vssd1 vccd1 vccd1 _3802_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4780_ _4104_/B _4778_/X _4779_/X _4999_/A1 vssd1 vssd1 vccd1 vccd1 _4780_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3731_ _3730_/B _3730_/C _4234_/A vssd1 vssd1 vccd1 vccd1 _3732_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6233_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3662_ _3623_/X _5374_/A _3660_/X _3661_/X _6074_/Q vssd1 vssd1 vccd1 vccd1 _3662_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5401_ _5400_/A _5400_/B _5507_/A vssd1 vssd1 vccd1 vccd1 _5401_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3679__A_N _6114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3508__B _6121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3593_ _5905_/Q _4034_/S _3592_/Y vssd1 vssd1 vccd1 vccd1 _3593_/X sky130_fd_sc_hd__o21a_1
X_5332_ _5448_/B _5332_/B vssd1 vssd1 vccd1 vccd1 _5332_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5263_ _5773_/A hold522/X _5245_/Y _5262_/X vssd1 vssd1 vccd1 vccd1 _5263_/X sky130_fd_sc_hd__a22o_1
X_4214_ _6025_/Q _3599_/X _3601_/X _5970_/Q _4213_/X vssd1 vssd1 vccd1 vccd1 _4217_/A
+ sky130_fd_sc_hd__a221o_1
X_5194_ _6242_/Q _5108_/Y _5129_/Y _5767_/B vssd1 vssd1 vccd1 vccd1 _5204_/B sky130_fd_sc_hd__a22o_1
X_4145_ _4146_/B _4145_/B vssd1 vssd1 vccd1 vccd1 _4147_/A sky130_fd_sc_hd__and2b_1
XANTENNA__5607__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5083__A1 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4076_ hold27/X _4075_/X _5296_/S vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__mux2_1
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3027_ _3203_/A _3203_/B vssd1 vssd1 vccd1 vccd1 _3113_/B sky130_fd_sc_hd__nor2_4
XANTENNA__4074__B _4104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4978_ _6217_/Q _5009_/A2 _4769_/Y _4976_/B _4977_/X vssd1 vssd1 vccd1 vccd1 _4978_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3929_ hold147/X hold98/X hold104/X hold216/X _5179_/S _3740_/S vssd1 vssd1 vccd1
+ vccd1 _3929_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4897__B2 _4895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4649__B2 _4474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3609__C1 _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4888__A1 _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4888__B2 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3312__A1 _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3312__B2 _5918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5950_ _6033_/CLK _5950_/D vssd1 vssd1 vccd1 vccd1 _5950_/Q sky130_fd_sc_hd__dfxtp_1
X_4901_ _4901_/A _4901_/B vssd1 vssd1 vccd1 vccd1 _4902_/B sky130_fd_sc_hd__and2_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5881_ _4094_/D _5875_/X _5876_/Y _5880_/X vssd1 vssd1 vccd1 vccd1 _5881_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_75_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4832_ _6057_/Q _5595_/S _5607_/B1 _4831_/X vssd1 vssd1 vccd1 vccd1 _4832_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3379__A1 _3434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4763_ _5595_/S _4763_/B vssd1 vssd1 vccd1 vccd1 _4763_/Y sky130_fd_sc_hd__nor2_2
X_4694_ hold510/X _4693_/X _5073_/S vssd1 vssd1 vccd1 vccd1 _4694_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3714_ _3562_/Y _3713_/Y _3090_/Y vssd1 vssd1 vccd1 vccd1 _3714_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4114__S _4115_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3645_ _6070_/Q _3655_/B vssd1 vssd1 vccd1 vccd1 _3645_/X sky130_fd_sc_hd__and2b_4
XFILLER_0_3_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout107_A _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3576_ _3513_/A _3571_/X _3559_/B _3552_/X vssd1 vssd1 vccd1 vccd1 _3577_/S sky130_fd_sc_hd__a211oi_4
X_6295_ _6299_/A vssd1 vssd1 vccd1 vccd1 _6295_/X sky130_fd_sc_hd__buf_1
X_5315_ _3523_/A _3329_/Y _3523_/B _3532_/B _5566_/S vssd1 vssd1 vccd1 vccd1 _5315_/X
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3551__A1 _5424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5246_ _5246_/A _5289_/S vssd1 vssd1 vccd1 vccd1 _5246_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3254__A _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4784__S _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5177_ _5023_/A _2979_/A _5086_/Y _5176_/X vssd1 vssd1 vccd1 vccd1 _5177_/X sky130_fd_sc_hd__a22o_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
X_4128_ _3405_/B _5330_/A _4127_/Y vssd1 vssd1 vccd1 vccd1 _4128_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3701__B _6176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4059_ _3556_/A _4055_/X _4058_/X _3457_/A vssd1 vssd1 vccd1 vccd1 _4059_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_66_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5359__A2 _5341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold590_A _5914_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5363__B _5363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4694__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3611__B _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_206 vssd1 vssd1 vccd1 vccd1 ci2406_z80_206/HI io_oeb[21] sky130_fd_sc_hd__conb_1
Xci2406_z80_217 vssd1 vssd1 vccd1 vccd1 io_out[7] ci2406_z80_217/LO sky130_fd_sc_hd__conb_1
XFILLER_0_69_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3058__B _3694_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold508 _6135_/Q vssd1 vssd1 vccd1 vccd1 hold508/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold519 _5236_/X vssd1 vssd1 vccd1 vccd1 _6129_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3430_ _5489_/D _3427_/X _3429_/Y hold300/X vssd1 vssd1 vccd1 vccd1 _3430_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3533__A1 _5837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3361_ hold56/X _3353_/X _3376_/B vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__a21o_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _4460_/A _5099_/X _5092_/X vssd1 vssd1 vccd1 vccd1 _5100_/Y sky130_fd_sc_hd__a21oi_1
X_6080_ _6170_/CLK _6080_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6080_/Q sky130_fd_sc_hd__dfrtp_1
X_5031_ _2960_/Y _6046_/Q _5030_/X _6073_/Q vssd1 vssd1 vccd1 vccd1 _5031_/X sky130_fd_sc_hd__a211o_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3292_ _3488_/B _3543_/B _3289_/Y _3395_/B _3291_/X vssd1 vssd1 vccd1 vccd1 _3294_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4089__A2 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3297__B1 _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5038__A1 _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3521__B _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4109__S _4115_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5933_ _6035_/CLK _5933_/D vssd1 vssd1 vccd1 vccd1 _5933_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_wb_clk_i _5978_/CLK vssd1 vssd1 vccd1 vccd1 _6129_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5864_ _6137_/Q _6115_/Q _5868_/S vssd1 vssd1 vccd1 vccd1 _5864_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4815_ _5538_/A _4815_/B vssd1 vssd1 vccd1 vccd1 _4815_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5795_ _5794_/B _5793_/X _5794_/Y hold371/X vssd1 vssd1 vccd1 vccd1 _5795_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5210__A1 _5116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3221__B1 _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4746_ _4485_/B _4416_/B _4737_/B _5424_/B vssd1 vssd1 vccd1 vccd1 _4746_/X sky130_fd_sc_hd__o2bb2a_1
X_4677_ _4677_/A _4677_/B vssd1 vssd1 vccd1 vccd1 _4677_/X sky130_fd_sc_hd__xor2_1
X_3628_ _5333_/B _3628_/B vssd1 vssd1 vccd1 vccd1 _3628_/X sky130_fd_sc_hd__or2_1
Xoutput39 _6245_/Q vssd1 vssd1 vccd1 vccd1 io_out[25] sky130_fd_sc_hd__buf_12
Xoutput17 _6296_/X vssd1 vssd1 vccd1 vccd1 io_oeb[27] sky130_fd_sc_hd__buf_12
Xoutput28 _6085_/Q vssd1 vssd1 vccd1 vccd1 io_out[15] sky130_fd_sc_hd__buf_12
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3559_ _3559_/A _3559_/B vssd1 vssd1 vccd1 vccd1 _5711_/A sky130_fd_sc_hd__nand2_1
X_5229_ _4398_/B _5218_/X _5220_/Y _5228_/X vssd1 vssd1 vccd1 vccd1 _5229_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6295__A _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4104__D_N _5107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4543__A _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold603_A _6237_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4004__A2 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5752__A2 _4943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3606__B _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5093__B _5093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5268__A1 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5313__S _5313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4600_ _5937_/Q _5920_/Q _5928_/Q _6028_/Q _4712_/S1 _4712_/S0 vssd1 vssd1 vccd1
+ vccd1 _4600_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5743__A2 _4895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5580_ _6159_/Q _5507_/Y _5508_/X vssd1 vssd1 vccd1 vccd1 _5582_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__4951__A0 _6157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4599__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4531_ _4531_/A _4531_/B vssd1 vssd1 vccd1 vccd1 _4531_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold316 _5847_/X vssd1 vssd1 vccd1 vccd1 _6245_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4462_ _3446_/A _4427_/A _4484_/A _3250_/D _3479_/A vssd1 vssd1 vccd1 vccd1 _4462_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold305 _5997_/Q vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
X_6201_ _6238_/CLK _6201_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6201_/Q sky130_fd_sc_hd__dfrtp_4
Xhold349 _6182_/Q vssd1 vssd1 vccd1 vccd1 hold349/X sky130_fd_sc_hd__dlygate4sd3_1
X_3413_ _3407_/X _3409_/X _3410_/Y _3412_/X _4485_/B vssd1 vssd1 vccd1 vccd1 _3413_/X
+ sky130_fd_sc_hd__o41a_1
Xhold338 _6129_/Q vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold327 _4128_/X vssd1 vssd1 vccd1 vccd1 _5915_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4393_ _4124_/A _4389_/X _4392_/X _4737_/B vssd1 vssd1 vccd1 vccd1 _4393_/X sky130_fd_sc_hd__o211a_1
X_3344_ _3539_/B hold38/X _3344_/S vssd1 vssd1 vccd1 vccd1 _3344_/X sky130_fd_sc_hd__mux2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6132_ _6192_/CLK _6132_/D vssd1 vssd1 vccd1 vccd1 _6132_/Q sky130_fd_sc_hd__dfxtp_1
X_6063_ _6206_/CLK _6063_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6063_/Q sky130_fd_sc_hd__dfrtp_2
X_3275_ _3275_/A _3275_/B vssd1 vssd1 vccd1 vccd1 _5216_/A sky130_fd_sc_hd__nand2_8
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5014_ _3270_/X _5011_/X _5013_/X _4824_/B vssd1 vssd1 vccd1 vccd1 _5014_/X sky130_fd_sc_hd__a22o_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5916_ _6144_/CLK _5916_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _5916_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_48_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5847_ _5773_/A _5846_/X _5836_/Y hold315/X vssd1 vssd1 vccd1 vccd1 _5847_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_29_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5778_ _6240_/Q hold448/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5778_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5734__A2 _4865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3745__A1 _5116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4729_ _4729_/A _4729_/B _4729_/C _4729_/D vssd1 vssd1 vccd1 vccd1 _4729_/X sky130_fd_sc_hd__or4_1
XANTENNA__5803__A2_N _5352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4302__S _4309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5360__C _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3681__B1 _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5308__S _5313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3595__S0 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3352__A _5216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3060_ _4486_/A _4406_/A vssd1 vssd1 vccd1 vccd1 _3511_/D sky130_fd_sc_hd__nor2_1
XANTENNA__5110__B1 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3071__B _3694_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5701_ _6187_/Q _6203_/Q _5701_/S vssd1 vssd1 vccd1 vccd1 _5701_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_85_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3962_ _6002_/Q _5963_/Q _3982_/S vssd1 vssd1 vccd1 vccd1 _3962_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3893_ _4223_/A _5053_/B vssd1 vssd1 vccd1 vccd1 _3893_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4911__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5632_ _5694_/A _5631_/X _4911_/Y vssd1 vssd1 vccd1 vccd1 _5632_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__5716__A2 _4779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4924__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5563_ _6058_/Q _5595_/S _5607_/B1 _5562_/X vssd1 vssd1 vccd1 vccd1 _5563_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3727__A1 _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4514_ _4512_/X _4514_/B vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5494_ _6240_/Q hold427/X _5497_/S vssd1 vssd1 vccd1 vccd1 _5494_/X sky130_fd_sc_hd__mux2_1
Xhold124 _5923_/Q vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 _6009_/Q vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 _5301_/X vssd1 vssd1 vccd1 vccd1 _6148_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 _6001_/Q vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5742__A _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold146 _4302_/X vssd1 vssd1 vccd1 vccd1 _5965_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 _5926_/Q vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ _4737_/A _4445_/B vssd1 vssd1 vccd1 vccd1 _4445_/Y sky130_fd_sc_hd__nor2_1
Xhold168 _5995_/Q vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
X_4376_ _5773_/A _5629_/A vssd1 vssd1 vccd1 vccd1 _5020_/S sky130_fd_sc_hd__nor2_4
Xhold179 _6151_/Q vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
X_6115_ _6119_/CLK _6115_/D vssd1 vssd1 vccd1 vccd1 _6115_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3327_ _4398_/A _3411_/B vssd1 vssd1 vccd1 vccd1 _3496_/C sky130_fd_sc_hd__nand2_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5652__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3258_ _3200_/A _3543_/B _3257_/X vssd1 vssd1 vccd1 vccd1 _3258_/X sky130_fd_sc_hd__o21ba_1
X_6046_ _6170_/CLK _6046_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6046_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4077__B _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3189_ _4398_/B _3540_/A vssd1 vssd1 vccd1 vccd1 _3543_/B sky130_fd_sc_hd__or2_4
XANTENNA__4792__S _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5168__B1 _3739_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4821__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5636__B _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3603__C _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3654__A0 _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5159__B1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3347__A _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4382__A1 _4451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4877__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4230_ _5926_/Q _3588_/X _3603_/X _6018_/Q vssd1 vssd1 vccd1 vccd1 _4230_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4161_ _4174_/B _4161_/B vssd1 vssd1 vccd1 vccd1 _5054_/C sky130_fd_sc_hd__xor2_1
XANTENNA__5634__A1 _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4437__A2 _3264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5095__C1 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4092_ _3488_/A _3543_/B _5498_/B _4065_/X vssd1 vssd1 vccd1 vccd1 _4092_/X sky130_fd_sc_hd__a31o_1
X_3112_ _3112_/A _3148_/B _4094_/D vssd1 vssd1 vccd1 vccd1 _4412_/B sky130_fd_sc_hd__and3_2
X_3043_ _3654_/S _4739_/A vssd1 vssd1 vccd1 vccd1 _4061_/C sky130_fd_sc_hd__nand2_4
XANTENNA__4842__C1 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4994_ _4990_/B _4993_/X _5011_/S vssd1 vssd1 vccd1 vccd1 _4994_/X sky130_fd_sc_hd__mux2_1
X_3945_ _4014_/A _4005_/B _3943_/X vssd1 vssd1 vccd1 vccd1 _3945_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5615_ _5616_/A _5616_/B vssd1 vssd1 vccd1 vccd1 _5615_/X sky130_fd_sc_hd__and2b_1
X_3876_ _4135_/A _4135_/B vssd1 vssd1 vccd1 vccd1 _5053_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout137_A _6165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5546_ _5566_/S _5544_/X _5545_/Y vssd1 vssd1 vccd1 vccd1 _5546_/X sky130_fd_sc_hd__o21a_1
X_5477_ _5477_/A vssd1 vssd1 vccd1 vccd1 _5477_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_14_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3581__C1 _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4787__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4428_ _5502_/D _4772_/C _4772_/D vssd1 vssd1 vccd1 vccd1 _5338_/C sky130_fd_sc_hd__or3_1
X_4359_ _4193_/X hold286/X _4363_/S vssd1 vssd1 vccd1 vccd1 _6023_/D sky130_fd_sc_hd__mux2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5625__A1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6029_ _6029_/CLK _6029_/D vssd1 vssd1 vccd1 vccd1 _6029_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_5_wb_clk_i _5978_/CLK vssd1 vssd1 vccd1 vccd1 _6102_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout74 _4239_/A vssd1 vssd1 vccd1 vccd1 _4223_/A sky130_fd_sc_hd__buf_4
Xfanout63 _5702_/A2 vssd1 vssd1 vccd1 vccd1 _5595_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout85 _3591_/Y vssd1 vssd1 vccd1 vccd1 _3739_/S sky130_fd_sc_hd__clkbuf_4
Xfanout96 _4418_/A vssd1 vssd1 vccd1 vccd1 _4094_/B sky130_fd_sc_hd__buf_4
XANTENNA__4697__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5313__A0 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5864__A1 _6115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3614__B _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3642__A3 _6113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3730_ _4234_/A _3730_/B _3730_/C vssd1 vssd1 vccd1 vccd1 _3730_/X sky130_fd_sc_hd__and3_1
XFILLER_0_27_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3661_ _3920_/A _5395_/A _3658_/X _6113_/Q vssd1 vssd1 vccd1 vccd1 _3661_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5400_ _5400_/A _5400_/B vssd1 vssd1 vccd1 vccd1 _5400_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_23_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3592_ _4461_/A _4034_/S vssd1 vssd1 vccd1 vccd1 _3592_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_42_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5331_ _6142_/Q _3995_/B _3998_/Y vssd1 vssd1 vccd1 vccd1 _5332_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5262_ hold506/X _5251_/Y _5252_/Y _6213_/Q _5261_/X vssd1 vssd1 vccd1 vccd1 _5262_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5855__B2 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4213_ hold72/A _3611_/X _3613_/X _5933_/Q vssd1 vssd1 vccd1 vccd1 _4213_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_76_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5193_ _6178_/Q _5104_/Y _5106_/Y _6210_/Q vssd1 vssd1 vccd1 vccd1 _5204_/A sky130_fd_sc_hd__a22o_1
X_4144_ _4250_/A _5246_/A vssd1 vssd1 vccd1 vccd1 _4146_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__6169__RESET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4075_ _6052_/Q _6053_/Q _4075_/S vssd1 vssd1 vccd1 vccd1 _4075_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3026_ _4417_/A _3180_/B vssd1 vssd1 vccd1 vccd1 _5502_/B sky130_fd_sc_hd__nor2_4
XANTENNA__4830__A2 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4074__C _5250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4977_ _6241_/Q _5008_/B vssd1 vssd1 vccd1 vccd1 _4977_/X sky130_fd_sc_hd__and2_1
X_3928_ hold17/X _4253_/A2 _3893_/Y _3927_/X vssd1 vssd1 vccd1 vccd1 _3928_/X sky130_fd_sc_hd__o22a_1
X_3859_ _3859_/A _3859_/B vssd1 vssd1 vccd1 vccd1 _3860_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5529_ _5528_/X _6055_/Q _5595_/S vssd1 vssd1 vccd1 vccd1 _5529_/X sky130_fd_sc_hd__mux2_1
XANTENNA__6298__A _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4649__A2 _4612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3434__B _3434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4980__S _5011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5782__A0 _6172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4585__A1 _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4888__A2 _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3360__A _6129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4900_ _4901_/A _4901_/B vssd1 vssd1 vccd1 vccd1 _4918_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4890__S _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5880_ input3/X _5890_/B vssd1 vssd1 vccd1 vccd1 _5880_/X sky130_fd_sc_hd__and2_1
XFILLER_0_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4831_ _6057_/Q _4764_/X _4829_/X _4830_/Y vssd1 vssd1 vccd1 vccd1 _4831_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4576__A1 _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3379__A2 _4486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4762_ _6048_/Q _4762_/B vssd1 vssd1 vccd1 vccd1 _4763_/B sky130_fd_sc_hd__and2_2
X_4693_ _6159_/Q _4620_/Y _4692_/X vssd1 vssd1 vccd1 vccd1 _4693_/X sky130_fd_sc_hd__o21a_1
X_3713_ _3713_/A _3713_/B vssd1 vssd1 vccd1 vccd1 _3713_/Y sky130_fd_sc_hd__nand2_1
X_3644_ _6072_/Q _6071_/Q _6073_/Q vssd1 vssd1 vccd1 vccd1 _3655_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_15_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3575_ _3513_/A _3571_/X _3559_/B vssd1 vssd1 vccd1 vccd1 _5021_/C sky130_fd_sc_hd__a21oi_1
X_6294_ _6299_/A vssd1 vssd1 vccd1 vccd1 _6294_/X sky130_fd_sc_hd__buf_1
X_5314_ _5314_/A _5566_/S vssd1 vssd1 vccd1 vccd1 _5314_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3551__A2 _4446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5245_ _5245_/A _5245_/B vssd1 vssd1 vccd1 vccd1 _5245_/Y sky130_fd_sc_hd__nor2_2
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ _5176_/A _5176_/B _5176_/C vssd1 vssd1 vccd1 vccd1 _5176_/X sky130_fd_sc_hd__or3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_4127_ _4124_/X _4126_/X _3405_/B vssd1 vssd1 vccd1 vccd1 _4127_/Y sky130_fd_sc_hd__a21oi_1
X_4058_ _4749_/A _4058_/B vssd1 vssd1 vccd1 vccd1 _4058_/X sky130_fd_sc_hd__or2_1
X_3009_ _4485_/A _3203_/B _3210_/A vssd1 vssd1 vccd1 vccd1 _3507_/C sky130_fd_sc_hd__nand3b_4
XFILLER_0_66_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4305__S _4309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5516__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5363__C _5363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5819__A1 _6241_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5819__B2 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4975__S _5020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_207 vssd1 vssd1 vccd1 vccd1 ci2406_z80_207/HI io_oeb[22] sky130_fd_sc_hd__conb_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4007__A0 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4558__A1 _4850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold509 _5258_/X vssd1 vssd1 vccd1 vccd1 _6135_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3360_ _6129_/Q _3368_/C vssd1 vssd1 vccd1 vccd1 _3376_/B sky130_fd_sc_hd__and2_1
XANTENNA__4730__A1 _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5372_/A _5372_/B _5029_/X _5479_/S vssd1 vssd1 vccd1 vccd1 _5030_/X sky130_fd_sc_hd__o31a_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3291_ _4483_/A _3193_/X _4116_/B _3545_/A _3709_/B vssd1 vssd1 vccd1 vccd1 _3291_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3297__A1 _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5038__A2 _6178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3521__C _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5443__C1 _6176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4246__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5932_ _6031_/CLK hold69/X vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__4797__A1 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4797__B2 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5863_ hold323/X _5836_/A _5862_/X _5245_/A vssd1 vssd1 vccd1 vccd1 _5863_/X sky130_fd_sc_hd__o22a_1
X_5794_ _5868_/S _5794_/B vssd1 vssd1 vccd1 vccd1 _5794_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_56_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4814_ _4814_/A _4814_/B _4814_/C vssd1 vssd1 vccd1 vccd1 _4814_/X sky130_fd_sc_hd__or3_1
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3221__A1 _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4745_ _5164_/A1 hold618/X _4927_/S _4438_/X vssd1 vssd1 vccd1 vccd1 _6072_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4676_ _4676_/A _4676_/B _4676_/C vssd1 vssd1 vccd1 vccd1 _4677_/B sky130_fd_sc_hd__and3_1
XFILLER_0_71_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3627_ _6135_/Q _3629_/B vssd1 vssd1 vccd1 vccd1 _3628_/B sky130_fd_sc_hd__and2_1
XFILLER_0_101_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4721__A1 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput29 _6086_/Q vssd1 vssd1 vccd1 vccd1 io_out[16] sky130_fd_sc_hd__buf_12
Xoutput18 _6297_/X vssd1 vssd1 vccd1 vccd1 io_oeb[28] sky130_fd_sc_hd__buf_12
X_3558_ _3457_/A _3555_/X _3557_/X vssd1 vssd1 vccd1 vccd1 _3559_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_101_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3489_ _3485_/Y _4613_/C _3488_/X _3476_/X _5424_/B vssd1 vssd1 vccd1 vccd1 _3523_/B
+ sky130_fd_sc_hd__o32a_1
X_5228_ _5225_/B _5228_/B vssd1 vssd1 vccd1 vccd1 _5228_/X sky130_fd_sc_hd__and2b_1
X_5159_ _5923_/Q _5200_/A2 _5200_/B1 _6031_/Q _5182_/S vssd1 vssd1 vccd1 vccd1 _5160_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA__5434__C1 _5341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4788__A1 _4787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3460__A1 _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4035__S _4035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4004__A3 _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3212__A1 _3713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3175__A _5502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5390__A _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4571__S0 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3622__B _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5440__A2 _5363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3451__A1 _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3987__C1 _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3069__B _4614_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4400__B1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4530_ _4514_/B _4516_/B _4512_/X vssd1 vssd1 vccd1 vccd1 _4531_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_13_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold317 _6246_/Q vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4461_ _4461_/A _4461_/B vssd1 vssd1 vccd1 vccd1 _6053_/D sky130_fd_sc_hd__xnor2_1
Xhold306 _4330_/X vssd1 vssd1 vccd1 vccd1 _5997_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6200_ _6203_/CLK _6200_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6200_/Q sky130_fd_sc_hd__dfrtp_4
Xhold339 _6091_/Q vssd1 vssd1 vccd1 vccd1 hold339/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3412_ _5502_/B _3479_/A _3477_/C _3412_/D vssd1 vssd1 vccd1 vccd1 _3412_/X sky130_fd_sc_hd__or4_1
Xhold328 _6082_/Q vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4392_ _4392_/A _4392_/B _4054_/X vssd1 vssd1 vccd1 vccd1 _4392_/X sky130_fd_sc_hd__or3b_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6131_ _6190_/CLK _6131_/D vssd1 vssd1 vccd1 vccd1 _6131_/Q sky130_fd_sc_hd__dfxtp_1
X_3343_ _3343_/A _3343_/B _3342_/X vssd1 vssd1 vccd1 vccd1 _3343_/Y sky130_fd_sc_hd__nor3b_1
XFILLER_0_0_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ _6218_/CLK _6062_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6062_/Q sky130_fd_sc_hd__dfrtp_2
X_3274_ _6038_/Q _4104_/B vssd1 vssd1 vccd1 vccd1 _3275_/B sky130_fd_sc_hd__nor2_2
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _6161_/Q _5012_/X _5013_/S vssd1 vssd1 vccd1 vccd1 _5013_/X sky130_fd_sc_hd__mux2_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout167_A _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5431__A2 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3442__A1 _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5915_ _6170_/CLK _5915_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _5915_/Q sky130_fd_sc_hd__dfrtp_1
X_5846_ _3707_/X _5837_/B _5837_/X _5845_/Y vssd1 vssd1 vccd1 vccd1 _5846_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2989_ _2989_/A vssd1 vssd1 vccd1 vccd1 _2989_/Y sky130_fd_sc_hd__inv_2
X_5777_ _6239_/Q hold488/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5777_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5195__B2 _6160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4942__A1 _4941_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4728_ _4728_/A _4728_/B _4728_/C _4772_/C vssd1 vssd1 vccd1 vccd1 _4729_/D sky130_fd_sc_hd__or4_1
X_4659_ _4699_/A _4659_/B vssd1 vssd1 vccd1 vccd1 _4676_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3426__C _3694_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4538__B _4538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3736__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_1_wb_clk_i_A _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3595__S1 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6235_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_54_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3424__A1 _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3961_ _5986_/Q _5994_/Q _3982_/S vssd1 vssd1 vccd1 vccd1 _3961_/X sky130_fd_sc_hd__mux2_1
X_5700_ _5687_/A _5691_/A _5698_/Y _5511_/X vssd1 vssd1 vccd1 vccd1 _5700_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_97_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4621__B1 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3424__B2 _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3892_ _4135_/C _3892_/B vssd1 vssd1 vccd1 vccd1 _5053_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4911__B _4915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5631_ hold454/X _5702_/A2 _5702_/B1 _5630_/X vssd1 vssd1 vccd1 vccd1 _5631_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5177__A1 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4403__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3808__A _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5562_ _6058_/Q _6192_/Q _5606_/S vssd1 vssd1 vccd1 vccd1 _5562_/X sky130_fd_sc_hd__mux2_1
X_4513_ _4575_/A _4512_/B _4512_/C vssd1 vssd1 vccd1 vccd1 _4514_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5493_ _6239_/Q hold398/X _5497_/S vssd1 vssd1 vccd1 vccd1 _5493_/X sky130_fd_sc_hd__mux2_1
Xhold125 _4194_/X vssd1 vssd1 vccd1 vccd1 _5923_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold103 _4334_/X vssd1 vssd1 vccd1 vccd1 _6001_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold114 _6002_/Q vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold158 _4243_/X vssd1 vssd1 vccd1 vccd1 _5926_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _4343_/X vssd1 vssd1 vccd1 vccd1 _6009_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 _5993_/Q vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
X_4444_ _4433_/B _5838_/B _4738_/A _4737_/A vssd1 vssd1 vccd1 vccd1 _4444_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5742__B _5771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4375_ _5629_/A vssd1 vssd1 vccd1 vccd1 _4375_/Y sky130_fd_sc_hd__inv_2
Xhold169 _5937_/Q vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
X_6114_ _6119_/CLK _6114_/D vssd1 vssd1 vccd1 vccd1 _6114_/Q sky130_fd_sc_hd__dfxtp_2
X_3326_ _4398_/A _3411_/B vssd1 vssd1 vccd1 vccd1 _3334_/B sky130_fd_sc_hd__and2_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ _6170_/CLK _6045_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6045_/Q sky130_fd_sc_hd__dfrtp_1
X_3257_ _4390_/A _4759_/A _3298_/A _3255_/X _3256_/X vssd1 vssd1 vccd1 vccd1 _3257_/X
+ sky130_fd_sc_hd__a311o_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5101__B2 _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3188_ _4398_/B _3540_/A vssd1 vssd1 vccd1 vccd1 _3713_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_95_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4374__A _5705_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3415__A1 _5918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5829_ hold591/X _5791_/X _5828_/X _5341_/A vssd1 vssd1 vccd1 vccd1 _5829_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_8_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3718__A _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4313__S _4318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4679__B1 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3406__A1 _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3406__B2 _3434_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4382__A2 _4391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3066__C _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4160_ _4219_/A _4143_/Y _4147_/A vssd1 vssd1 vccd1 vccd1 _4161_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__3363__A _5216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3111_ _3777_/A _3643_/A _4433_/B _5489_/C _5356_/A vssd1 vssd1 vccd1 vccd1 _3111_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4893__S _4926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4091_ _3112_/A _4077_/X _4090_/X _5220_/A vssd1 vssd1 vccd1 vccd1 _5120_/A sky130_fd_sc_hd__a22o_4
X_3042_ _3777_/A _4735_/A vssd1 vssd1 vccd1 vccd1 _3193_/C sky130_fd_sc_hd__nor2_4
XANTENNA__4842__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6205__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4993_ _6202_/Q _6068_/Q _6038_/Q vssd1 vssd1 vccd1 vccd1 _4993_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3944_ _3944_/A _3944_/B vssd1 vssd1 vccd1 vccd1 _4005_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3875_ _4250_/A _3875_/B vssd1 vssd1 vccd1 vccd1 _4135_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5614_ _5602_/A _5685_/B _5603_/X vssd1 vssd1 vccd1 vccd1 _5616_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5545_ _5538_/A _5566_/S _5670_/A vssd1 vssd1 vccd1 vccd1 _5545_/Y sky130_fd_sc_hd__a21oi_1
X_5476_ _3959_/A _5475_/X _5487_/S vssd1 vssd1 vccd1 vccd1 _5477_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5322__A1 _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4427_ _4427_/A _4427_/B _4427_/C _4427_/D vssd1 vssd1 vccd1 vccd1 _4429_/B sky130_fd_sc_hd__or4_1
X_4358_ _4180_/X hold186/X _4363_/S vssd1 vssd1 vccd1 vccd1 _6022_/D sky130_fd_sc_hd__mux2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4289_ _4226_/X hold166/X _4291_/S vssd1 vssd1 vccd1 vccd1 _4289_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5086__B1 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4508__S0 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _4038_/A _3309_/B vssd1 vssd1 vccd1 vccd1 _4731_/S sky130_fd_sc_hd__nand2_2
XANTENNA__5625__A2 _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6028_ _6110_/CLK _6028_/D vssd1 vssd1 vccd1 vccd1 _6028_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4308__S _4309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5647__B _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout53 _5020_/S vssd1 vssd1 vccd1 vccd1 _4927_/S sky130_fd_sc_hd__buf_6
Xfanout64 _4761_/X vssd1 vssd1 vccd1 vccd1 _5702_/A2 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout86 _4118_/Y vssd1 vssd1 vccd1 vccd1 _4119_/B sky130_fd_sc_hd__buf_4
XFILLER_0_51_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3572__B1 _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5313__A1 hold636/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5077__B1 _4750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3630__B _6172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5838__A _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6050__RESET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3660_ _6135_/Q _3650_/X _3659_/X _3624_/Y vssd1 vssd1 vccd1 vccd1 _3660_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_15_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3591_ _3591_/A _4034_/S vssd1 vssd1 vccd1 vccd1 _3591_/Y sky130_fd_sc_hd__nor2_1
X_5330_ _5330_/A _5330_/B vssd1 vssd1 vccd1 vccd1 _5348_/S sky130_fd_sc_hd__or2_1
X_5261_ _6155_/Q _5253_/Y _5254_/Y _6237_/Q _5260_/X vssd1 vssd1 vccd1 vccd1 _5261_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5855__A2 _5836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4212_ hold141/X _4211_/X _4262_/S vssd1 vssd1 vccd1 vccd1 _4212_/X sky130_fd_sc_hd__mux2_1
X_5192_ _5023_/A hold388/X _5086_/Y _5191_/X vssd1 vssd1 vccd1 vccd1 _5192_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_44_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6171_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4143_ _5246_/A vssd1 vssd1 vccd1 vccd1 _4143_/Y sky130_fd_sc_hd__inv_2
X_4074_ _6038_/Q _4104_/B _5250_/A _5250_/B vssd1 vssd1 vccd1 vccd1 _4075_/S sky130_fd_sc_hd__or4b_1
X_3025_ _3777_/A _4417_/B vssd1 vssd1 vccd1 vccd1 _3180_/B sky130_fd_sc_hd__or2_2
XFILLER_0_92_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5240__A0 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4976_ _4990_/A _4976_/B vssd1 vssd1 vccd1 vccd1 _4976_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5791__A1 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3927_ _4223_/A _3926_/X _3573_/B vssd1 vssd1 vccd1 vccd1 _3927_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3251__C1 _4439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3268__A _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3858_ _3848_/B _3854_/X _3899_/B _3857_/X vssd1 vssd1 vccd1 vccd1 _3859_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3789_ _4034_/S _3745_/X _3787_/X _3788_/X vssd1 vssd1 vccd1 vccd1 _3789_/X sky130_fd_sc_hd__a22o_2
XANTENNA__5543__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5528_ _6189_/Q _5606_/S _4790_/X vssd1 vssd1 vccd1 vccd1 _5528_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_14_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3715__B _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5459_ hold576/X _3377_/X _5365_/S _5458_/X vssd1 vssd1 vccd1 vccd1 _5459_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3434__C _5875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5470__B1 _5484_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4273__A1 _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4830_ _5551_/A _4815_/B _4764_/X vssd1 vssd1 vccd1 vccd1 _4830_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4472__A _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4761_ _4761_/A _4761_/B vssd1 vssd1 vccd1 vccd1 _4761_/X sky130_fd_sc_hd__or2_2
X_4692_ hold510/X _4612_/X _4691_/Y _4611_/A _4619_/X vssd1 vssd1 vccd1 vccd1 _4692_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3712_ _3545_/Y _3710_/X _3711_/Y _3545_/A _5502_/A vssd1 vssd1 vccd1 vccd1 _3712_/Y
+ sky130_fd_sc_hd__a221oi_4
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3643_ _3643_/A _3643_/B vssd1 vssd1 vccd1 vccd1 _3657_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5313_ input8/X hold636/X _5313_/S vssd1 vssd1 vccd1 vccd1 _6161_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_11_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3574_ _4034_/S _3573_/B _3573_/C _4461_/A vssd1 vssd1 vccd1 vccd1 _3574_/Y sky130_fd_sc_hd__o31ai_2
X_6293_ _6299_/A vssd1 vssd1 vccd1 vccd1 _6293_/X sky130_fd_sc_hd__buf_1
X_5244_ _5250_/A _5250_/B _4409_/X vssd1 vssd1 vccd1 vccd1 _5245_/B sky130_fd_sc_hd__o21a_1
XANTENNA__3839__A1 _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ _6176_/Q _5104_/Y _5129_/Y _6216_/Q _5174_/X vssd1 vssd1 vccd1 vccd1 _5176_/C
+ sky130_fd_sc_hd__a221o_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_4126_ _5502_/A _4126_/B _4613_/C vssd1 vssd1 vccd1 vccd1 _4126_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4057_ _5424_/A _4446_/B _4737_/B vssd1 vssd1 vccd1 vccd1 _4058_/B sky130_fd_sc_hd__o21ai_1
X_3008_ _3210_/A _3203_/B _3148_/C vssd1 vssd1 vccd1 vccd1 _3150_/A sky130_fd_sc_hd__and3_1
XFILLER_0_93_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4959_ _4990_/A _4963_/B vssd1 vssd1 vccd1 vccd1 _4959_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3775__A0 _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3148__D _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4321__S _4327_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_61_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold576_A _6177_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xci2406_z80_208 vssd1 vssd1 vccd1 vccd1 ci2406_z80_208/HI io_oeb[23] sky130_fd_sc_hd__conb_1
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5755__A1 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5755__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4730__A2 _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _4483_/A _3290_/B _3334_/A vssd1 vssd1 vccd1 vccd1 _3290_/X sky130_fd_sc_hd__or3_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5062__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3297__A2 _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3521__D _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5931_ _6035_/CLK _5931_/D vssd1 vssd1 vccd1 vccd1 _5931_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5862_ _3926_/X _5834_/X _5837_/X _5861_/X vssd1 vssd1 vccd1 vccd1 _5862_/X sky130_fd_sc_hd__o22a_1
X_5793_ _6236_/Q _5791_/X _5792_/X _5764_/B vssd1 vssd1 vccd1 vccd1 _5793_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5746__A1 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5746__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4813_ _6156_/Q _5008_/B _4811_/X _4999_/A1 vssd1 vssd1 vccd1 vccd1 _4814_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4744_ _5164_/A1 _5333_/B _4927_/S _4743_/X vssd1 vssd1 vccd1 vccd1 _4744_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3221__A2 _6127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4675_ _4647_/A _4647_/C _4658_/Y _4647_/B vssd1 vssd1 vccd1 vccd1 _4676_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout112_A _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3626_ _5333_/B _6113_/Q vssd1 vssd1 vccd1 vccd1 _3629_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_101_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4182__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput19 _6298_/X vssd1 vssd1 vccd1 vccd1 io_oeb[29] sky130_fd_sc_hd__buf_12
X_3557_ _3545_/Y _3547_/X _3556_/Y _3541_/X vssd1 vssd1 vccd1 vccd1 _3557_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3980__S _4035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5227_ _4398_/B _3353_/B _5217_/A _5226_/X vssd1 vssd1 vccd1 vccd1 _5227_/X sky130_fd_sc_hd__a22o_1
X_3488_ _3488_/A _3488_/B _4614_/D vssd1 vssd1 vccd1 vccd1 _3488_/X sky130_fd_sc_hd__or3_1
X_5158_ _6015_/Q _5200_/A2 _5200_/B1 _5948_/Q _4256_/S vssd1 vssd1 vccd1 vccd1 _5160_/A
+ sky130_fd_sc_hd__o221a_1
X_4109_ hold91/X _3737_/X _4115_/S vssd1 vssd1 vccd1 vccd1 _5907_/D sky130_fd_sc_hd__mux2_1
X_5089_ _4460_/A _4094_/B _4094_/C _4077_/X vssd1 vssd1 vccd1 vccd1 _5089_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_66_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4824__B _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4316__S _4318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5737__A1 _4116_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5737__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3212__A2 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4571__S1 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5425__B1 _5426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5610__S _5705_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3451__A2 _4043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5728__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5728__A1 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4750__A _4750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4460_ _4460_/A _5875_/A _4460_/C _5341_/A vssd1 vssd1 vccd1 vccd1 _4461_/B sky130_fd_sc_hd__and4_1
Xhold307 _6132_/Q vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold318 _5851_/X vssd1 vssd1 vccd1 vccd1 _6246_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3411_ _4726_/A _3411_/B _3543_/A _3411_/D vssd1 vssd1 vccd1 vccd1 _3412_/D sky130_fd_sc_hd__or4_1
X_4391_ _6127_/Q _4391_/B vssd1 vssd1 vccd1 vccd1 _4392_/B sky130_fd_sc_hd__nor2_1
Xhold329 _4849_/X vssd1 vssd1 vccd1 vccd1 _6082_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3342_ _6164_/Q _4497_/S _3344_/S vssd1 vssd1 vccd1 vccd1 _3342_/X sky130_fd_sc_hd__mux2_1
X_6130_ _6130_/CLK _6130_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6130_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6061_ _6119_/CLK _6061_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6061_/Q sky130_fd_sc_hd__dfrtp_4
X_3273_ _6052_/Q _6051_/Q vssd1 vssd1 vccd1 vccd1 _5011_/S sky130_fd_sc_hd__or2_4
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _6069_/Q _5012_/B vssd1 vssd1 vccd1 vccd1 _5012_/X sky130_fd_sc_hd__xor2_1
XANTENNA__3675__C1 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3690__A2 _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5520__S _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5914_ _6144_/CLK _5914_/D vssd1 vssd1 vccd1 vccd1 _5914_/Q sky130_fd_sc_hd__dfxtp_1
X_5845_ _5845_/A vssd1 vssd1 vccd1 vccd1 _5845_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5719__A1 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5719__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5776_ _6238_/Q hold437/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5776_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2988_ _6160_/Q vssd1 vssd1 vccd1 vccd1 _4570_/B sky130_fd_sc_hd__inv_2
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4727_ _4727_/A _4727_/B _4727_/C vssd1 vssd1 vccd1 vccd1 _4729_/C sky130_fd_sc_hd__or3_1
X_4658_ _4699_/A _4659_/B vssd1 vssd1 vccd1 vccd1 _4658_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4155__B1 _3615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3609_ _2966_/Y _3724_/S _3608_/X _3616_/B vssd1 vssd1 vccd1 vccd1 _3609_/Y sky130_fd_sc_hd__a211oi_1
X_4589_ _6211_/Q _4879_/B _4589_/S vssd1 vssd1 vccd1 vccd1 _4591_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4458__A1 _3694_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6259_ _6259_/CLK _6259_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6259_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4394__B1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4241__S0 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4449__A1 _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4449__B2 _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5110__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5464__A2_N _5363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3960_ _3597_/X _3959_/A _3539_/Y vssd1 vssd1 vccd1 vccd1 _3960_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3424__A2 _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4082__C1 _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3891_ _4135_/A _4135_/B _3874_/X vssd1 vssd1 vccd1 vccd1 _3892_/B sky130_fd_sc_hd__a21o_1
X_5630_ _6181_/Q _6197_/Q _5701_/S vssd1 vssd1 vccd1 vccd1 _5630_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4924__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5561_ _2993_/A _5560_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _5561_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5492_ _6238_/Q hold349/X _5497_/S vssd1 vssd1 vccd1 vccd1 _5492_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4512_ _4575_/A _4512_/B _4512_/C vssd1 vssd1 vccd1 vccd1 _4512_/X sky130_fd_sc_hd__and3_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold104 _5985_/Q vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 _5903_/Q vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 _4335_/X vssd1 vssd1 vccd1 vccd1 _6002_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 _5931_/Q vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 _5925_/Q vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold148 _4325_/X vssd1 vssd1 vccd1 vccd1 _5993_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ _4441_/X _4442_/X _2957_/Y vssd1 vssd1 vccd1 vccd1 _4443_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5515__S _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4374_ _5705_/S _5762_/A vssd1 vssd1 vccd1 vccd1 _5629_/A sky130_fd_sc_hd__or2_4
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6113_ _6119_/CLK _6113_/D vssd1 vssd1 vccd1 vccd1 _6113_/Q sky130_fd_sc_hd__dfxtp_4
X_3325_ _3290_/B _3314_/X _4427_/B _3498_/A vssd1 vssd1 vccd1 vccd1 _3325_/X sky130_fd_sc_hd__o31a_1
XANTENNA__3543__B _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5637__B1 _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6044_ _6060_/CLK _6044_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6044_/Q sky130_fd_sc_hd__dfrtp_1
X_3256_ _3302_/A _3184_/A _5093_/B _3542_/B _3196_/B vssd1 vssd1 vccd1 vccd1 _3256_/X
+ sky130_fd_sc_hd__a32o_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3663__A2 _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4860__A1 _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3187_ _4417_/A _3187_/B vssd1 vssd1 vccd1 vccd1 _4045_/A sky130_fd_sc_hd__or2_2
XANTENNA__4374__B _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3415__A2 _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5828_ _6243_/Q _5352_/A _5457_/A hold468/X vssd1 vssd1 vccd1 vccd1 _5828_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_76_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5168__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5759_ _3926_/X _5771_/S _5742_/Y _5758_/X vssd1 vssd1 vccd1 vccd1 _5759_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout92_A _5007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold660 _6005_/Q vssd1 vssd1 vccd1 vccd1 hold660/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold656_A _6131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4603__A1 _4895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3909__A _6172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5159__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4504__S _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3342__A1 _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3204__A_N _3434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3110_ _3249_/A _3210_/C vssd1 vssd1 vccd1 vccd1 _4445_/B sky130_fd_sc_hd__or2_4
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5095__A1 _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4090_ _3539_/A _4084_/X _4086_/X _4089_/X _4618_/B vssd1 vssd1 vccd1 vccd1 _4090_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5070__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4475__A _6129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3041_ _3507_/C _4051_/B _3249_/B _3643_/B vssd1 vssd1 vccd1 vccd1 _3041_/Y sky130_fd_sc_hd__a211oi_1
XANTENNA__4842__B2 _4836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4992_ _6218_/Q _5009_/A2 _4769_/Y _4990_/B _4991_/X vssd1 vssd1 vccd1 vccd1 _4992_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3943_ _4005_/A _3944_/A _3944_/B vssd1 vssd1 vccd1 vccd1 _3943_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_46_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3874_ _4234_/A _3875_/B vssd1 vssd1 vccd1 vccd1 _3874_/X sky130_fd_sc_hd__and2_1
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5613_ _5613_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5616_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__3538__B _6166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5544_ _5543_/X _6056_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _5544_/X sky130_fd_sc_hd__mux2_1
X_5475_ _5472_/X _5474_/X _5475_/S vssd1 vssd1 vccd1 vccd1 _5475_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3581__A1 _3513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4426_ _4426_/A _4728_/C _4483_/B _4614_/C vssd1 vssd1 vccd1 vccd1 _4427_/D sky130_fd_sc_hd__or4_1
XFILLER_0_1_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4357_ _4165_/X hold201/X _4363_/S vssd1 vssd1 vccd1 vccd1 _4357_/X sky130_fd_sc_hd__mux2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _4211_/X hold265/X _4291_/S vssd1 vssd1 vccd1 vccd1 _5949_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5086__A1 _5120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4508__S1 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3308_ _3303_/X _3304_/X _3307_/Y _3540_/A vssd1 vssd1 vccd1 vccd1 _3321_/B sky130_fd_sc_hd__a31o_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ _6111_/CLK _6027_/D vssd1 vssd1 vccd1 vccd1 _6027_/Q sky130_fd_sc_hd__dfxtp_1
X_3239_ _3777_/A _5356_/A _3643_/A vssd1 vssd1 vccd1 vccd1 _3239_/X sky130_fd_sc_hd__or3b_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4833__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4324__S _4327_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout54 _5705_/S vssd1 vssd1 vccd1 vccd1 _5566_/S sky130_fd_sc_hd__buf_6
Xfanout65 _3579_/Y vssd1 vssd1 vccd1 vccd1 _3988_/A sky130_fd_sc_hd__buf_4
Xfanout87 _4118_/Y vssd1 vssd1 vccd1 vccd1 _5694_/A sky130_fd_sc_hd__buf_4
Xfanout76 _5698_/B vssd1 vssd1 vccd1 vccd1 _5685_/B sky130_fd_sc_hd__clkbuf_8
Xfanout98 _4765_/Y vssd1 vssd1 vccd1 vccd1 _5606_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5849__A0 _6115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3572__A1 _3513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold490 _6201_/Q vssd1 vssd1 vccd1 vccd1 _5679_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4994__S _5011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6211__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5077__B2 _4391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5838__B _5838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4683__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3590_ _5297_/A _4132_/A vssd1 vssd1 vccd1 vccd1 _4035_/S sky130_fd_sc_hd__nor2_4
X_5260_ _4157_/Y _5259_/B _5248_/Y _5259_/Y vssd1 vssd1 vccd1 vccd1 _5260_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_50_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4211_ _4209_/X _4210_/X _4242_/S vssd1 vssd1 vccd1 vccd1 _4211_/X sky130_fd_sc_hd__mux2_2
X_5191_ _6217_/Q _5129_/Y _5188_/X _5190_/X vssd1 vssd1 vccd1 vccd1 _5191_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_76_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4142_ _4142_/A _4142_/B vssd1 vssd1 vccd1 vccd1 _5246_/A sky130_fd_sc_hd__nand2_2
XANTENNA__3079__B1 _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4073_ _4058_/B _4062_/X _4072_/X _4618_/B vssd1 vssd1 vccd1 vccd1 _5250_/B sky130_fd_sc_hd__o22a_4
X_3024_ _3112_/A _4094_/D _3203_/B vssd1 vssd1 vccd1 vccd1 _4417_/B sky130_fd_sc_hd__or3b_4
XFILLER_0_92_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_13_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6032_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4975_ hold365/X _4974_/X _5020_/S vssd1 vssd1 vccd1 vccd1 _4975_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3926_ _3925_/X hold388/X _3958_/S vssd1 vssd1 vccd1 vccd1 _3926_/X sky130_fd_sc_hd__mux2_4
XANTENNA_fanout142_A hold652/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5791__A2 _5352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3857_ _3639_/X _3855_/A _3856_/Y _5024_/B vssd1 vssd1 vccd1 vccd1 _3857_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3983__S _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3788_ hold7/X _4253_/A2 _3671_/B vssd1 vssd1 vccd1 vccd1 _3788_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_6_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_25_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5527_ _5540_/B _5527_/B vssd1 vssd1 vccd1 vccd1 _5527_/Y sky130_fd_sc_hd__nor2_1
X_5458_ _6233_/Q _5340_/Y _5457_/X _5341_/A vssd1 vssd1 vccd1 vccd1 _5458_/X sky130_fd_sc_hd__o211a_1
X_5389_ _5389_/A _5389_/B vssd1 vssd1 vccd1 vccd1 _5392_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3434__D _3434_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4409_ _4460_/A _4407_/X _4408_/X _4618_/B vssd1 vssd1 vccd1 vccd1 _4409_/X sky130_fd_sc_hd__a22o_2
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5004__A _6160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3609__A2 _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5658__B _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold619_A _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5231__B2 _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4989__S _5020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4737__B _4737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4258__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4472__B _4779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3233__B1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4760_ _3483_/X _4760_/B _4760_/C _4760_/D vssd1 vssd1 vccd1 vccd1 _4761_/B sky130_fd_sc_hd__and4b_1
XANTENNA__6200__RESET_B fanout184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4691_ _4691_/A _4691_/B vssd1 vssd1 vccd1 vccd1 _4691_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__4899__S _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3711_ _4759_/B _3711_/B vssd1 vssd1 vccd1 vccd1 _3711_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3642_ _5024_/A _6135_/Q _6113_/Q _3848_/B _3641_/X vssd1 vssd1 vccd1 vccd1 _5374_/A
+ sky130_fd_sc_hd__o41a_2
X_5312_ input7/X hold630/X _5313_/S vssd1 vssd1 vccd1 vccd1 _6160_/D sky130_fd_sc_hd__mux2_1
X_3573_ _4034_/S _3573_/B _3573_/C vssd1 vssd1 vccd1 vccd1 _3573_/X sky130_fd_sc_hd__or3_2
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4928__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5243_ _3517_/A _5242_/X _3252_/B vssd1 vssd1 vccd1 vccd1 _5243_/X sky130_fd_sc_hd__o21ba_1
X_5174_ _6200_/Q _5119_/Y _5173_/X _5109_/Y vssd1 vssd1 vccd1 vccd1 _5174_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3832__A _3832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_4125_ _4772_/C _4483_/B _4125_/C vssd1 vssd1 vccd1 vccd1 _4126_/B sky130_fd_sc_hd__or3_1
XANTENNA__5461__A1 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4056_ _4056_/A _4056_/B vssd1 vssd1 vccd1 vccd1 _4749_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3007_ _4739_/A _3193_/A _6259_/Q _6258_/Q vssd1 vssd1 vccd1 vccd1 _3182_/A sky130_fd_sc_hd__or4bb_4
XFILLER_0_78_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3072__A_N _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4958_ hold343/X _4957_/X _5020_/S vssd1 vssd1 vccd1 vccd1 _4958_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4972__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3909_ _6172_/Q _3909_/B vssd1 vssd1 vccd1 vccd1 _4005_/A sky130_fd_sc_hd__or2_2
X_4889_ _6195_/Q _4767_/X _4886_/X _4888_/X vssd1 vssd1 vccd1 vccd1 _4889_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3775__A1 _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4602__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4724__B1 _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3461__B _3503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_209 vssd1 vssd1 vccd1 vccd1 ci2406_z80_209/HI io_out[32] sky130_fd_sc_hd__conb_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5452__B2 _3864_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4638__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5755__A2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3518__A1 _3513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5443__A1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4246__A2 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5930_ _6014_/CLK hold55/X vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__dfxtp_1
X_5861_ _6118_/Q _5860_/X _5869_/S vssd1 vssd1 vccd1 vccd1 _5861_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5792_ _6236_/Q _5352_/A _5457_/A hold441/X vssd1 vssd1 vccd1 vccd1 _5792_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__5746__A2 _4915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4812_ _6206_/Q _4768_/Y _4769_/Y _4805_/B _4815_/B vssd1 vssd1 vccd1 vccd1 _4814_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4743_ _5838_/A _4738_/X _4739_/X _4742_/X vssd1 vssd1 vccd1 vccd1 _4743_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3827__A _6116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5518__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4674_ _4703_/A _4674_/B vssd1 vssd1 vccd1 vccd1 _4677_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3625_ _6070_/Q _6072_/Q vssd1 vssd1 vccd1 vccd1 _5024_/B sky130_fd_sc_hd__and2b_2
XFILLER_0_101_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout105_A _5424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3556_ _3556_/A _3709_/B vssd1 vssd1 vccd1 vccd1 _3556_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_24_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5761__B _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5226_ _3540_/A _5218_/X _5220_/Y hold517/X vssd1 vssd1 vccd1 vccd1 _5226_/X sky130_fd_sc_hd__a22o_1
X_3487_ _4485_/B _4618_/C vssd1 vssd1 vccd1 vccd1 _4614_/D sky130_fd_sc_hd__nand2_1
X_5157_ _5157_/A _5157_/B vssd1 vssd1 vccd1 vccd1 _5157_/X sky130_fd_sc_hd__or2_1
XFILLER_0_98_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5088_ _5129_/A vssd1 vssd1 vccd1 vccd1 _5088_/Y sky130_fd_sc_hd__inv_2
X_4108_ hold86/X _3668_/X _4115_/S vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__mux2_1
XANTENNA__5489__A _6165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4039_ _5489_/B _4614_/B vssd1 vssd1 vccd1 vccd1 _4040_/B sky130_fd_sc_hd__and2_1
XANTENNA__6193__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5737__A2 _4879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4945__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4332__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3175__C _3488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5189__B1 _5186_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5728__A2 _4836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4400__A2 _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3647__A _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold308 _5241_/X vssd1 vssd1 vccd1 vccd1 _6132_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold319 _6093_/Q vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3410_ _4038_/A _3237_/Y _3324_/A vssd1 vssd1 vccd1 vccd1 _3410_/Y sky130_fd_sc_hd__a21oi_1
X_4390_ _4390_/A _4406_/A vssd1 vssd1 vccd1 vccd1 _4392_/A sky130_fd_sc_hd__nor2_1
X_3341_ _3343_/B _3344_/S vssd1 vssd1 vccd1 vccd1 _3341_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5073__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4478__A _4478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__B1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6060_ _6060_/CLK _6060_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6060_/Q sky130_fd_sc_hd__dfrtp_4
X_3272_ _3272_/A _3272_/B vssd1 vssd1 vccd1 vccd1 _4104_/B sky130_fd_sc_hd__nor2_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _5007_/B _5010_/X _5011_/S vssd1 vssd1 vccd1 vccd1 _5011_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3675__B1 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3690__A3 _6114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5102__A _5185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5913_ _6152_/CLK hold59/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dfxtp_1
X_5844_ _6114_/Q _5843_/X _5869_/S vssd1 vssd1 vccd1 vccd1 _5845_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_29_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5775_ _6237_/Q hold492/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5775_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_2987_ _6158_/Q vssd1 vssd1 vccd1 vccd1 _4538_/B sky130_fd_sc_hd__inv_2
XFILLER_0_44_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4726_ _4726_/A _4726_/B _4726_/C _4726_/D vssd1 vssd1 vccd1 vccd1 _4727_/C sky130_fd_sc_hd__or4_1
X_4657_ _6215_/Q _4943_/B _4714_/S vssd1 vssd1 vccd1 vccd1 _4659_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3608_ _3573_/C _3986_/A2 _3584_/X _3585_/X _2965_/Y vssd1 vssd1 vccd1 vccd1 _3608_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_101_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4588_ _4587_/X _4586_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4879_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_12_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3539_ _3539_/A _3539_/B _4726_/D vssd1 vssd1 vccd1 vccd1 _3539_/Y sky130_fd_sc_hd__nand3_4
X_6258_ _6259_/CLK _6258_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6258_/Q sky130_fd_sc_hd__dfrtp_4
X_5209_ _5209_/A _5209_/B _5209_/C vssd1 vssd1 vccd1 vccd1 _5209_/X sky130_fd_sc_hd__or3_1
X_6189_ _6190_/CLK _6189_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6189_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4327__S _4327_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold601_A _6179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3467__A _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4449__A2 _3488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5621__S _5705_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__6044__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3409__B1 _3488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3424__A3 _3434_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3890_ _4250_/A _3890_/B vssd1 vssd1 vccd1 vccd1 _4135_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5068__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5031__C1 _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5560_ _5558_/X _5559_/Y _5670_/A vssd1 vssd1 vccd1 vccd1 _5560_/X sky130_fd_sc_hd__mux2_1
X_5491_ _6237_/Q hold412/X _5497_/S vssd1 vssd1 vccd1 vccd1 _5491_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_38_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6060_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4511_ _6206_/Q _4805_/B _4589_/S vssd1 vssd1 vccd1 vccd1 _4512_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_26_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold105 _4316_/X vssd1 vssd1 vccd1 vccd1 _5985_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4442_ _3715_/B _4412_/A _4056_/A _4412_/B _3715_/Y vssd1 vssd1 vccd1 vccd1 _4442_/X
+ sky130_fd_sc_hd__a311o_1
Xhold116 _5892_/Q vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _4227_/X vssd1 vssd1 vccd1 vccd1 _5925_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold127 _3416_/X vssd1 vssd1 vccd1 vccd1 _5903_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold149 _5981_/Q vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4373_ _3392_/A _4457_/B _3433_/X hold619/X vssd1 vssd1 vccd1 vccd1 _4373_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_95_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3324_ _3324_/A _3324_/B vssd1 vssd1 vccd1 vccd1 _4427_/B sky130_fd_sc_hd__nand2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6112_ _6144_/CLK _6112_/D vssd1 vssd1 vccd1 vccd1 _6112_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__5637__A1 _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6043_ _6175_/CLK _6043_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6043_/Q sky130_fd_sc_hd__dfrtp_1
X_3255_ _3396_/A _3246_/A _3254_/Y _3395_/B _3251_/X vssd1 vssd1 vccd1 vccd1 _3255_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5531__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3186_ _4417_/A _3187_/B vssd1 vssd1 vccd1 vccd1 _4483_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout172_A input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5767__A _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3415__A3 _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5827_ hold595/X _5826_/X _5832_/S vssd1 vssd1 vccd1 vccd1 _6242_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3287__A _4043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5758_ _4119_/A _4976_/B _4691_/Y _5762_/C vssd1 vssd1 vccd1 vccd1 _5758_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3179__A2 _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4709_ _6160_/Q _4620_/Y _4708_/X vssd1 vssd1 vccd1 vccd1 _4709_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5689_ _5690_/A _5690_/B vssd1 vssd1 vccd1 vccd1 _5691_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4128__A1 _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4679__A2 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5876__A1 _5341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold650 _5350_/X vssd1 vssd1 vccd1 vccd1 _6172_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 _6042_/Q vssd1 vssd1 vccd1 vccd1 hold661/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5007__A _5007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold384_A _6119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold649_A _6172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4064__B1 _3694_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4520__S _4598_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5867__B2 _5245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5619__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4827__C1 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5095__A2 _4391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3040_ _3777_/A _5356_/A vssd1 vssd1 vccd1 vccd1 _3643_/B sky130_fd_sc_hd__or2_2
XANTENNA__4475__B _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4991_ _6242_/Q _5008_/B vssd1 vssd1 vccd1 vccd1 _4991_/X sky130_fd_sc_hd__and2_1
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3942_ _6141_/Q _4007_/S vssd1 vssd1 vccd1 vccd1 _3944_/B sky130_fd_sc_hd__xnor2_1
X_3873_ _3873_/A _3873_/B _3873_/C vssd1 vssd1 vccd1 vccd1 _3875_/B sky130_fd_sc_hd__or3_2
XFILLER_0_18_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5612_ _5602_/A _5611_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _5612_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5555__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3538__C _4726_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5543_ _4119_/B _5542_/X _4805_/Y vssd1 vssd1 vccd1 vccd1 _5543_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__5307__A0 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_15_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5858__A1 _3864_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5474_ _6155_/Q _6154_/Q _5474_/C _5474_/D vssd1 vssd1 vccd1 vccd1 _5474_/X sky130_fd_sc_hd__or4_1
X_4425_ _3643_/B _4614_/B _3167_/B _4484_/A vssd1 vssd1 vccd1 vccd1 _4427_/C sky130_fd_sc_hd__a211o_1
X_4356_ _4150_/X hold151/X _4363_/S vssd1 vssd1 vccd1 vccd1 _4356_/X sky130_fd_sc_hd__mux2_1
X_3307_ _3307_/A _3307_/B vssd1 vssd1 vccd1 vccd1 _3307_/Y sky130_fd_sc_hd__nor2_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4287_ _4193_/X hold275/X _4291_/S vssd1 vssd1 vccd1 vccd1 _4287_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5086__A2 _5107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ _6034_/CLK _6026_/D vssd1 vssd1 vccd1 vccd1 _6026_/Q sky130_fd_sc_hd__dfxtp_1
X_3238_ _3694_/C _3643_/B vssd1 vssd1 vccd1 vccd1 _3238_/Y sky130_fd_sc_hd__nor2_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3169_ _4486_/A _3192_/B vssd1 vssd1 vccd1 vccd1 _4439_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_55_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout55 _3346_/Y vssd1 vssd1 vccd1 vccd1 _5705_/S sky130_fd_sc_hd__buf_6
XFILLER_0_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout99 _4765_/Y vssd1 vssd1 vccd1 vccd1 _5701_/S sky130_fd_sc_hd__buf_4
XFILLER_0_64_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout88 _4116_/Y vssd1 vssd1 vccd1 vccd1 _4119_/A sky130_fd_sc_hd__buf_4
XFILLER_0_36_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout77 _3717_/X vssd1 vssd1 vccd1 vccd1 _4234_/A sky130_fd_sc_hd__clkbuf_8
Xfanout66 _5711_/X vssd1 vssd1 vccd1 vccd1 _5762_/C sky130_fd_sc_hd__buf_4
XANTENNA_hold599_A _6239_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4340__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold480 _6065_/Q vssd1 vssd1 vccd1 vccd1 hold480/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold491 _5684_/X vssd1 vssd1 vccd1 vccd1 _6201_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5077__A2 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4726__D _4726_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3245__D1 _4451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4683__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4210_ hold234/X hold68/X hold171/X hold70/X _5182_/S _5200_/B1 vssd1 vssd1 vccd1
+ vccd1 _4210_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5190_ _6159_/Q _5121_/Y _5187_/X _5189_/X vssd1 vssd1 vccd1 vccd1 _5190_/X sky130_fd_sc_hd__a211o_1
X_4141_ hold270/X _4292_/B _4364_/A hold122/X _4140_/X vssd1 vssd1 vccd1 vccd1 _4142_/B
+ sky130_fd_sc_hd__o221a_1
X_4072_ _4460_/A _4069_/X _4071_/X _4415_/A _4094_/D vssd1 vssd1 vccd1 vccd1 _4072_/X
+ sky130_fd_sc_hd__a32o_1
X_3023_ _4728_/A _3484_/A _3488_/A vssd1 vssd1 vccd1 vccd1 _4426_/A sky130_fd_sc_hd__or3_1
XANTENNA__5776__A0 _6238_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4974_ _4973_/X _6158_/Q _5704_/S vssd1 vssd1 vccd1 vccd1 _4974_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3925_ _6159_/Q _3924_/X _6074_/Q vssd1 vssd1 vccd1 vccd1 _3925_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3251__A1 _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5764__B _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3856_ _5024_/A _3899_/A vssd1 vssd1 vccd1 vccd1 _3856_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3787_ _3597_/X _3758_/Y _3759_/X _3786_/Y vssd1 vssd1 vccd1 vccd1 _3787_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4751__A1 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5526_ _5526_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5527_/B sky130_fd_sc_hd__and2_1
X_5457_ _5457_/A _5457_/B _5457_/C vssd1 vssd1 vccd1 vccd1 _5457_/X sky130_fd_sc_hd__or3_1
XANTENNA__4503__A1 input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4408_ _4391_/B _4054_/X _4749_/A vssd1 vssd1 vccd1 vccd1 _4408_/X sky130_fd_sc_hd__a21o_1
X_5388_ _5388_/A _5388_/B vssd1 vssd1 vccd1 vccd1 _5389_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4339_ hold208/X _3737_/X _4345_/S vssd1 vssd1 vccd1 vccd1 _6005_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6009_ _6029_/CLK _6009_/D vssd1 vssd1 vccd1 vccd1 _6009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3490__A1 _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4335__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3242__A1 _6174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4742__A1 _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5207__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4430__B1 _4446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3710_ _5093_/A _3246_/A _3246_/B _3543_/Y _3709_/Y vssd1 vssd1 vccd1 vccd1 _3710_/X
+ sky130_fd_sc_hd__o311a_1
X_4690_ _4677_/A _4677_/B _4703_/A vssd1 vssd1 vccd1 vccd1 _4691_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3641_ _3635_/X _3636_/Y _3848_/B _3640_/X vssd1 vssd1 vccd1 vccd1 _3641_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3385__A _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3572_ _3513_/A _3571_/X _4963_/A vssd1 vssd1 vccd1 vccd1 _3573_/C sky130_fd_sc_hd__a21oi_4
X_5311_ input6/X hold635/X _5313_/S vssd1 vssd1 vccd1 vccd1 _6159_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_51_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5242_ _6134_/D _6134_/Q vssd1 vssd1 vccd1 vccd1 _5242_/X sky130_fd_sc_hd__and2b_1
XANTENNA__4497__A0 _6205_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5173_ _3879_/X _4210_/X _5169_/X _5172_/X _5185_/S _5116_/A vssd1 vssd1 vccd1 vccd1
+ _5173_/X sky130_fd_sc_hd__mux4_2
XANTENNA__5105__A _5120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4124_ _4124_/A _4124_/B _4446_/A _5424_/B vssd1 vssd1 vccd1 vccd1 _4124_/X sky130_fd_sc_hd__or4_1
Xinput1 io_in[24] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4944__A _6239_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4055_ _3694_/C _4054_/X _4053_/X vssd1 vssd1 vccd1 vccd1 _4055_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5461__A2 _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3006_ _6259_/Q _6258_/Q vssd1 vssd1 vccd1 vccd1 _4486_/A sky130_fd_sc_hd__nand2_8
XANTENNA__3472__B2 _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4957_ _4956_/X _6157_/Q _5704_/S vssd1 vssd1 vccd1 vccd1 _4957_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4421__B1 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3908_ _6172_/Q _3909_/B vssd1 vssd1 vccd1 vccd1 _4014_/A sky130_fd_sc_hd__nor2_1
X_4888_ _6161_/Q _5008_/B _4881_/X _4999_/A1 _4887_/X vssd1 vssd1 vccd1 vccd1 _4888_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3839_ _6173_/Q _3699_/Y _3912_/C _3838_/Y vssd1 vssd1 vccd1 vccd1 _3840_/B sky130_fd_sc_hd__o22a_1
XANTENNA__4724__A1 _5164_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5509_ _2957_/Y _3370_/B _5220_/A vssd1 vssd1 vccd1 vccd1 _5509_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold631_A _6156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4638__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4191__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3933__A _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5140__A1 _5164_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3151__B1 _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4764__A _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5443__A2 _5343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5860_ _6136_/Q _6114_/Q _5868_/S vssd1 vssd1 vccd1 vccd1 _5860_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_75_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4811_ _4805_/B _4810_/X _4963_/A vssd1 vssd1 vccd1 vccd1 _4811_/X sky130_fd_sc_hd__mux2_1
X_5791_ _5762_/A _5352_/A _5773_/B vssd1 vssd1 vccd1 vccd1 _5791_/X sky130_fd_sc_hd__o21a_2
XFILLER_0_28_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4742_ _4415_/A _4732_/X _4741_/X _4118_/A vssd1 vssd1 vccd1 vccd1 _4742_/X sky130_fd_sc_hd__a22o_1
X_4673_ _4699_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _4674_/B sky130_fd_sc_hd__or2_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3624_ _6073_/Q _5460_/S vssd1 vssd1 vccd1 vccd1 _3624_/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_98_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4706__B2 _4474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4182__A2 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3265__D _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3555_ _5362_/B _5424_/C _3554_/X vssd1 vssd1 vccd1 vccd1 _3555_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5534__S _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3486_ _4772_/C _4483_/A _4483_/B vssd1 vssd1 vccd1 vccd1 _4613_/C sky130_fd_sc_hd__or3_1
XANTENNA__5131__A1 _6205_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5225_ _6076_/Q _5225_/B vssd1 vssd1 vccd1 vccd1 _5225_/X sky130_fd_sc_hd__and2b_1
XANTENNA__5131__B2 _6189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5156_ _5895_/Q _3591_/A _3739_/S _6007_/Q _5179_/S vssd1 vssd1 vccd1 vccd1 _5157_/B
+ sky130_fd_sc_hd__o221a_1
X_5087_ _5107_/A _5107_/B vssd1 vssd1 vccd1 vccd1 _5129_/A sky130_fd_sc_hd__or2_2
X_4107_ _5297_/A _4263_/A vssd1 vssd1 vccd1 vccd1 _4115_/S sky130_fd_sc_hd__nor2_4
X_4038_ _4038_/A _4038_/B _4070_/B vssd1 vssd1 vccd1 vccd1 _4416_/A sky130_fd_sc_hd__and3_1
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5989_ _6144_/CLK _5989_/D vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__4945__B2 _4943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3381__B1 _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4556__S0 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4881__A0 _4879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3987__A2 _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4759__A _4759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold309 _6080_/Q vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__dlygate4sd3_1
X_3340_ _3343_/B _3344_/S vssd1 vssd1 vccd1 vccd1 _3340_/X sky130_fd_sc_hd__and2b_1
XANTENNA__3382__B _3383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _6203_/Q _6069_/Q _6038_/Q vssd1 vssd1 vccd1 vccd1 _5010_/X sky130_fd_sc_hd__mux2_1
X_3271_ _4124_/B _3205_/B _4999_/A1 vssd1 vssd1 vccd1 vccd1 _3275_/A sky130_fd_sc_hd__a21o_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3427__A1 _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5912_ _6010_/CLK _5912_/D vssd1 vssd1 vccd1 vccd1 _5912_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5843_ _6118_/Q _6136_/Q _5868_/S vssd1 vssd1 vccd1 vccd1 _5843_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3838__A _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4388__C1 _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5774_ _6236_/Q hold441/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5774_/X sky130_fd_sc_hd__mux2_1
X_2986_ _6156_/Q vssd1 vssd1 vccd1 vccd1 _4507_/B sky130_fd_sc_hd__inv_2
XFILLER_0_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4725_ _4739_/A _4725_/B vssd1 vssd1 vccd1 vccd1 _4725_/X sky130_fd_sc_hd__or2_1
X_4656_ _4655_/X _4654_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4943_/B sky130_fd_sc_hd__mux2_2
XANTENNA__3276__C _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3607_ hold189/X hold217/X _3724_/S vssd1 vssd1 vccd1 vccd1 _3607_/X sky130_fd_sc_hd__mux2_1
X_4587_ hold106/X hold168/X _6003_/Q _5964_/Q _5076_/A0 _4272_/B vssd1 vssd1 vccd1
+ vccd1 _4587_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_101_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5264__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3538_ _3539_/A _6166_/Q _4726_/D vssd1 vssd1 vccd1 vccd1 _3573_/B sky130_fd_sc_hd__and3_2
XANTENNA__3573__A _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3469_ _4445_/B _4759_/A vssd1 vssd1 vccd1 vccd1 _3469_/Y sky130_fd_sc_hd__nor2_2
X_6257_ _6259_/CLK _6257_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6257_/Q sky130_fd_sc_hd__dfrtp_1
X_5208_ _5899_/Q _3591_/A _3739_/S _6011_/Q _5179_/S vssd1 vssd1 vccd1 vccd1 _5209_/C
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3666__A1 _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6188_ _6190_/CLK _6188_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6188_/Q sky130_fd_sc_hd__dfrtp_4
X_5139_ _5139_/A _5139_/B vssd1 vssd1 vccd1 vccd1 _5139_/X sky130_fd_sc_hd__or2_1
XFILLER_0_79_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6208_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3418__A1 _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4091__B2 _5220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4343__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3748__A _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3467__B _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4518__S _4596_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3409__A1 _6048_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4082__A1 _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4909__A1 _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5873__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5490_ _6236_/Q hold371/X _5497_/S vssd1 vssd1 vccd1 vccd1 _5490_/X sky130_fd_sc_hd__mux2_1
X_4510_ _4509_/X _4508_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4805_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold117 _3669_/X vssd1 vssd1 vccd1 vccd1 _5892_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ _3654_/S _4731_/S _4440_/X vssd1 vssd1 vccd1 vccd1 _4441_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_41_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold106 _5987_/Q vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 _5960_/Q vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 _5982_/Q vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4372_ hold242/X _4261_/X _4372_/S vssd1 vssd1 vccd1 vccd1 _4372_/X sky130_fd_sc_hd__mux2_1
X_6111_ _6111_/CLK hold26/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3323_ _4398_/A _4051_/B _3323_/C vssd1 vssd1 vccd1 vccd1 _3324_/B sky130_fd_sc_hd__or3_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5637__A2 _6197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6042_ _6119_/CLK _6042_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6042_/Q sky130_fd_sc_hd__dfrtp_1
X_3254_ _3543_/B _5498_/B vssd1 vssd1 vccd1 vccd1 _3254_/Y sky130_fd_sc_hd__nand2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3185_ _3543_/A _4385_/A _3185_/C vssd1 vssd1 vccd1 vccd1 _3200_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_95_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5847__A1_N _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_44_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4073__B2 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5826_ _5825_/X _3959_/Y _5831_/S vssd1 vssd1 vccd1 vccd1 _5826_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5757_ hold565/X _5741_/Y _5756_/X _5767_/A vssd1 vssd1 vccd1 vccd1 _5757_/X sky130_fd_sc_hd__o22a_1
X_2969_ _6171_/Q vssd1 vssd1 vccd1 vccd1 _2969_/Y sky130_fd_sc_hd__inv_2
X_4708_ _5764_/B _4706_/X _4707_/X vssd1 vssd1 vccd1 vccd1 _4708_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4781__C1 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3584__B1 _3671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5688_ _5682_/B _5682_/C _5678_/Y vssd1 vssd1 vccd1 vccd1 _5690_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_71_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4128__A2 _5330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4639_ _6022_/Q _5967_/Q _6014_/Q _5947_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4639_/X sky130_fd_sc_hd__mux4_1
Xhold651 _6173_/Q vssd1 vssd1 vccd1 vccd1 hold651/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3887__A1 _3795_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold640 _6253_/Q vssd1 vssd1 vccd1 vccd1 hold640/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout78_A _3717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4338__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5023__A _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold544_A _6197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5677__B _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5013__A0 _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5564__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5867__A2 _5836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3644__C _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4827__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4772__A _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4055__A1 _3694_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4990_ _4990_/A _4990_/B vssd1 vssd1 vccd1 vccd1 _4990_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3941_ _5024_/A _6141_/Q _6119_/Q _3848_/B _3940_/X vssd1 vssd1 vccd1 vccd1 _5372_/A
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3872_ _3795_/C _3869_/X _3871_/X vssd1 vssd1 vccd1 vccd1 _3873_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5611_ _5610_/X _5605_/X _5670_/A vssd1 vssd1 vccd1 vccd1 _5611_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5542_ _5541_/X _6056_/Q _5595_/S vssd1 vssd1 vccd1 vccd1 _5542_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5473_ _6157_/Q _6156_/Q _6161_/Q _6160_/Q vssd1 vssd1 vccd1 vccd1 _5474_/D sky130_fd_sc_hd__or4_1
XFILLER_0_1_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4424_ _5502_/B _4727_/B _4729_/A _4424_/D vssd1 vssd1 vccd1 vccd1 _5338_/B sky130_fd_sc_hd__or4_1
X_4355_ _4355_/A _4364_/B vssd1 vssd1 vccd1 vccd1 _4363_/S sky130_fd_sc_hd__or2_4
X_3306_ _3306_/A _4445_/B _3306_/C vssd1 vssd1 vccd1 vccd1 _3307_/B sky130_fd_sc_hd__and3_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _4180_/X hold224/X _4291_/S vssd1 vssd1 vccd1 vccd1 _5947_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5086__A3 _5085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5491__A0 _6237_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6025_ _6035_/CLK _6025_/D vssd1 vssd1 vccd1 vccd1 _6025_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _3654_/S _3237_/B vssd1 vssd1 vccd1 vccd1 _3237_/Y sky130_fd_sc_hd__xnor2_4
X_3168_ _3477_/A _4460_/C _3168_/C _3479_/A vssd1 vssd1 vccd1 vccd1 _3281_/A sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_0_wb_clk_i_A _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3099_ _4094_/D _3654_/S vssd1 vssd1 vccd1 vccd1 _3203_/D sky130_fd_sc_hd__nand2_2
XFILLER_0_76_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xci2406_z80_190 vssd1 vssd1 vccd1 vccd1 ci2406_z80_190/HI io_oeb[5] sky130_fd_sc_hd__conb_1
XFILLER_0_91_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5809_ _6239_/Q _5791_/X _5808_/X _5764_/B vssd1 vssd1 vccd1 vccd1 _5809_/X sky130_fd_sc_hd__a22o_1
Xfanout78 _3717_/X vssd1 vssd1 vccd1 vccd1 _4219_/A sky130_fd_sc_hd__buf_2
XFILLER_0_64_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout89 _3539_/Y vssd1 vssd1 vccd1 vccd1 _4253_/A2 sky130_fd_sc_hd__clkbuf_8
Xfanout67 _4926_/S vssd1 vssd1 vccd1 vccd1 _5609_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__5546__A1 _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold494_A _6046_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold481 _4667_/X vssd1 vssd1 vccd1 vccd1 _6065_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold470 _6206_/Q vssd1 vssd1 vccd1 vccd1 hold470/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 _6221_/Q vssd1 vssd1 vccd1 vccd1 hold492/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4037__A1 _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5170__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4140_ _5920_/Q _4132_/A _4346_/A _6012_/Q vssd1 vssd1 vccd1 vccd1 _4140_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4486__B _4486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3079__A2 _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4071_ _4061_/A _4061_/C _4070_/Y _4056_/A vssd1 vssd1 vccd1 vccd1 _4071_/X sky130_fd_sc_hd__a31o_1
X_3022_ _4737_/A _3022_/B vssd1 vssd1 vccd1 vccd1 _4726_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ _5694_/A _4972_/X _4959_/Y vssd1 vssd1 vccd1 vccd1 _4973_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_58_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3924_ _3624_/Y _5373_/B _3918_/X _3923_/X vssd1 vssd1 vccd1 vccd1 _3924_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5528__A1 _6189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3855_ _3855_/A _5448_/A vssd1 vssd1 vccd1 vccd1 _3899_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3786_ _3597_/X _3785_/A _4253_/A2 vssd1 vssd1 vccd1 vccd1 _3786_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_22_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6206_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5525_ _5526_/A _5526_/B vssd1 vssd1 vccd1 vccd1 _5540_/B sky130_fd_sc_hd__nor2_1
X_5456_ _6177_/Q _5352_/Y _5354_/B _2990_/Y vssd1 vssd1 vccd1 vccd1 _5457_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4407_ _5502_/B _4391_/B _4043_/C _4406_/Y _3477_/C vssd1 vssd1 vccd1 vccd1 _4407_/X
+ sky130_fd_sc_hd__a32o_1
X_5387_ _5387_/A _5387_/B vssd1 vssd1 vccd1 vccd1 _5388_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4338_ hold130/X _3668_/X _4345_/S vssd1 vssd1 vccd1 vccd1 _4338_/X sky130_fd_sc_hd__mux2_1
X_4269_ hold175/X _4226_/X _4271_/S vssd1 vssd1 vccd1 vccd1 _4269_/X sky130_fd_sc_hd__mux2_1
X_6008_ _6029_/CLK _6008_/D vssd1 vssd1 vccd1 vccd1 _6008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4351__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5182__S _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5207__B1 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5758__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5758__A1 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4430__B2 _3193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4430__A1 _3488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3640_ _5024_/B _3628_/X _3636_/A _3639_/X vssd1 vssd1 vccd1 vccd1 _3640_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3385__B _4486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4733__A2 _4433_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3571_ _3457_/A _3560_/X _3565_/X _3567_/Y vssd1 vssd1 vccd1 vccd1 _3571_/X sky130_fd_sc_hd__a211o_2
X_5310_ input5/X hold629/X _5313_/S vssd1 vssd1 vccd1 vccd1 _6158_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5143__C1 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5241_ hold307/X _5107_/A _5875_/A vssd1 vssd1 vccd1 vccd1 _5241_/X sky130_fd_sc_hd__mux2_1
X_5172_ _5172_/A _5172_/B vssd1 vssd1 vccd1 vccd1 _5172_/X sky130_fd_sc_hd__or2_1
XANTENNA__5105__B _5105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4123_ _4697_/S _4122_/X _5296_/S vssd1 vssd1 vccd1 vccd1 _5914_/D sky130_fd_sc_hd__mux2_1
Xinput2 io_in[25] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_2
X_4054_ _4737_/A _4618_/A _4054_/C vssd1 vssd1 vccd1 vccd1 _4054_/X sky130_fd_sc_hd__and3_1
XANTENNA__4944__B _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3005_ _6259_/Q _6258_/Q vssd1 vssd1 vccd1 vccd1 _4038_/B sky130_fd_sc_hd__and2_1
XANTENNA__5749__B2 _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5749__A1 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4960__A _6240_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4956_ _5694_/A _4955_/X _4943_/Y vssd1 vssd1 vccd1 vccd1 _4956_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4972__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3907_ _6140_/Q _6141_/Q _3906_/B _5046_/A vssd1 vssd1 vccd1 vccd1 _3909_/B sky130_fd_sc_hd__o31a_1
X_4887_ _4776_/Y _4901_/B _4882_/X _4824_/B vssd1 vssd1 vccd1 vccd1 _4887_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3838_ _6173_/Q _6176_/Q vssd1 vssd1 vccd1 vccd1 _3838_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_46_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4185__B1 _3615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3769_ _3647_/C _3767_/Y _3768_/X vssd1 vssd1 vccd1 vccd1 _3769_/X sky130_fd_sc_hd__o21ba_1
X_5508_ _5507_/A _5507_/B hold52/X vssd1 vssd1 vccd1 vccd1 _5508_/X sky130_fd_sc_hd__a21o_2
X_5439_ _5437_/X _5438_/X _5363_/C _5435_/X vssd1 vssd1 vccd1 vccd1 _5439_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_0_69_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout60_A _4763_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5685__B _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3652__C _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5428__B1 _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5243__B1_N _3252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4764__B _6050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4256__S _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4651__A1 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4810_ _6190_/Q _6056_/Q _6038_/Q vssd1 vssd1 vccd1 vccd1 _4810_/X sky130_fd_sc_hd__mux2_1
X_5790_ _5327_/B _5790_/B _5790_/C _5790_/D vssd1 vssd1 vccd1 vccd1 _5831_/S sky130_fd_sc_hd__and4b_4
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4741_ _3203_/B _4483_/A _4740_/X _4739_/A _3334_/B vssd1 vssd1 vccd1 vccd1 _4741_/X
+ sky130_fd_sc_hd__a221o_1
X_4672_ _4699_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _4703_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4706__A2 _4612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3623_ _6073_/Q _5460_/S vssd1 vssd1 vccd1 vccd1 _3623_/X sky130_fd_sc_hd__and2_1
XFILLER_0_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3554_ _3554_/A _4046_/B vssd1 vssd1 vccd1 vccd1 _3554_/X sky130_fd_sc_hd__or2_1
X_3485_ _4613_/B vssd1 vssd1 vccd1 vccd1 _3485_/Y sky130_fd_sc_hd__inv_2
XANTENNA__5116__A _5116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5224_ _5217_/Y _5223_/X _3540_/A _3353_/B vssd1 vssd1 vccd1 vccd1 _6124_/D sky130_fd_sc_hd__a2bb2o_1
X_5155_ _5999_/Q _3591_/A _3740_/S _5960_/Q _4256_/S vssd1 vssd1 vccd1 vccd1 _5157_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5086_ _5120_/A _5107_/A _5085_/B _5023_/A vssd1 vssd1 vccd1 vccd1 _5086_/Y sky130_fd_sc_hd__a31oi_4
X_4106_ hold367/X _4105_/X _5296_/S vssd1 vssd1 vccd1 vccd1 _4106_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_79_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4037_ _3210_/C _3622_/C _4053_/A _4118_/A vssd1 vssd1 vccd1 vccd1 _4037_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5988_ _6151_/CLK _5988_/D vssd1 vssd1 vccd1 vccd1 _5988_/Q sky130_fd_sc_hd__dfxtp_1
X_4939_ _4990_/A _4938_/Y _4928_/Y vssd1 vssd1 vccd1 vccd1 _4939_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_93_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3381__A1 _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4556__S1 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4865__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4633__B2 _4474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xmax_cap97 _3488_/A vssd1 vssd1 vccd1 vccd1 _3395_/B sky130_fd_sc_hd__buf_2
Xmax_cap75 _3577_/S vssd1 vssd1 vccd1 vccd1 _3986_/A2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4804__S _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4936__A2 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4149__B1 _3671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4759__B _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3270_ _4771_/A _4771_/B _4771_/C vssd1 vssd1 vccd1 vccd1 _3270_/X sky130_fd_sc_hd__and3b_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4872__A1 _6160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3675__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4872__B2 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_34_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_88_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5911_ _6029_/CLK hold99/X vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__3427__A2 _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5842_ hold336/X _5836_/A _5841_/X _5773_/A vssd1 vssd1 vccd1 vccd1 _5842_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5773_ _5773_/A _5773_/B vssd1 vssd1 vccd1 vccd1 _5789_/S sky130_fd_sc_hd__or2_4
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3838__B _6176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2985_ _6157_/Q vssd1 vssd1 vccd1 vccd1 _4522_/B sky130_fd_sc_hd__inv_2
XFILLER_0_56_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4724_ _5164_/A1 _6070_/Q _4927_/S _4450_/X vssd1 vssd1 vccd1 vccd1 _4724_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_71_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4655_ _6023_/Q _5968_/Q _6015_/Q _5948_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4655_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_71_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3276__D _4439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3606_ _3968_/A _3616_/B _3793_/D vssd1 vssd1 vccd1 vccd1 _4292_/B sky130_fd_sc_hd__or3_1
X_4586_ hold76/X hold58/X hold118/X hold227/X _5076_/A0 _4272_/B vssd1 vssd1 vccd1
+ vccd1 _4586_/X sky130_fd_sc_hd__mux4_1
XANTENNA_fanout110_A _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3537_ _4460_/A _4497_/S _4726_/D vssd1 vssd1 vccd1 vccd1 _3671_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_58_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6256_ _6256_/CLK _6256_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6256_/Q sky130_fd_sc_hd__dfrtp_1
X_3468_ _5362_/B _3713_/A _3543_/B _4390_/A _4765_/A vssd1 vssd1 vccd1 vccd1 _3468_/X
+ sky130_fd_sc_hd__a2111o_1
X_6187_ _6242_/CLK _6187_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6187_/Q sky130_fd_sc_hd__dfrtp_1
X_3399_ _3405_/B _3399_/B vssd1 vssd1 vccd1 vccd1 _3399_/X sky130_fd_sc_hd__or2_1
X_5207_ _6003_/Q _3591_/A _3740_/S _5964_/Q _4256_/S vssd1 vssd1 vccd1 vccd1 _5209_/B
+ sky130_fd_sc_hd__o221a_1
X_5138_ _6197_/Q _5119_/Y _5121_/Y _6155_/Q _5137_/X vssd1 vssd1 vccd1 vccd1 _5139_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_98_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5069_ hold15/X _4173_/B _5073_/S vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__mux2_1
XANTENNA__3418__A2 _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5040__A1 _6116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5040__B2 _6114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3764__A _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3339__D1 _6130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5500__C1 _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4534__S _4596_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5031__A1 _2960_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6053__RESET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4440_ _3277_/A _4070_/B _4731_/S _4439_/X _3421_/Y vssd1 vssd1 vccd1 vccd1 _4440_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold107 _4318_/X vssd1 vssd1 vccd1 vccd1 _5987_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 _5899_/Q vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 _4313_/X vssd1 vssd1 vccd1 vccd1 _5982_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4371_ hold225/X _4242_/X _4372_/S vssd1 vssd1 vccd1 vccd1 _4371_/X sky130_fd_sc_hd__mux2_1
X_6110_ _6110_/CLK hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3322_ _3319_/Y _3320_/Y _3321_/X _4077_/A vssd1 vssd1 vccd1 vccd1 _3343_/B sky130_fd_sc_hd__a31o_1
XFILLER_0_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ _6119_/CLK _6041_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6041_/Q sky130_fd_sc_hd__dfrtp_1
X_3253_ _5498_/B vssd1 vssd1 vccd1 vccd1 _3328_/B sky130_fd_sc_hd__inv_2
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _3184_/A _3411_/D vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__or2_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_47_wb_clk_i _5978_/CLK vssd1 vssd1 vccd1 vccd1 _6190_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__5270__A1 _6157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5270__B2 _6239_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5825_ hold332/X _5794_/Y _5824_/X _5794_/B vssd1 vssd1 vccd1 vccd1 _5825_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout158_A _5245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5756_ _3864_/Y _5771_/S _5742_/Y _5755_/X vssd1 vssd1 vccd1 vccd1 _5756_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_44_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2968_ _3405_/B vssd1 vssd1 vccd1 vccd1 _2968_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5687_ _5687_/A _5687_/B vssd1 vssd1 vccd1 vccd1 _5690_/A sky130_fd_sc_hd__or2_1
X_4707_ hold423/X _5762_/A _4619_/X vssd1 vssd1 vccd1 vccd1 _4707_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4781__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4638_ hold66/A hold54/A _5922_/Q _6030_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4638_/X sky130_fd_sc_hd__mux4_1
Xhold630 _6160_/Q vssd1 vssd1 vccd1 vccd1 hold630/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3336__A1 _3302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4569_ hold559/X _4568_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _4569_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold652 _6130_/Q vssd1 vssd1 vccd1 vccd1 hold652/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold641 _5879_/X vssd1 vssd1 vccd1 vccd1 _6253_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5089__A1 _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6239_ _6243_/CLK _6239_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6239_/Q sky130_fd_sc_hd__dfstp_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4354__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5261__A1 _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5261__B2 _6237_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4695__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3575__A1 _3513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5185__S _5185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3878__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4264__S _4271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3940_ _3639_/X _3935_/Y _3939_/X _5024_/B _3938_/X vssd1 vssd1 vccd1 vccd1 _3940_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3263__B1 _5424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3871_ _3582_/Y _3870_/X _3968_/A vssd1 vssd1 vccd1 vccd1 _3871_/X sky130_fd_sc_hd__o21a_1
XANTENNA__5884__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5610_ _5609_/X _5602_/A _5705_/S vssd1 vssd1 vccd1 vccd1 _5610_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_45_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3566__A1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5541_ _6190_/Q _5606_/S _4806_/X vssd1 vssd1 vccd1 vccd1 _5541_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_81_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5472_ _5050_/B _5330_/B _5471_/X vssd1 vssd1 vccd1 vccd1 _5472_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4423_ _4129_/B _4422_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _6044_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4354_ _4261_/X hold294/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4354_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3305_ _4433_/B _3713_/B _5838_/B _3286_/Y vssd1 vssd1 vccd1 vccd1 _3307_/A sky130_fd_sc_hd__a22o_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6024_ _6031_/CLK _6024_/D vssd1 vssd1 vccd1 vccd1 _6024_/Q sky130_fd_sc_hd__dfxtp_1
X_4285_ _4165_/X hold283/X _4291_/S vssd1 vssd1 vccd1 vccd1 _5946_/D sky130_fd_sc_hd__mux2_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4818__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _6178_/Q _6172_/Q _4739_/A vssd1 vssd1 vccd1 vccd1 _3237_/B sky130_fd_sc_hd__mux2_2
XANTENNA__4963__A _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3167_ _4728_/A _3167_/B vssd1 vssd1 vccd1 vccd1 _3479_/A sky130_fd_sc_hd__or2_2
X_3098_ _4485_/A _3125_/C vssd1 vssd1 vccd1 vccd1 _4433_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5794__A _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_191 vssd1 vssd1 vccd1 vccd1 ci2406_z80_191/HI io_oeb[6] sky130_fd_sc_hd__conb_1
X_5808_ hold488/X _5457_/A _5352_/Y _2989_/Y vssd1 vssd1 vccd1 vccd1 _5808_/X sky130_fd_sc_hd__a22o_1
Xfanout68 _4926_/S vssd1 vssd1 vccd1 vccd1 _5704_/S sky130_fd_sc_hd__clkbuf_8
Xfanout57 _4766_/Y vssd1 vssd1 vccd1 vccd1 _4815_/B sky130_fd_sc_hd__buf_4
Xfanout79 _3594_/Y vssd1 vssd1 vccd1 vccd1 _4256_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_91_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5739_ hold583/X _5714_/Y _5738_/X _5023_/A vssd1 vssd1 vccd1 vccd1 _5739_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_17_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4601__S0 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold471 _5724_/X vssd1 vssd1 vccd1 vccd1 _6206_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold460 _6195_/Q vssd1 vssd1 vccd1 vccd1 _5602_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold493 _5775_/X vssd1 vssd1 vccd1 vccd1 _6221_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4349__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold482 _6141_/Q vssd1 vssd1 vccd1 vccd1 hold482/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5034__A _6135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4668__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4745__B1 _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5209__A _5209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5846__A1_N _3707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3671__B _3671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4486__C _5424_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4070_ _4124_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _4070_/Y sky130_fd_sc_hd__nand2_1
X_3021_ _3426_/A _3135_/B _4417_/A _4051_/B vssd1 vssd1 vccd1 vccd1 _3488_/A sky130_fd_sc_hd__nor4_4
XANTENNA__3399__A _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4972_ _6066_/Q _5702_/A2 _5607_/B1 _4971_/X vssd1 vssd1 vccd1 vccd1 _4972_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_19_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3236__A0 _6178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3923_ _3921_/A _3645_/X _3922_/X _6118_/Q _3920_/X vssd1 vssd1 vccd1 vccd1 _3923_/X
+ sky130_fd_sc_hd__a221o_1
X_3854_ _3855_/A _5448_/A vssd1 vssd1 vccd1 vccd1 _3854_/X sky130_fd_sc_hd__or2_1
XFILLER_0_18_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5528__A2 _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3785_ _3785_/A vssd1 vssd1 vccd1 vccd1 _3785_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4200__A2 _3588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5524_ _5524_/A _5524_/B vssd1 vssd1 vccd1 vccd1 _5526_/B sky130_fd_sc_hd__xnor2_1
X_5455_ _2990_/Y _5317_/A _5454_/Y vssd1 vssd1 vccd1 vccd1 _5457_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4406_ _4406_/A _4446_/B vssd1 vssd1 vccd1 vccd1 _4406_/Y sky130_fd_sc_hd__nor2_1
X_5386_ _5386_/A _5386_/B vssd1 vssd1 vccd1 vccd1 _5388_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4337_ _5297_/A _4364_/A vssd1 vssd1 vccd1 vccd1 _4345_/S sky130_fd_sc_hd__nor2_4
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4268_ hold68/X _4211_/X _4271_/S vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__mux2_1
X_6007_ _6152_/CLK _6007_/D vssd1 vssd1 vccd1 vccd1 _6007_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3475__B1 _4446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3219_ _3268_/B _4770_/A vssd1 vssd1 vccd1 vccd1 _4771_/A sky130_fd_sc_hd__and2b_1
X_4199_ hold70/X _3611_/X _3613_/X hold68/X _4198_/X vssd1 vssd1 vccd1 vccd1 _4202_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3102__A _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3772__A _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold290 _6051_/Q vssd1 vssd1 vccd1 vccd1 _3272_/B sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4258__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5758__A2 _4976_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4430__A2 _4759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3570_ _3535_/X _3671_/B _3539_/Y _3569_/Y _5023_/A vssd1 vssd1 vccd1 vccd1 _5297_/A
+ sky130_fd_sc_hd__a41o_4
XANTENNA__4733__A3 _4759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5143__B1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5240_ _3591_/A _5239_/X _5296_/S vssd1 vssd1 vccd1 vccd1 _6131_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_11_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5171_ _5924_/Q _5200_/A2 _4255_/S _6032_/Q _5182_/S vssd1 vssd1 vccd1 vccd1 _5172_/B
+ sky130_fd_sc_hd__o221a_1
X_4122_ _2967_/A _4120_/Y _4121_/X _3272_/A vssd1 vssd1 vccd1 vccd1 _4122_/X sky130_fd_sc_hd__a22o_1
X_4053_ _4053_/A _4061_/D vssd1 vssd1 vccd1 vccd1 _4053_/X sky130_fd_sc_hd__and2_1
Xinput3 io_in[26] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
X_3004_ _5356_/A _3643_/A vssd1 vssd1 vccd1 vccd1 _3135_/B sky130_fd_sc_hd__or2_4
XFILLER_0_93_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4955_ _6065_/Q _5702_/A2 _5607_/B1 _4954_/X vssd1 vssd1 vccd1 vccd1 _4955_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4960__B _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3906_ _6140_/Q _3906_/B vssd1 vssd1 vccd1 vccd1 _3911_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5548__S _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4886_ _6211_/Q _5009_/A2 _4769_/Y _4879_/B _4815_/B vssd1 vssd1 vccd1 vccd1 _4886_/X
+ sky130_fd_sc_hd__a221o_1
X_3837_ hold222/X _3836_/X _4035_/S vssd1 vssd1 vccd1 vccd1 _3837_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3768_ _5024_/B _3763_/Y _3767_/A _3639_/X vssd1 vssd1 vccd1 vccd1 _3768_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_14_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5507_ _5507_/A _5507_/B vssd1 vssd1 vccd1 vccd1 _5507_/Y sky130_fd_sc_hd__nand2_4
X_3699_ _6136_/Q _6137_/Q _6138_/Q vssd1 vssd1 vccd1 vccd1 _3699_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5438_ _6175_/Q _5026_/A _5436_/X _5025_/A _5330_/B vssd1 vssd1 vccd1 vccd1 _5438_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5369_ _5368_/X _6170_/Q _5484_/S vssd1 vssd1 vccd1 vccd1 _5369_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout53_A _5020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4362__S _4363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5901__RESET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3384__C1 _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3923__B2 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5676__A1 _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5428__A1 _3785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4537__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4100__A1 _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_output34_A _6090_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3677__A _5209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4740_ _3488_/B _4759_/A _4125_/C _4429_/X vssd1 vssd1 vccd1 vccd1 _4740_/X sky130_fd_sc_hd__a211o_1
X_4671_ _6216_/Q _4963_/B _4714_/S vssd1 vssd1 vccd1 vccd1 _4673_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_71_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3622_ _4118_/A _4094_/B _3622_/C vssd1 vssd1 vccd1 vccd1 _3958_/S sky130_fd_sc_hd__and3_4
XFILLER_0_3_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3553_ _3457_/A _3551_/X _3549_/X vssd1 vssd1 vccd1 vccd1 _3559_/A sky130_fd_sc_hd__o21ai_2
X_3484_ _3484_/A _3488_/A _3488_/B vssd1 vssd1 vccd1 vccd1 _4613_/B sky130_fd_sc_hd__or3_1
XANTENNA__5667__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5223_ _4077_/A _5221_/X _5222_/Y _5218_/X vssd1 vssd1 vccd1 vccd1 _5223_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5154_ hold404/X _5104_/Y _5119_/Y _6199_/Q vssd1 vssd1 vccd1 vccd1 _5163_/C sky130_fd_sc_hd__a22o_1
X_4105_ _3272_/A _6053_/Q _4105_/S vssd1 vssd1 vccd1 vccd1 _4105_/X sky130_fd_sc_hd__mux2_1
X_5085_ _5107_/A _5085_/B vssd1 vssd1 vccd1 vccd1 _5122_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4036_ _4124_/A _4036_/B vssd1 vssd1 vccd1 vccd1 _4053_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5987_ _6102_/CLK _5987_/D vssd1 vssd1 vccd1 vccd1 _5987_/Q sky130_fd_sc_hd__dfxtp_1
X_4938_ _6064_/Q _5702_/A2 _5607_/B1 _4937_/X vssd1 vssd1 vccd1 vccd1 _4938_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4869_ _6060_/Q _4856_/A _4824_/B vssd1 vssd1 vccd1 vccd1 _4869_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_30 _5218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4910__S _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5202__S0 _5185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold567_A _6174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4865__B _4865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4357__S _4363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4633__A2 _4612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4554__A_N _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4397__A1 _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4820__S _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4121__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4857__C1 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4267__S _4271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4872__A2 _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5821__A1 _3926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5910_ _6029_/CLK _5910_/D vssd1 vssd1 vccd1 vccd1 _5910_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5841_ _3664_/X _5834_/X _5837_/X _5840_/X vssd1 vssd1 vccd1 vccd1 _5841_/X sky130_fd_sc_hd__o22a_1
X_5772_ hold554/X _5771_/X _5772_/S vssd1 vssd1 vccd1 vccd1 _5772_/X sky130_fd_sc_hd__mux2_1
X_2984_ _6154_/Q vssd1 vssd1 vccd1 vccd1 _2984_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_90_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4723_ _5767_/A hold458/X _4721_/X _4722_/X vssd1 vssd1 vccd1 vccd1 _4723_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_8_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4654_ hold82/A _5931_/Q _5923_/Q _6031_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4654_/X sky130_fd_sc_hd__mux4_1
X_4585_ _4219_/A _6161_/Q _4589_/S vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_71_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3605_ _3988_/A _3983_/S _3982_/S vssd1 vssd1 vccd1 vccd1 _3605_/X sky130_fd_sc_hd__and3_4
XANTENNA__4560__A1 _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout103_A _3377_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3536_ _4460_/A _4497_/S _4726_/D vssd1 vssd1 vccd1 vccd1 _3536_/X sky130_fd_sc_hd__and3_1
X_6255_ _6259_/CLK _6255_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6255_/Q sky130_fd_sc_hd__dfrtp_1
X_5206_ _6179_/Q _5104_/Y _5122_/Y _6195_/Q vssd1 vssd1 vccd1 vccd1 _5206_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5561__S _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3467_ _4765_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3711_/B sky130_fd_sc_hd__nor2_2
X_6186_ _6242_/CLK _6186_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6186_/Q sky130_fd_sc_hd__dfrtp_1
X_3398_ _3439_/B _3457_/A vssd1 vssd1 vccd1 vccd1 _3399_/B sky130_fd_sc_hd__nor2_1
X_5137_ _6173_/Q _5104_/Y _5109_/Y _5136_/X vssd1 vssd1 vccd1 vccd1 _5137_/X sky130_fd_sc_hd__a22o_1
X_5068_ hold36/X _4157_/Y _5073_/S vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__mux2_1
X_4019_ hold408/X _4021_/B _3646_/X _4018_/X vssd1 vssd1 vccd1 vccd1 _4019_/X sky130_fd_sc_hd__a31o_1
XANTENNA__3418__A3 _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3823__A0 _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4640__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4067__B1 _4750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4082__A3 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4116__A _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5031__A2 _6046_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4550__S _4596_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3593__A2 _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold108 _6007_/Q vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ hold183/X _4226_/X _4372_/S vssd1 vssd1 vccd1 vccd1 _4370_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4542__A1 _4836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold119 _4035_/X vssd1 vssd1 vccd1 vccd1 _5899_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3321_ _5424_/B _3321_/B vssd1 vssd1 vccd1 vccd1 _3321_/X sky130_fd_sc_hd__or2_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6040_ _6175_/CLK _6040_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6040_/Q sky130_fd_sc_hd__dfrtp_1
X_3252_ _6050_/Q _3252_/B vssd1 vssd1 vccd1 vccd1 _5498_/B sky130_fd_sc_hd__or2_4
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3183_ _4486_/A _4051_/B _3182_/B _3182_/A vssd1 vssd1 vccd1 vccd1 _3185_/C sky130_fd_sc_hd__o22a_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_16_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6031_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_5824_ _6242_/Q _5791_/X _5823_/X _5764_/B vssd1 vssd1 vccd1 vccd1 _5824_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_76_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5022__A2 _3496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5755_ _4119_/A _4963_/B _4677_/X _5762_/C vssd1 vssd1 vccd1 vccd1 _5755_/X sky130_fd_sc_hd__o22a_1
X_2967_ _2967_/A vssd1 vssd1 vccd1 vccd1 _4461_/A sky130_fd_sc_hd__inv_2
X_5686_ _6202_/Q _5698_/B vssd1 vssd1 vccd1 vccd1 _5687_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4706_ hold423/X _4612_/B _5762_/B _4474_/X vssd1 vssd1 vccd1 vccd1 _4706_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4781__B2 _4779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4637_ hold454/X _4636_/Y _5073_/S vssd1 vssd1 vccd1 vccd1 _4637_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold620 _4373_/X vssd1 vssd1 vccd1 vccd1 _6038_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 _6156_/Q vssd1 vssd1 vccd1 vccd1 hold631/X sky130_fd_sc_hd__dlygate4sd3_1
X_4568_ _6159_/Q _4567_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4568_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold642 _6164_/Q vssd1 vssd1 vccd1 vccd1 _3382_/A sky130_fd_sc_hd__buf_1
Xhold653 _6164_/Q vssd1 vssd1 vccd1 vccd1 hold653/X sky130_fd_sc_hd__dlygate4sd3_1
X_4499_ _4575_/A _4498_/B _4498_/C vssd1 vssd1 vccd1 vccd1 _4500_/B sky130_fd_sc_hd__a21o_1
X_3519_ _3511_/X _3519_/B _3519_/C vssd1 vssd1 vccd1 vccd1 _3519_/X sky130_fd_sc_hd__and3b_1
XANTENNA__5089__A2 _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6238_ _6238_/CLK _6238_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6238_/Q sky130_fd_sc_hd__dfstp_2
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ _6170_/CLK _6169_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6169_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4049__B1 _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4695__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5466__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4370__S _4372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5788__A0 _6178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3870_ _5896_/Q _6008_/Q _3885_/S vssd1 vssd1 vccd1 vccd1 _3870_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5540_ _5540_/A _5540_/B _5538_/Y vssd1 vssd1 vccd1 vccd1 _5540_/X sky130_fd_sc_hd__or3b_1
XANTENNA__6203__RESET_B fanout184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5471_ _5484_/S _5467_/X _5470_/Y _5330_/B vssd1 vssd1 vccd1 vccd1 _5471_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_53_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4422_ _4410_/B _4415_/X _4419_/X _4421_/X _5317_/A vssd1 vssd1 vccd1 vccd1 _4422_/X
+ sky130_fd_sc_hd__o41a_1
XANTENNA__5712__B1 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4353_ _4242_/X hold246/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4353_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4284_ _4150_/X hold270/X _4291_/S vssd1 vssd1 vccd1 vccd1 _5945_/D sky130_fd_sc_hd__mux2_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3304_ _5424_/A _3563_/A _3221_/X vssd1 vssd1 vccd1 vccd1 _3304_/X sky130_fd_sc_hd__a21o_1
X_6023_ _6035_/CLK _6023_/D vssd1 vssd1 vccd1 vccd1 _6023_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _3268_/B _4770_/B vssd1 vssd1 vccd1 vccd1 _4771_/B sky130_fd_sc_hd__or2_2
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4963__B _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3166_ _4486_/A _3249_/A vssd1 vssd1 vccd1 vccd1 _3167_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5779__A0 _6241_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3097_ _3303_/A _3563_/A vssd1 vssd1 vccd1 vccd1 _3097_/Y sky130_fd_sc_hd__nand2_2
XANTENNA_fanout170_A fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5243__A2 _5242_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xci2406_z80_192 vssd1 vssd1 vccd1 vccd1 ci2406_z80_192/HI io_oeb[7] sky130_fd_sc_hd__conb_1
X_5807_ hold593/X _5806_/X _5832_/S vssd1 vssd1 vccd1 vccd1 _6238_/D sky130_fd_sc_hd__mux2_1
X_3999_ _5046_/A _6120_/Q vssd1 vssd1 vccd1 vccd1 _3999_/X sky130_fd_sc_hd__or2_1
Xfanout69 _3885_/S vssd1 vssd1 vccd1 vccd1 _3982_/S sky130_fd_sc_hd__buf_4
XFILLER_0_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout58 _3270_/X vssd1 vssd1 vccd1 vccd1 _4999_/A1 sky130_fd_sc_hd__clkbuf_8
X_5738_ _4030_/Y _5715_/B _5715_/Y _5737_/X vssd1 vssd1 vccd1 vccd1 _5738_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4754__A1 _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5669_ _5668_/X _5658_/A _5705_/S vssd1 vssd1 vccd1 vccd1 _5670_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold472 _6226_/Q vssd1 vssd1 vccd1 vccd1 hold472/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold450 _6203_/Q vssd1 vssd1 vccd1 vccd1 _5698_/A sky130_fd_sc_hd__buf_1
Xhold461 _5612_/X vssd1 vssd1 vccd1 vccd1 _6195_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4601__S1 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold483 _5288_/X vssd1 vssd1 vccd1 vccd1 _6141_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 _6046_/Q vssd1 vssd1 vccd1 vccd1 hold494/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout83_A _3739_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold647_A _5936_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4365__S _4372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4668__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3796__A2 _3588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4745__A1 _5164_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5813__A2_N _5352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5458__C1 _5341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5828__A2_N _5352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3020_ _3210_/A _3203_/B _4485_/A vssd1 vssd1 vccd1 vccd1 _4051_/B sky130_fd_sc_hd__or3_4
X_4971_ _6184_/Q _4970_/X _5701_/S vssd1 vssd1 vccd1 vccd1 _4971_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3236__A1 _6172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3922_ _3921_/A _3646_/X _3921_/Y _3645_/X vssd1 vssd1 vccd1 vccd1 _3922_/X sky130_fd_sc_hd__a211o_1
X_3853_ _3811_/A _3811_/B _3809_/A vssd1 vssd1 vccd1 vccd1 _5448_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3619__S _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3784_ _3783_/X _3761_/B _3958_/S vssd1 vssd1 vccd1 vccd1 _3785_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5523_ _5524_/A _5524_/B vssd1 vssd1 vccd1 vccd1 _5540_/A sky130_fd_sc_hd__nor2_1
X_5454_ _6177_/Q _5352_/A _5354_/Y vssd1 vssd1 vccd1 vccd1 _5454_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4405_ _5790_/D _4404_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _6042_/D sky130_fd_sc_hd__mux2_1
X_5385_ _5385_/A _5385_/B vssd1 vssd1 vccd1 vccd1 _5389_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4336_ _4034_/X hold263/X _4336_/S vssd1 vssd1 vccd1 vccd1 _6003_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_10_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4267_ hold159/X _4193_/X _4271_/S vssd1 vssd1 vccd1 vccd1 _4267_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_31_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6243_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4198_ _6024_/Q _3599_/X _3601_/X _5969_/Q vssd1 vssd1 vccd1 vccd1 _4198_/X sky130_fd_sc_hd__a22o_1
X_6006_ _6006_/CLK _6006_/D vssd1 vssd1 vccd1 vccd1 _6006_/Q sky130_fd_sc_hd__dfxtp_1
X_3218_ _3234_/A _3218_/B _3234_/B _3218_/D vssd1 vssd1 vccd1 vccd1 _4770_/A sky130_fd_sc_hd__nand4_4
X_3149_ _3507_/C _3210_/C vssd1 vssd1 vccd1 vccd1 _4618_/A sky130_fd_sc_hd__nor2_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6125__RESET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5152__A1 _6157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3772__B _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4586__S0 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold280 _6168_/Q vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3163__B1 _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold291 _4458_/X vssd1 vssd1 vccd1 vccd1 _6051_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5455__A2 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5207__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4124__A _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5654__S _5705_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5391__A1 _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3941__A2 _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5170_ _6016_/Q _5200_/A2 _4255_/S _5949_/Q _4256_/S vssd1 vssd1 vccd1 vccd1 _5172_/A
+ sky130_fd_sc_hd__o221a_1
X_4121_ _4474_/A _4121_/B vssd1 vssd1 vccd1 vccd1 _4121_/X sky130_fd_sc_hd__or2_1
X_4052_ _5360_/D vssd1 vssd1 vccd1 vccd1 _4061_/D sky130_fd_sc_hd__inv_2
Xinput4 io_in[27] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_2
X_3003_ _5356_/A _3643_/A vssd1 vssd1 vccd1 vccd1 _3052_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4957__A1 _6157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4954_ _6183_/Q _4953_/X _5701_/S vssd1 vssd1 vccd1 vccd1 _4954_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3905_ _6139_/Q _3910_/C vssd1 vssd1 vccd1 vccd1 _3906_/B sky130_fd_sc_hd__and2_1
XANTENNA__4709__A1 _6160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4885_ _4885_/A _4885_/B vssd1 vssd1 vccd1 vccd1 _4901_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3836_ _4034_/S _3835_/X _3834_/X vssd1 vssd1 vccd1 vccd1 _3836_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_15_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5382__A1 _6046_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3767_ _3767_/A _3767_/B vssd1 vssd1 vccd1 vccd1 _3767_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5506_ _5503_/X _5504_/X _5505_/X _5501_/X vssd1 vssd1 vccd1 vccd1 _5506_/X sky130_fd_sc_hd__o31a_1
X_3698_ _6136_/Q _6137_/Q _6138_/Q vssd1 vssd1 vccd1 vccd1 _3910_/C sky130_fd_sc_hd__o21a_1
XANTENNA__3592__B _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5437_ _2978_/A _3192_/B _3646_/X _3824_/X _3825_/X vssd1 vssd1 vccd1 vccd1 _5437_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_2_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5368_ _6230_/Q _6174_/Q _5773_/B vssd1 vssd1 vccd1 vccd1 _5368_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4319_ _5297_/A _4319_/B vssd1 vssd1 vccd1 vccd1 _4327_/S sky130_fd_sc_hd__or2_4
XFILLER_0_10_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5299_ hold132/X _3737_/X _5305_/S vssd1 vssd1 vccd1 vccd1 _6146_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5437__A2 _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2952__A _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold512_A _6189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4879__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5125__A1 _6172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5125__B2 _6236_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4119__A _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4939__A1 _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4553__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4670_ _4669_/X _4668_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4963_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5364__B2 _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4789__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3621_ _3988_/A _3619_/X _3610_/X vssd1 vssd1 vccd1 vccd1 _5249_/A sky130_fd_sc_hd__o21ai_4
X_3552_ _3457_/A _3551_/X _3549_/X vssd1 vssd1 vccd1 vccd1 _3552_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_24_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3483_ _3483_/A _4727_/B _5338_/A _3483_/D vssd1 vssd1 vccd1 vccd1 _3483_/X sky130_fd_sc_hd__or4_1
X_5222_ _5225_/B _5228_/B _5222_/C vssd1 vssd1 vccd1 vccd1 _5222_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__3678__A1 _5116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5153_ _6207_/Q _5106_/Y _5129_/Y _6215_/Q vssd1 vssd1 vccd1 vccd1 _5163_/B sky130_fd_sc_hd__a22o_1
X_4104_ _6038_/Q _4104_/B _5120_/A _5107_/A vssd1 vssd1 vccd1 vccd1 _4105_/S sky130_fd_sc_hd__or4b_1
X_5084_ _5085_/B vssd1 vssd1 vccd1 vccd1 _5107_/B sky130_fd_sc_hd__inv_2
X_4035_ hold118/X _4034_/X _4035_/S vssd1 vssd1 vccd1 vccd1 _4035_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5986_ _6010_/CLK _5986_/D vssd1 vssd1 vccd1 vccd1 _5986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4937_ _6182_/Q _4936_/X _5701_/S vssd1 vssd1 vccd1 vccd1 _4937_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4868_ _4865_/B _4867_/X _5011_/S vssd1 vssd1 vccd1 vccd1 _4868_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_31 _5218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_20 _3517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5355__B2 _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3819_ _3699_/Y _3818_/X _6173_/Q vssd1 vssd1 vccd1 vccd1 _3820_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_62_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4799_ _6189_/Q _4815_/B _4798_/X vssd1 vssd1 vccd1 vccd1 _4799_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3380__A_N _4486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5202__S1 _5116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3108__A _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3841__A1 _6117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4397__A2 _6127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5346__A1 _5705_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3018__A _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4857__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5840_ _6113_/Q _5839_/X _5869_/S vssd1 vssd1 vccd1 vccd1 _5840_/X sky130_fd_sc_hd__mux2_1
X_5771_ _4030_/Y _5770_/X _5771_/S vssd1 vssd1 vccd1 vccd1 _5771_/X sky130_fd_sc_hd__mux2_1
X_2983_ _6155_/Q vssd1 vssd1 vccd1 vccd1 _4493_/B sky130_fd_sc_hd__inv_2
XFILLER_0_68_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4722_ _6161_/Q _4620_/Y _5073_/S vssd1 vssd1 vccd1 vccd1 _4722_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4653_ hold520/X _4652_/Y _5073_/S vssd1 vssd1 vccd1 vccd1 _4653_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4584_ hold552/X _4583_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _4584_/X sky130_fd_sc_hd__mux2_1
X_3604_ _3968_/A _3616_/B _3982_/S vssd1 vssd1 vccd1 vccd1 _4346_/A sky130_fd_sc_hd__or3_1
X_3535_ _6043_/Q _5834_/C _5740_/A _5834_/B vssd1 vssd1 vccd1 vccd1 _3535_/X sky130_fd_sc_hd__or4b_2
XFILLER_0_12_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3466_ _3525_/C _3466_/B vssd1 vssd1 vccd1 vccd1 _3466_/Y sky130_fd_sc_hd__nor2_1
X_6254_ _6259_/CLK _6254_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6254_/Q sky130_fd_sc_hd__dfrtp_1
X_5205_ _5767_/A _2980_/A _5086_/Y _5204_/X vssd1 vssd1 vccd1 vccd1 _5205_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_58_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6185_ _6242_/CLK _6185_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6185_/Q sky130_fd_sc_hd__dfrtp_1
X_3397_ _3394_/Y _3396_/X _4485_/B vssd1 vssd1 vccd1 vccd1 _3397_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5136_ _3678_/X _5105_/B _5135_/X vssd1 vssd1 vccd1 vccd1 _5136_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3520__B1 _3503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5067_ hold21/X _4143_/Y _5073_/S vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__mux2_1
X_4018_ _5046_/A _3648_/A _3650_/X _5384_/B vssd1 vssd1 vccd1 vccd1 _4018_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5289__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5969_ _6033_/CLK _5969_/D vssd1 vssd1 vccd1 vccd1 _5969_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3110__B _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4368__S _4372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5500__A1 _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4067__A1 _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3301__A _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5567__A1 _6158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4116__B _4116_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold109 _4341_/X vssd1 vssd1 vccd1 vccd1 _6007_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3750__B1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3320_ _5918_/Q _3320_/B vssd1 vssd1 vccd1 vccd1 _3320_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3446_/A _3276_/A _4483_/A _4439_/B _3250_/X vssd1 vssd1 vccd1 vccd1 _3251_/X
+ sky130_fd_sc_hd__a2111o_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ _3182_/A _3182_/B vssd1 vssd1 vccd1 vccd1 _3411_/D sky130_fd_sc_hd__nor2_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5823_ _6242_/Q _5352_/A _5457_/A hold472/X vssd1 vssd1 vccd1 vccd1 _5823_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5754_ hold571/X _5741_/Y _5753_/X _5767_/A vssd1 vssd1 vccd1 vccd1 _5754_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2966_ _2966_/A vssd1 vssd1 vccd1 vccd1 _2966_/Y sky130_fd_sc_hd__inv_2
X_5685_ _5685_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5687_/A sky130_fd_sc_hd__and2_1
X_4705_ _4705_/A _4705_/B vssd1 vssd1 vccd1 vccd1 _5762_/B sky130_fd_sc_hd__xor2_1
X_4636_ _4493_/B _4619_/X _4635_/Y vssd1 vssd1 vccd1 vccd1 _4636_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4042__A _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4977__A _6241_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3336__A3 _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold610 _4744_/X vssd1 vssd1 vccd1 vccd1 _6071_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 _6259_/Q vssd1 vssd1 vccd1 vccd1 hold621/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold632 _6155_/Q vssd1 vssd1 vccd1 vccd1 hold632/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 _6142_/Q vssd1 vssd1 vccd1 vccd1 hold654/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5730__B2 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4567_ _4565_/X _4566_/X _5872_/A vssd1 vssd1 vccd1 vccd1 _4567_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold643 _6126_/Q vssd1 vssd1 vccd1 vccd1 hold643/X sky130_fd_sc_hd__dlygate4sd3_1
X_4498_ _4575_/A _4498_/B _4498_/C vssd1 vssd1 vccd1 vccd1 _4498_/X sky130_fd_sc_hd__and3_1
X_3518_ _3513_/A _3508_/C hold611/X vssd1 vssd1 vccd1 vccd1 _3518_/Y sky130_fd_sc_hd__o21bai_1
X_6237_ _6242_/CLK _6237_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6237_/Q sky130_fd_sc_hd__dfstp_2
XANTENNA__5494__A0 _6240_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3449_ _4735_/A _3446_/A _3448_/Y _4398_/B vssd1 vssd1 vccd1 vccd1 _3449_/X sky130_fd_sc_hd__o211a_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ _6171_/CLK hold39/X fanout173/X vssd1 vssd1 vccd1 vccd1 _6168_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _5122_/A _5129_/B vssd1 vssd1 vccd1 vccd1 _5119_/Y sky130_fd_sc_hd__nor2_2
X_6099_ _6208_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5549__A1 _6157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3121__A _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2960__A _6178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5721__B2 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5485__B1 _5363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4826__S _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5511__A _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3799__B1 _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5470_ _5468_/X _5469_/X _5484_/S vssd1 vssd1 vccd1 vccd1 _5470_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4421_ _4053_/X _4054_/X _4749_/B _4618_/B vssd1 vssd1 vccd1 vccd1 _4421_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5712__A1 _4116_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4352_ _4226_/X hold230/X _4354_/S vssd1 vssd1 vccd1 vccd1 _4352_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5476__A0 _3959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4283_ _4292_/B _4364_/B vssd1 vssd1 vccd1 vccd1 _4291_/S sky130_fd_sc_hd__or2_4
X_3303_ _3303_/A _3303_/B vssd1 vssd1 vccd1 vccd1 _3303_/X sky130_fd_sc_hd__or2_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6022_ _6030_/CLK _6022_/D vssd1 vssd1 vccd1 vccd1 _6022_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3206__A _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _3234_/A _3234_/B _3234_/C _3234_/D vssd1 vssd1 vccd1 vccd1 _4770_/B sky130_fd_sc_hd__and4_2
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5421__A _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3165_ _4118_/B _4486_/B vssd1 vssd1 vccd1 vccd1 _3168_/C sky130_fd_sc_hd__or2_1
X_3096_ _3203_/A _4094_/D _3125_/C vssd1 vssd1 vccd1 vccd1 _3713_/A sky130_fd_sc_hd__or3_4
XFILLER_0_89_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout163_A hold588/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_193 vssd1 vssd1 vccd1 vccd1 ci2406_z80_193/HI io_oeb[8] sky130_fd_sc_hd__conb_1
X_5806_ _5805_/X _3785_/Y _5831_/S vssd1 vssd1 vccd1 vccd1 _5806_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3998_ _3998_/A _5370_/B vssd1 vssd1 vccd1 vccd1 _3998_/Y sky130_fd_sc_hd__nand2_1
Xfanout59 _5707_/S vssd1 vssd1 vccd1 vccd1 _5672_/S sky130_fd_sc_hd__buf_6
X_5737_ _4116_/Y _4879_/B _4594_/Y _5762_/C vssd1 vssd1 vccd1 vccd1 _5737_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2949_ _4094_/D vssd1 vssd1 vccd1 vccd1 _3148_/C sky130_fd_sc_hd__inv_2
XFILLER_0_32_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5668_ _5667_/X _6158_/Q _5704_/S vssd1 vssd1 vccd1 vccd1 _5668_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5703__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5599_ _5598_/X _5593_/X _5670_/A vssd1 vssd1 vccd1 vccd1 _5599_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4619_ _4617_/X _4618_/X _4497_/S vssd1 vssd1 vccd1 vccd1 _4619_/X sky130_fd_sc_hd__o21a_4
Xhold451 _5707_/X vssd1 vssd1 vccd1 vccd1 _6203_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold462 _6041_/Q vssd1 vssd1 vccd1 vccd1 _5790_/C sky130_fd_sc_hd__clkbuf_2
Xhold440 _5321_/X vssd1 vssd1 vccd1 vccd1 _6164_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 _5780_/X vssd1 vssd1 vccd1 vccd1 _6226_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 _6114_/Q vssd1 vssd1 vccd1 vccd1 hold484/X sky130_fd_sc_hd__buf_1
XANTENNA__3190__A1 _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold495 _4453_/X vssd1 vssd1 vccd1 vccd1 _6046_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout76_A _5698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2955__A _3302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5050__B _5050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4442__A1 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5155__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_1_wb_clk_i _5978_/CLK vssd1 vssd1 vccd1 vccd1 _6010_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__4410__A _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5170__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_43_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4681__A1 _4538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4970_ _6200_/Q _4815_/B _4961_/X _4969_/X vssd1 vssd1 vccd1 vccd1 _4970_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4984__A2 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3921_ _3921_/A _3950_/B vssd1 vssd1 vccd1 vccd1 _3921_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4291__S _4291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3852_ _3899_/A _3852_/B vssd1 vssd1 vccd1 vccd1 _3855_/A sky130_fd_sc_hd__and2_1
XFILLER_0_73_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3783_ _4507_/B _3782_/X _6074_/Q vssd1 vssd1 vccd1 vccd1 _3783_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5522_ _6155_/Q _5507_/Y _5508_/X vssd1 vssd1 vccd1 vccd1 _5524_/B sky130_fd_sc_hd__o21ai_1
X_5453_ hold616/X _5452_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _5453_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5416__A _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5384_ _5384_/A _5384_/B vssd1 vssd1 vccd1 vccd1 _5385_/B sky130_fd_sc_hd__xor2_1
X_4404_ _5250_/B _4410_/B _5317_/A vssd1 vssd1 vccd1 vccd1 _4404_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4335_ _3979_/X hold114/X _4336_/S vssd1 vssd1 vccd1 vccd1 _4335_/X sky130_fd_sc_hd__mux2_1
X_4266_ hold54/X _4180_/X _4271_/S vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__mux2_1
X_4197_ _4145_/B _4174_/X _4195_/X _4196_/X vssd1 vssd1 vccd1 vccd1 _4207_/A sky130_fd_sc_hd__a31oi_2
X_3217_ _3211_/Y _3212_/X _3215_/Y _3216_/X _3457_/A vssd1 vssd1 vccd1 vccd1 _3218_/D
+ sky130_fd_sc_hd__a41o_1
X_6005_ _6146_/CLK _6005_/D vssd1 vssd1 vccd1 vccd1 _6005_/Q sky130_fd_sc_hd__dfxtp_1
X_3148_ _3210_/A _3148_/B _3148_/C _3210_/C vssd1 vssd1 vccd1 vccd1 _3554_/A sky130_fd_sc_hd__or4_4
XANTENNA__4990__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3079_ _3148_/C _4398_/A _3507_/C _3210_/A vssd1 vssd1 vccd1 vccd1 _3079_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_37_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold270 _5945_/Q vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4586__S1 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3163__A1 _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5763__B1_N _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold281 _5318_/X vssd1 vssd1 vccd1 vccd1 _6162_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 _5996_/Q vssd1 vssd1 vccd1 vccd1 _2966_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4663__B2 _4474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5860__A0 _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3941__A3 _6119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5143__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4120_ _4963_/A _4121_/B _4474_/A vssd1 vssd1 vccd1 vccd1 _4120_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__4286__S _4291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4051_ _4725_/B _4051_/B _4056_/A vssd1 vssd1 vccd1 vccd1 _5360_/D sky130_fd_sc_hd__or3_2
Xinput5 io_in[28] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_2
X_3002_ _3539_/A _3389_/B hold92/X _4077_/A vssd1 vssd1 vccd1 vccd1 _3268_/B sky130_fd_sc_hd__o31a_1
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4953_ _6199_/Q _4815_/B _4945_/X _4952_/X vssd1 vssd1 vccd1 vccd1 _4953_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_86_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3904_ _3894_/A _6140_/Q _6118_/Q _3848_/B _3903_/X vssd1 vssd1 vccd1 vccd1 _5373_/B
+ sky130_fd_sc_hd__o41a_2
X_4884_ _6054_/Q _6055_/Q _6058_/Q _6059_/Q vssd1 vssd1 vccd1 vccd1 _4885_/B sky130_fd_sc_hd__and4_1
XANTENNA__4709__A2 _4620_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3835_ hold197/X hold163/X hold237/X hold112/X _5179_/S _3740_/S vssd1 vssd1 vccd1
+ vccd1 _3835_/X sky130_fd_sc_hd__mux4_2
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3766_ _3687_/A _3687_/B _3684_/A vssd1 vssd1 vccd1 vccd1 _3767_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5505_ _6127_/Q _3396_/D _3711_/B _4044_/B _3334_/B vssd1 vssd1 vccd1 vccd1 _5505_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5436_ hold573/X _5375_/B _5460_/S vssd1 vssd1 vccd1 vccd1 _5436_/X sky130_fd_sc_hd__mux2_1
X_3697_ _3645_/X _3695_/B _3696_/X _6114_/Q _3693_/X vssd1 vssd1 vccd1 vccd1 _3704_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5367_ hold651/X _5366_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _6173_/D sky130_fd_sc_hd__mux2_1
X_5298_ hold84/X _3668_/X _5305_/S vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__mux2_1
X_4318_ _4034_/X hold106/X _4318_/S vssd1 vssd1 vccd1 vccd1 _4318_/X sky130_fd_sc_hd__mux2_1
X_4249_ _4249_/A _4249_/B vssd1 vssd1 vccd1 vccd1 _4250_/B sky130_fd_sc_hd__or2_1
XFILLER_0_97_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__6206__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold338_A _6129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4879__B _4879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3384__A1 _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5490__S _5497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4895__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4119__B _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4834__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4495__S0 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3620_ _3988_/A _3619_/X _3610_/X vssd1 vssd1 vccd1 vccd1 _3620_/X sky130_fd_sc_hd__o21a_1
X_3551_ _5424_/A _4446_/B _5424_/C _3563_/A _3550_/X vssd1 vssd1 vccd1 vccd1 _3551_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3482_ _4739_/A _4614_/B _4729_/A _4094_/B _4439_/B vssd1 vssd1 vccd1 vccd1 _3483_/D
+ sky130_fd_sc_hd__a2111o_1
X_5221_ _5225_/B _5228_/B _5222_/C vssd1 vssd1 vccd1 vccd1 _5221_/X sky130_fd_sc_hd__or3_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5152_ _6157_/Q _5121_/Y _5122_/Y _6191_/Q vssd1 vssd1 vccd1 vccd1 _5163_/A sky130_fd_sc_hd__a22o_1
X_4103_ _4094_/D _4077_/X _4102_/X _5220_/A vssd1 vssd1 vccd1 vccd1 _5107_/A sky130_fd_sc_hd__a22o_4
XANTENNA__4627__A1 _4915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5083_ _4618_/B _5080_/Y _5081_/X _5082_/X _5220_/A vssd1 vssd1 vccd1 vccd1 _5085_/B
+ sky130_fd_sc_hd__o221a_4
X_4034_ _4032_/X _4033_/X _4034_/S vssd1 vssd1 vccd1 vccd1 _4034_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_78_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5985_ _6006_/CLK _5985_/D vssd1 vssd1 vccd1 vccd1 _5985_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ _6198_/Q _4815_/B _4930_/X _4935_/X vssd1 vssd1 vccd1 vccd1 _4936_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_86_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4867_ _6194_/Q _6060_/Q _5216_/A vssd1 vssd1 vccd1 vccd1 _4867_/X sky130_fd_sc_hd__mux2_1
XANTENNA_21 _3434_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_32 _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_10 _4418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3818_ _6136_/Q _6137_/Q _6138_/Q vssd1 vssd1 vccd1 vccd1 _3818_/X sky130_fd_sc_hd__or3_1
XFILLER_0_62_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4798_ _6205_/Q _4768_/Y _4791_/X _4797_/X vssd1 vssd1 vccd1 vccd1 _4798_/X sky130_fd_sc_hd__a211o_1
X_3749_ _5894_/Q _6006_/Q _3982_/S vssd1 vssd1 vccd1 vccd1 _3749_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_100_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5419_ _6159_/Q _6158_/Q vssd1 vssd1 vccd1 vccd1 _5420_/B sky130_fd_sc_hd__nand2_1
XANTENNA__3823__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap56 _4768_/Y vssd1 vssd1 vccd1 vccd1 _5009_/A2 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5043__B2 _6115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5043__A1 _6117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5594__A2 _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3357__A1 _3370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4857__B2 _4850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4468__S0 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5770_ hold554/X _5713_/Y _5769_/X _5762_/A vssd1 vssd1 vccd1 vccd1 _5770_/X sky130_fd_sc_hd__o22a_1
X_2982_ _6046_/Q vssd1 vssd1 vccd1 vccd1 _5479_/S sky130_fd_sc_hd__inv_2
XFILLER_0_8_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4721_ _5764_/B _4719_/X _4720_/X vssd1 vssd1 vccd1 vccd1 _4721_/X sky130_fd_sc_hd__a21o_1
X_4652_ _4507_/B _4619_/X _4651_/Y vssd1 vssd1 vccd1 vccd1 _4652_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3603_ _3988_/A _3983_/S _3724_/S vssd1 vssd1 vccd1 vccd1 _3603_/X sky130_fd_sc_hd__and3_4
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4583_ _6160_/Q _4582_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4583_/X sky130_fd_sc_hd__mux2_1
X_3534_ _5740_/A _5834_/C vssd1 vssd1 vccd1 vccd1 _5790_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3465_ _4750_/A _5507_/B _4485_/B vssd1 vssd1 vccd1 vccd1 _3466_/B sky130_fd_sc_hd__o21a_1
X_6253_ _6259_/CLK _6253_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6253_/Q sky130_fd_sc_hd__dfrtp_1
X_5204_ _5204_/A _5204_/B _5204_/C _5204_/D vssd1 vssd1 vccd1 vccd1 _5204_/X sky130_fd_sc_hd__or4_1
XANTENNA__5424__A _5424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6184_ _6242_/CLK _6184_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6184_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3520__A1 _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3396_ _3396_/A _5502_/D _3545_/A _3396_/D vssd1 vssd1 vccd1 vccd1 _3396_/X sky130_fd_sc_hd__or4_1
X_5135_ _5116_/A _4164_/X _5185_/S _5134_/X vssd1 vssd1 vccd1 vccd1 _5135_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5066_ hold3/X _3990_/B _5296_/S vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__mux2_1
XFILLER_0_79_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5273__A1 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4017_ _6120_/Q _4021_/B vssd1 vssd1 vccd1 vccd1 _5044_/A sky130_fd_sc_hd__and2_1
XFILLER_0_94_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5968_ _6035_/CLK _5968_/D vssd1 vssd1 vccd1 vccd1 _5968_/Q sky130_fd_sc_hd__dfxtp_1
X_4919_ _6155_/Q _5013_/S vssd1 vssd1 vccd1 vccd1 _4919_/X sky130_fd_sc_hd__or2_1
X_5899_ _6152_/CLK _5899_/D vssd1 vssd1 vccd1 vccd1 _5899_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5328__A2 _3496_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4536__A0 _6157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3339__A1 _5918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2958__A _6174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5500__A2 _5313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4067__A2 _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3750__A1 _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3250_ _5502_/A _3277_/A _4094_/B _3250_/D vssd1 vssd1 vccd1 vccd1 _3250_/X sky130_fd_sc_hd__or4_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _4737_/A _4486_/A _4417_/B vssd1 vssd1 vccd1 vccd1 _4385_/A sky130_fd_sc_hd__or3_2
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5255__A1 _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5255__B2 _6236_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4294__S _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5822_ _2990_/A _5821_/X _5832_/S vssd1 vssd1 vccd1 vccd1 _5822_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5753_ _3832_/Y _5771_/S _5742_/Y _5752_/X vssd1 vssd1 vccd1 vccd1 _5753_/X sky130_fd_sc_hd__o22a_1
X_4704_ _4703_/A _4703_/B _4703_/C _4705_/A vssd1 vssd1 vccd1 vccd1 _4716_/B sky130_fd_sc_hd__a31o_1
XANTENNA__5419__A _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4230__A2 _3588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2965_ _5957_/Q vssd1 vssd1 vccd1 vccd1 _2965_/Y sky130_fd_sc_hd__inv_2
X_5684_ _5679_/A _5625_/Y _5683_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _5684_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5853__S _5869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4635_ _5764_/B _4633_/X _4634_/X vssd1 vssd1 vccd1 vccd1 _4635_/Y sky130_fd_sc_hd__a21oi_1
Xhold600 _5812_/X vssd1 vssd1 vccd1 vccd1 _6239_/D sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_25_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6119_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_4566_ hold559/X input6/X _4596_/S vssd1 vssd1 vccd1 vccd1 _4566_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold611 _6170_/Q vssd1 vssd1 vccd1 vccd1 hold611/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4977__B _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold644 _5230_/X vssd1 vssd1 vccd1 vccd1 _6126_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3517_ _3517_/A _3517_/B _3517_/C _3508_/X vssd1 vssd1 vccd1 vccd1 _3519_/B sky130_fd_sc_hd__or4b_1
XANTENNA__4469__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold622 _5891_/X vssd1 vssd1 vccd1 vccd1 _6259_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 _6258_/Q vssd1 vssd1 vccd1 vccd1 hold633/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold655 _5293_/X vssd1 vssd1 vccd1 vccd1 _6142_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4497_ _6205_/Q _4789_/B _4497_/S vssd1 vssd1 vccd1 vccd1 _4498_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_40_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6236_ _6242_/CLK _6236_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6236_/Q sky130_fd_sc_hd__dfstp_2
X_3448_ _4737_/A _4398_/C vssd1 vssd1 vccd1 vccd1 _3448_/Y sky130_fd_sc_hd__nor2_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ _6167_/CLK _6167_/D fanout173/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dfrtp_1
X_3379_ _3434_/B _4486_/B _3208_/A _4460_/A vssd1 vssd1 vccd1 vccd1 _3392_/A sky130_fd_sc_hd__o211a_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _5120_/A _5185_/S vssd1 vssd1 vccd1 vccd1 _5129_/B sky130_fd_sc_hd__or2_1
XANTENNA__5798__A1_N _6237_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6098_ _6148_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
X_5049_ _5031_/X _5039_/X _5048_/X _5026_/A _2960_/Y vssd1 vssd1 vccd1 vccd1 _5050_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_94_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_2_3__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4932__S _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5511__B _5629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5237__B2 _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5237__A1 _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4748__B1 _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3971__A1 _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4420_ _4124_/B _3097_/Y _5838_/B _4618_/C _3469_/Y vssd1 vssd1 vccd1 vccd1 _4749_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5712__A2 _5711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4289__S _4291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4920__B1 _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4351_ _4211_/X hold266/X _4354_/S vssd1 vssd1 vccd1 vccd1 _6016_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4282_ hold110/X _4261_/X _4282_/S vssd1 vssd1 vccd1 vccd1 _4282_/X sky130_fd_sc_hd__mux2_1
X_3302_ _3302_/A _5838_/C vssd1 vssd1 vccd1 vccd1 _3303_/B sky130_fd_sc_hd__or2_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ _6034_/CLK _6021_/D vssd1 vssd1 vccd1 vccd1 _6021_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3206__B _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _3211_/Y _3212_/X _3231_/X _3337_/D _3457_/A vssd1 vssd1 vccd1 vccd1 _3234_/D
+ sky130_fd_sc_hd__a41o_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5421__B _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3164_ _3210_/C _3622_/C _3163_/X _4485_/B vssd1 vssd1 vccd1 vccd1 _3164_/Y sky130_fd_sc_hd__o31ai_1
X_3095_ _3249_/A _3125_/C vssd1 vssd1 vccd1 vccd1 _3563_/A sky130_fd_sc_hd__or2_2
XFILLER_0_76_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5848__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout156_A _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xci2406_z80_194 vssd1 vssd1 vccd1 vccd1 ci2406_z80_194/HI io_oeb[9] sky130_fd_sc_hd__conb_1
X_5805_ hold349/X _5794_/Y _5804_/X _5794_/B vssd1 vssd1 vccd1 vccd1 _5805_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_91_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3997_ _3998_/A _5370_/B vssd1 vssd1 vccd1 vccd1 _3997_/X sky130_fd_sc_hd__or2_1
XFILLER_0_91_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5736_ hold550/X _5714_/Y _5735_/X _5023_/A vssd1 vssd1 vccd1 vccd1 _5736_/X sky130_fd_sc_hd__o22a_1
X_2948_ _3203_/B vssd1 vssd1 vccd1 vccd1 _3148_/B sky130_fd_sc_hd__inv_2
X_5667_ _5694_/A _5666_/X _4959_/Y vssd1 vssd1 vccd1 vccd1 _5667_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4618_ _4618_/A _4618_/B _4618_/C vssd1 vssd1 vccd1 vccd1 _4618_/X sky130_fd_sc_hd__and3_1
X_5598_ _5597_/X _2996_/A _5705_/S vssd1 vssd1 vccd1 vccd1 _5598_/X sky130_fd_sc_hd__mux2_1
Xhold441 _6220_/Q vssd1 vssd1 vccd1 vccd1 hold441/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold430 _5784_/X vssd1 vssd1 vccd1 vccd1 _6230_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold452 _6207_/Q vssd1 vssd1 vccd1 vccd1 hold452/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _4403_/X vssd1 vssd1 vccd1 vccd1 _6041_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4549_ _4547_/Y _4548_/X _4565_/S vssd1 vssd1 vccd1 vccd1 _4549_/X sky130_fd_sc_hd__mux2_1
Xhold474 _6235_/Q vssd1 vssd1 vccd1 vccd1 hold474/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 _5140_/X vssd1 vssd1 vccd1 vccd1 _6114_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 _6077_/Q vssd1 vssd1 vccd1 vccd1 _5222_/C sky130_fd_sc_hd__clkbuf_2
XANTENNA__3190__A2 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4927__S _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5467__A1 _6178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6219_ _6219_/CLK _6219_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6219_/Q sky130_fd_sc_hd__dfstp_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3132__A _3694_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4978__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3953__A1 _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5493__S _5497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5155__B1 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4410__B _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4837__S _5216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3741__S _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4681__A2 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5630__A1 _6197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3920_ _3920_/A _5397_/B vssd1 vssd1 vccd1 vccd1 _3920_/X sky130_fd_sc_hd__and2_1
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3851_ _6139_/Q _3851_/B _3851_/C vssd1 vssd1 vccd1 vccd1 _3852_/B sky130_fd_sc_hd__or3_1
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3782_ _3624_/Y _5375_/A _3781_/X vssd1 vssd1 vccd1 vccd1 _3782_/X sky130_fd_sc_hd__a21bo_1
X_5521_ _5514_/A _5520_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _6188_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_14_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5452_ _5363_/X _5447_/X _5451_/X _5326_/X _3864_/Y vssd1 vssd1 vccd1 vccd1 _5452_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5416__B _6160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4403_ _5790_/C _4402_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _4403_/X sky130_fd_sc_hd__mux2_1
X_5383_ _6135_/Q _5383_/B vssd1 vssd1 vccd1 vccd1 _5385_/A sky130_fd_sc_hd__xnor2_1
X_4334_ _3930_/X hold102/X _4336_/S vssd1 vssd1 vccd1 vccd1 _4334_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4265_ hold78/X _4165_/X _4271_/S vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__mux2_1
X_6004_ _6010_/CLK _6004_/D vssd1 vssd1 vccd1 vccd1 _6004_/Q sky130_fd_sc_hd__dfxtp_1
X_4196_ _4143_/Y _4157_/Y _4173_/B _4187_/B _4219_/A vssd1 vssd1 vccd1 vccd1 _4196_/X
+ sky130_fd_sc_hd__o41a_1
X_3216_ _3540_/A _4446_/A _3543_/B _5362_/B _3439_/B vssd1 vssd1 vccd1 vccd1 _3216_/X
+ sky130_fd_sc_hd__o221a_1
X_3147_ _4391_/B _3074_/Y _4094_/B _3143_/Y _3052_/A vssd1 vssd1 vccd1 vccd1 _3158_/A
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_96_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4990__B _4990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5578__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4482__S _4598_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3078_ _4739_/A _3249_/B vssd1 vssd1 vccd1 vccd1 _3131_/B sky130_fd_sc_hd__or2_1
XFILLER_0_64_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6259_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5719_ _4119_/A _4789_/B _4501_/X _5762_/C vssd1 vssd1 vccd1 vccd1 _5719_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3699__B1 _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3163__A2 _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 _5994_/Q vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 _5898_/Q vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 _5951_/Q vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 _4329_/X vssd1 vssd1 vccd1 vccd1 _5996_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold652_A _6130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4663__A2 _4612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5860__A1 _6114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3871__B1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5488__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4887__C1 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5252__A _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4567__S _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4794__C _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4050_ _4037_/X _4048_/X _4049_/X _4415_/A _3112_/A vssd1 vssd1 vccd1 vccd1 _4050_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__4103__B2 _5220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 io_in[29] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_2
X_3001_ _3001_/A vssd1 vssd1 vccd1 vccd1 _6047_/D sky130_fd_sc_hd__inv_2
XANTENNA__3862__A0 _4538_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5851__B2 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _4999_/A1 _4947_/X _4951_/X _4824_/B vssd1 vssd1 vccd1 vccd1 _4952_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_52_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3903_ _3639_/X _3900_/A _3900_/Y _3901_/X _3902_/X vssd1 vssd1 vccd1 vccd1 _3903_/X
+ sky130_fd_sc_hd__a221o_1
X_4883_ _6056_/Q _6057_/Q _6060_/Q _6061_/Q vssd1 vssd1 vccd1 vccd1 _4885_/A sky130_fd_sc_hd__and4_1
X_3834_ hold19/X _4253_/A2 _3803_/Y _3833_/Y _3671_/B vssd1 vssd1 vccd1 vccd1 _3834_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_15_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3765_ _3765_/A _3765_/B vssd1 vssd1 vccd1 vccd1 _3767_/A sky130_fd_sc_hd__and2_1
X_3696_ _3646_/X _3695_/B _3695_/Y _3645_/X vssd1 vssd1 vccd1 vccd1 _3696_/X sky130_fd_sc_hd__a211o_1
X_5504_ _3484_/A _4427_/B _4439_/X _4038_/A vssd1 vssd1 vccd1 vccd1 _5504_/X sky130_fd_sc_hd__o31a_1
X_5435_ hold404/X _5872_/A _5365_/S _5434_/X vssd1 vssd1 vccd1 vccd1 _5435_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5861__S _5869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5366_ _3707_/X _5326_/X _5363_/X _5365_/X vssd1 vssd1 vccd1 vccd1 _5366_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5297_ _5297_/A _5297_/B vssd1 vssd1 vccd1 vccd1 _5305_/S sky130_fd_sc_hd__nor2_4
X_4317_ _3979_/X hold161/X _4318_/S vssd1 vssd1 vccd1 vccd1 _4317_/X sky130_fd_sc_hd__mux2_1
X_4248_ _5952_/Q _3605_/X _3615_/X _6035_/Q _4247_/X vssd1 vssd1 vccd1 vccd1 _4249_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5842__B2 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4179_ hold100/X hold54/X hold186/X hold66/X _5182_/S _4255_/S vssd1 vssd1 vccd1
+ vccd1 _4179_/X sky130_fd_sc_hd__mux4_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold400_A _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4581__A1 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3384__A2 _5313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5771__S _5771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4895__B _4895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4636__A2 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4192__S0 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3844__A0 _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5011__S _5011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3320__A _5918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4495__S1 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5349__A0 _3664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5247__A _5250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3550_ _3303_/A _3554_/A _4046_/B vssd1 vssd1 vccd1 vccd1 _3550_/X sky130_fd_sc_hd__a21o_1
XANTENNA__6056__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5220_ _5220_/A _5222_/C vssd1 vssd1 vccd1 vccd1 _5220_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3481_ _4615_/B _4614_/C vssd1 vssd1 vccd1 vccd1 _5338_/A sky130_fd_sc_hd__or2_1
X_5151_ _5023_/A _2977_/A _5086_/Y _5150_/X vssd1 vssd1 vccd1 vccd1 _5151_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4297__S _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5082_ _4124_/B _3097_/Y _4087_/X _4391_/B vssd1 vssd1 vccd1 vccd1 _5082_/X sky130_fd_sc_hd__a22o_1
X_4102_ _3539_/A _4099_/X _4101_/X _4618_/B vssd1 vssd1 vccd1 vccd1 _4102_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5824__A1 _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5824__B2 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3214__B _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4033_ hold168/X hold58/X hold106/X hold76/X _5179_/S _3740_/S vssd1 vssd1 vccd1
+ vccd1 _4033_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5984_ _6029_/CLK _5984_/D vssd1 vssd1 vccd1 vccd1 _5984_/Q sky130_fd_sc_hd__dfxtp_1
X_4935_ _4999_/A1 _4932_/X _4934_/X _4824_/B vssd1 vssd1 vccd1 vccd1 _4935_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_74_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5856__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_22 _3959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4866_ _6060_/Q _4764_/X _4763_/B vssd1 vssd1 vccd1 vccd1 _4866_/X sky130_fd_sc_hd__a21o_1
XANTENNA_11 _3477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3817_ _6136_/Q _6137_/Q _6138_/Q _3912_/B vssd1 vssd1 vccd1 vccd1 _3817_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_0_55_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4797_ _4999_/A1 _4793_/X _4796_/Y _4824_/B vssd1 vssd1 vccd1 vccd1 _4797_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_33 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3748_ _3983_/S _3748_/B vssd1 vssd1 vccd1 vccd1 _3748_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__4061__A _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3679_ _6114_/Q _5333_/B vssd1 vssd1 vccd1 vccd1 _3683_/B sky130_fd_sc_hd__and2b_1
X_5418_ _6159_/Q _6158_/Q vssd1 vssd1 vccd1 vccd1 _5474_/C sky130_fd_sc_hd__or2_1
X_5349_ _3664_/X _5348_/X _5487_/S vssd1 vssd1 vccd1 vccd1 _5349_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3405__A _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4670__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5200__C1 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5503__B1 _4043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5006__S _5020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5806__A1 _3785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4845__S _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output32_A _6089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4490__B1 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3293__B2 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4468__S1 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2981_ _6176_/Q vssd1 vssd1 vccd1 vccd1 _5445_/A sky130_fd_sc_hd__inv_2
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4720_ hold458/X _5762_/A _4619_/X vssd1 vssd1 vccd1 vccd1 _4720_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3596__A2 _3513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4651_ _5764_/B _4649_/X _4650_/X vssd1 vssd1 vccd1 vccd1 _4651_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3602_ _3968_/A _3983_/S _3724_/S vssd1 vssd1 vccd1 vccd1 _4319_/B sky130_fd_sc_hd__or3_1
XFILLER_0_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4582_ _4580_/X _4581_/X _5762_/A vssd1 vssd1 vccd1 vccd1 _4582_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_52_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3533_ _3531_/Y _5837_/A _3533_/S vssd1 vssd1 vccd1 vccd1 _5834_/C sky130_fd_sc_hd__mux2_2
XFILLER_0_52_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3209__B _5838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6252_ _6259_/CLK _6252_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6252_/Q sky130_fd_sc_hd__dfrtp_1
X_3464_ _3496_/C _5424_/C _3333_/B vssd1 vssd1 vccd1 vccd1 _5507_/B sky130_fd_sc_hd__o21ai_4
X_6183_ _6235_/CLK _6183_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6183_/Q sky130_fd_sc_hd__dfrtp_1
X_5203_ _6194_/Q _5122_/Y _5202_/X _5109_/Y vssd1 vssd1 vccd1 vccd1 _5204_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_58_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5424__B _5424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5134_ _5209_/A _5134_/B _5134_/C vssd1 vssd1 vccd1 vccd1 _5134_/X sky130_fd_sc_hd__or3_1
XFILLER_0_58_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3225__A _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3395_ _6048_/Q _3395_/B _6050_/Q vssd1 vssd1 vccd1 vccd1 _3396_/D sky130_fd_sc_hd__and3b_1
XANTENNA__3520__A2 _5314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5065_ hold1/X _3970_/B _5296_/S vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__mux2_1
XFILLER_0_74_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4016_ _4008_/Y _4015_/X _6173_/Q vssd1 vssd1 vccd1 vccd1 _5384_/B sky130_fd_sc_hd__mux2_1
XANTENNA__3284__A1 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_2__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2__f_wb_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5050__A_N _5052_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5967_ _6111_/CLK _5967_/D vssd1 vssd1 vccd1 vccd1 _5967_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5586__S _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4918_ _6063_/Q _4918_/B vssd1 vssd1 vccd1 vccd1 _4918_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5898_ _6010_/CLK _5898_/D vssd1 vssd1 vccd1 vccd1 _5898_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4849_ hold328/X _4848_/X _4927_/S vssd1 vssd1 vccd1 vccd1 _4849_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_99_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_23_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout99_A _4765_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3135__A _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5496__S _5497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ _4486_/A _3180_/B vssd1 vssd1 vccd1 vccd1 _3477_/C sky130_fd_sc_hd__nor2_2
XFILLER_0_28_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5821_ _5820_/X _3926_/X _5831_/S vssd1 vssd1 vccd1 vccd1 _5821_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5752_ _4119_/A _4943_/B _4662_/X _5762_/C vssd1 vssd1 vccd1 vccd1 _5752_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3919__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2964_ hold50/A vssd1 vssd1 vccd1 vccd1 _2964_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5419__B _6158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4703_ _4703_/A _4703_/B _4703_/C vssd1 vssd1 vccd1 vccd1 _4705_/B sky130_fd_sc_hd__and3_1
XFILLER_0_44_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5683_ _5670_/A _5681_/Y _5682_/X _5629_/Y _5676_/X vssd1 vssd1 vccd1 vccd1 _5683_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4634_ hold454/X _5762_/A _4619_/X vssd1 vssd1 vccd1 vccd1 _4634_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_44_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4518__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 _6179_/Q vssd1 vssd1 vccd1 vccd1 hold601/X sky130_fd_sc_hd__dlygate4sd3_1
X_4565_ _4563_/Y _4564_/X _4565_/S vssd1 vssd1 vccd1 vccd1 _4565_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold612 _3518_/Y vssd1 vssd1 vccd1 vccd1 _3519_/C sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3726__C1 _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold623 _6157_/Q vssd1 vssd1 vccd1 vccd1 hold623/X sky130_fd_sc_hd__dlygate4sd3_1
X_3516_ _3510_/X _3511_/X _3516_/C _3516_/D vssd1 vssd1 vccd1 vccd1 _3516_/X sky130_fd_sc_hd__and4bb_1
Xhold645 _6095_/Q vssd1 vssd1 vccd1 vccd1 _3502_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 _5889_/X vssd1 vssd1 vccd1 vccd1 _6258_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4496_ _4495_/X _4494_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4789_/B sky130_fd_sc_hd__mux2_2
Xhold656 _6131_/Q vssd1 vssd1 vccd1 vccd1 hold656/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6235_ _6235_/CLK _6235_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6235_/Q sky130_fd_sc_hd__dfstp_1
X_3447_ _3395_/B _5498_/B _3543_/A vssd1 vssd1 vccd1 vccd1 _3447_/X sky130_fd_sc_hd__a21o_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6166_ _6167_/CLK _6166_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6166_/Q sky130_fd_sc_hd__dfrtp_4
X_3378_ _4497_/S _3461_/A hold653/X _4725_/B vssd1 vssd1 vccd1 vccd1 _3378_/Y sky130_fd_sc_hd__o31ai_2
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5117_ _5209_/A _4133_/X _5105_/B _5116_/X vssd1 vssd1 vccd1 vccd1 _5117_/X sky130_fd_sc_hd__a211o_1
X_6097_ _6148_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
X_5048_ _5384_/A _5384_/B _5034_/X _5047_/X vssd1 vssd1 vccd1 vccd1 _5048_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_94_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3121__C _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3965__C1 _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5080__A _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4540__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4424__A _5502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4748__A1 _5164_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3739__S _3739_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4350_ _4193_/X hold289/X _4354_/S vssd1 vssd1 vccd1 vccd1 _6015_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3301_ _4124_/A _3301_/B vssd1 vssd1 vccd1 vccd1 _5838_/C sky130_fd_sc_hd__and2_2
X_4281_ hold64/X _4242_/X _4282_/S vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__mux2_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ _6110_/CLK _6020_/D vssd1 vssd1 vccd1 vccd1 _6020_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _3540_/A _5424_/A vssd1 vssd1 vccd1 vccd1 _3337_/D sky130_fd_sc_hd__or2_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _4070_/B _4036_/B _3446_/A vssd1 vssd1 vccd1 vccd1 _3163_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3503__A _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3094_ _3507_/C _3125_/C vssd1 vssd1 vccd1 vccd1 _3303_/A sky130_fd_sc_hd__or2_2
XANTENNA__4987__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5804_ _6238_/Q _5791_/X _5803_/X _5764_/B vssd1 vssd1 vccd1 vccd1 _5804_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_9_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_195 vssd1 vssd1 vccd1 vccd1 ci2406_z80_195/HI io_oeb[10] sky130_fd_sc_hd__conb_1
XFILLER_0_91_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3996_ _6071_/Q _6120_/Q vssd1 vssd1 vccd1 vccd1 _5370_/B sky130_fd_sc_hd__xor2_1
XANTENNA_fanout149_A _4725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5864__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5735_ _3959_/Y _5715_/B _5715_/Y _5734_/X vssd1 vssd1 vccd1 vccd1 _5735_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_29_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2947_ _3112_/A vssd1 vssd1 vccd1 vccd1 _3203_/A sky130_fd_sc_hd__inv_2
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5666_ _6066_/Q _5702_/A2 _5702_/B1 _5665_/X vssd1 vssd1 vccd1 vccd1 _5666_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_60_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5164__A1 _5164_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4617_ _4729_/A _4424_/D _4760_/B _4617_/D vssd1 vssd1 vccd1 vccd1 _4617_/X sky130_fd_sc_hd__and4bb_2
Xhold420 _5268_/X vssd1 vssd1 vccd1 vccd1 _6137_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5597_ _5596_/X _6060_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _5597_/X sky130_fd_sc_hd__mux2_1
Xhold442 _5774_/X vssd1 vssd1 vccd1 vccd1 _6220_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold453 _5727_/X vssd1 vssd1 vccd1 vccd1 _6207_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold431 _6192_/Q vssd1 vssd1 vccd1 vccd1 hold431/X sky130_fd_sc_hd__dlygate4sd3_1
X_4548_ _3556_/A _6058_/Q _4564_/S vssd1 vssd1 vccd1 vccd1 _4548_/X sky130_fd_sc_hd__mux2_1
Xhold464 _6217_/Q vssd1 vssd1 vccd1 vccd1 hold464/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 _5789_/X vssd1 vssd1 vccd1 vccd1 _6235_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold486 _6212_/Q vssd1 vssd1 vccd1 vccd1 hold486/X sky130_fd_sc_hd__dlygate4sd3_1
X_4479_ _5875_/B _5872_/B _4479_/C vssd1 vssd1 vccd1 vccd1 _4596_/S sky130_fd_sc_hd__and3_4
X_6218_ _6218_/CLK _6218_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6218_/Q sky130_fd_sc_hd__dfstp_1
Xhold497 _5233_/X vssd1 vssd1 vccd1 vccd1 hold497/X sky130_fd_sc_hd__dlygate4sd3_1
X_6149_ _6149_/CLK hold61/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__dfxtp_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4978__B2 _4976_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3132__B _5502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3323__A _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4969__A1 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4853__S _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3042__B _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3850_ _3851_/B _3851_/C _6139_/Q vssd1 vssd1 vccd1 vccd1 _3899_/A sky130_fd_sc_hd__o21ai_1
X_3781_ _3645_/X _3778_/B _3780_/X _3776_/X vssd1 vssd1 vccd1 vccd1 _3781_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3993__A _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5520_ _5519_/X _5514_/X _5670_/A vssd1 vssd1 vccd1 vccd1 _5520_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5146__A1 _3745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5451_ _5025_/A _5449_/X _5450_/X _3646_/X _5330_/B vssd1 vssd1 vccd1 vccd1 _5451_/X
+ sky130_fd_sc_hd__a2111o_1
X_4402_ _5250_/A _4410_/B _5317_/A vssd1 vssd1 vccd1 vccd1 _4402_/X sky130_fd_sc_hd__o21a_1
X_5382_ _6046_/Q _5380_/X _5381_/Y vssd1 vssd1 vccd1 vccd1 _5382_/X sky130_fd_sc_hd__o21a_1
X_4333_ _3880_/X hold264/X _4336_/S vssd1 vssd1 vccd1 vccd1 _6000_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4264_ hold239/X _4150_/X _4271_/S vssd1 vssd1 vccd1 vccd1 _5928_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3215_ _5838_/B _4759_/A vssd1 vssd1 vccd1 vccd1 _3215_/Y sky130_fd_sc_hd__nand2_1
X_6003_ _6152_/CLK _6003_/D vssd1 vssd1 vccd1 vccd1 _6003_/Q sky130_fd_sc_hd__dfxtp_1
X_4195_ _4195_/A _4195_/B vssd1 vssd1 vccd1 vccd1 _4195_/X sky130_fd_sc_hd__and2_1
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3146_ _3208_/B _4085_/B vssd1 vssd1 vccd1 vccd1 _3154_/B sky130_fd_sc_hd__nor2_1
X_3077_ _3507_/C _3187_/B _3182_/B _3070_/A vssd1 vssd1 vccd1 vccd1 _3077_/X sky130_fd_sc_hd__a31o_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5718_ hold578/X _5714_/Y _5717_/X _5023_/A vssd1 vssd1 vccd1 vccd1 _5718_/X sky130_fd_sc_hd__o22a_1
X_3979_ _3977_/X _3978_/X _4034_/S vssd1 vssd1 vccd1 vccd1 _3979_/X sky130_fd_sc_hd__mux2_2
XANTENNA__5137__A1 _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5649_ _5660_/B _5649_/B vssd1 vssd1 vccd1 vccd1 _5649_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__3699__A1 _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold250 _5972_/Q vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold261 _4326_/X vssd1 vssd1 vccd1 vccd1 _5994_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold294 _6019_/Q vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _5946_/Q vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold272 _3980_/X vssd1 vssd1 vccd1 vccd1 _5898_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4239__A _4239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3871__A1 _3582_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2982__A _6046_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4124__D _5424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5128__A1 _5164_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3318__A _4116_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4848__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3053__A _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput7 io_in[30] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
X_3000_ input9/X vssd1 vssd1 vccd1 vccd1 _6121_/D sky130_fd_sc_hd__inv_2
XANTENNA__5851__A2 _5836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4583__S _4598_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4951_ _6157_/Q _4950_/Y _5013_/S vssd1 vssd1 vccd1 vccd1 _4951_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3902_ _6071_/Q _3898_/A _5024_/B vssd1 vssd1 vccd1 vccd1 _3902_/X sky130_fd_sc_hd__o21a_1
X_4882_ _6059_/Q _6060_/Q _4854_/B _6061_/Q vssd1 vssd1 vccd1 vccd1 _4882_/X sky130_fd_sc_hd__a31o_1
X_3833_ _3597_/X _3832_/A _4253_/A2 vssd1 vssd1 vccd1 vccd1 _3833_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3378__B1 _4725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4612__A _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3764_ _6137_/Q _3764_/B _3764_/C vssd1 vssd1 vccd1 vccd1 _3765_/B sky130_fd_sc_hd__or3_1
XFILLER_0_6_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3695_ _3950_/B _3695_/B vssd1 vssd1 vccd1 vccd1 _3695_/Y sky130_fd_sc_hd__nor2_1
X_5503_ _3479_/A _4484_/A _5502_/X _4043_/C vssd1 vssd1 vccd1 vccd1 _5503_/X sky130_fd_sc_hd__o31a_1
X_5434_ _6231_/Q _5340_/Y _5433_/X _5341_/A vssd1 vssd1 vccd1 vccd1 _5434_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_2_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5365_ _5359_/X _5364_/X _5365_/S vssd1 vssd1 vccd1 vccd1 _5365_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4316_ _3930_/X hold104/X _4318_/S vssd1 vssd1 vccd1 vccd1 _4316_/X sky130_fd_sc_hd__mux2_1
X_5296_ hold23/X _5250_/B _5296_/S vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__mux2_1
X_4247_ _5927_/Q _3588_/X _3603_/X _6019_/Q vssd1 vssd1 vccd1 vccd1 _4247_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5842__A2 _5836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4178_ hold15/X _4253_/A2 _3786_/Y _4177_/Y _3671_/B vssd1 vssd1 vccd1 vccd1 _4178_/X
+ sky130_fd_sc_hd__o221a_1
X_3129_ _3148_/C _4398_/A _3113_/B _3128_/X vssd1 vssd1 vccd1 vccd1 _3129_/X sky130_fd_sc_hd__o31a_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3837__S _4035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold595_A _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4869__B1 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3541__B1 _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5530__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5294__B1 _5250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5247__B _5250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3480_ _4726_/C _3709_/B vssd1 vssd1 vccd1 vccd1 _4614_/C sky130_fd_sc_hd__or2_1
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5150_ _5150_/A _5150_/B _5150_/C vssd1 vssd1 vccd1 vccd1 _5150_/X sky130_fd_sc_hd__or3_1
XFILLER_0_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5081_ _3302_/A _3143_/Y _4036_/B _3457_/A vssd1 vssd1 vccd1 vccd1 _5081_/X sky130_fd_sc_hd__a31o_1
X_4101_ _3127_/B _4087_/X _4100_/X _4058_/X vssd1 vssd1 vccd1 vccd1 _4101_/X sky130_fd_sc_hd__a211o_1
X_4032_ hold3/X _4253_/A2 _3993_/Y _4031_/Y vssd1 vssd1 vccd1 vccd1 _4032_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4088__B2 _3694_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_1__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_leaf_9_wb_clk_i/A
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5037__B1 _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5588__A1 _6160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5983_ _6149_/CLK _5983_/D vssd1 vssd1 vccd1 vccd1 _5983_/Q sky130_fd_sc_hd__dfxtp_1
X_4934_ _6156_/Q _4933_/X _5013_/S vssd1 vssd1 vccd1 vccd1 _4934_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_19_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6111_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4260__A1 _5116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _3959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4865_ _4990_/A _4865_/B vssd1 vssd1 vccd1 vccd1 _4865_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_12 _6121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3816_ _6136_/Q _6137_/Q _6138_/Q vssd1 vssd1 vccd1 vccd1 _3912_/C sky130_fd_sc_hd__a21o_1
X_4796_ _4823_/C _4796_/B vssd1 vssd1 vccd1 vccd1 _4796_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_34 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3747_ hold74/A hold94/A _3982_/S vssd1 vssd1 vccd1 vccd1 _3748_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5760__B2 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3771__A0 _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3678_ _5116_/A _3674_/X _3677_/X vssd1 vssd1 vccd1 vccd1 _3678_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_100_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5417_ _5417_/A _5417_/B vssd1 vssd1 vccd1 vccd1 _5423_/A sky130_fd_sc_hd__xnor2_1
X_5348_ _5337_/X _5347_/X _5348_/S vssd1 vssd1 vccd1 vccd1 _5348_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3405__B _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5279_ _3890_/B _4219_/B _5289_/S vssd1 vssd1 vccd1 vccd1 _5279_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4079__A1 _4439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold343_A _6089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4951__S _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3794__C _3795_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5200__B1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5751__B2 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3762__B1 _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3817__A1 _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4490__A1 _5341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2980_ _2980_/A vssd1 vssd1 vccd1 vccd1 _2980_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4650_ hold520/X _5762_/A _4619_/X vssd1 vssd1 vccd1 vccd1 _4650_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_83_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4162__A _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput10 io_in[33] vssd1 vssd1 vccd1 vccd1 _6134_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3601_ _3988_/A _3616_/B _3982_/S vssd1 vssd1 vccd1 vccd1 _3601_/X sky130_fd_sc_hd__and3_4
X_4581_ hold552/X input7/X _4596_/S vssd1 vssd1 vccd1 vccd1 _4581_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3532_ _5362_/A _3532_/B vssd1 vssd1 vccd1 vccd1 _5837_/A sky130_fd_sc_hd__or2_2
X_6251_ _6251_/CLK _6251_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6251_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3463_ _3463_/A _4759_/A vssd1 vssd1 vccd1 vccd1 _4750_/A sky130_fd_sc_hd__nor2_2
X_6182_ _6238_/CLK _6182_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6182_/Q sky130_fd_sc_hd__dfrtp_1
X_5202_ _3978_/X _4241_/X _5198_/X _5201_/X _5185_/S _5116_/A vssd1 vssd1 vccd1 vccd1
+ _5202_/X sky130_fd_sc_hd__mux4_2
XANTENNA__5424__C _5424_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5133_ _5921_/Q _5200_/A2 _5200_/B1 _6029_/Q _5182_/S vssd1 vssd1 vccd1 vccd1 _5134_/C
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3225__B _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3394_ _4618_/C _5093_/B _5093_/A vssd1 vssd1 vccd1 vccd1 _3394_/Y sky130_fd_sc_hd__a21oi_1
X_5064_ hold17/X _3890_/B _5073_/S vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__mux2_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4015_ _4005_/A _5390_/B _4014_/X _4013_/A vssd1 vssd1 vccd1 vccd1 _4015_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4481__B2 _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5966_ _6034_/CLK _5966_/D vssd1 vssd1 vccd1 vccd1 _5966_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3036__A2 _5502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4917_ _6063_/Q _4918_/B vssd1 vssd1 vccd1 vccd1 _4948_/C sky130_fd_sc_hd__and2_1
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3895__B _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5897_ _6029_/CLK _5897_/D vssd1 vssd1 vccd1 vccd1 _5897_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_74_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4848_ _4847_/X _6058_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _4848_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5733__B2 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4779_ _4963_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _4779_/X sky130_fd_sc_hd__or2_1
XFILLER_0_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5497__A0 _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4946__S _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4067__A4 _4439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5724__B2 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3326__A _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5820_ hold380/X _5794_/Y _5819_/X _5794_/B vssd1 vssd1 vccd1 vccd1 _5820_/X sky130_fd_sc_hd__a22o_1
X_5751_ hold557/X _5741_/Y _5750_/X _5767_/A vssd1 vssd1 vccd1 vccd1 _5751_/X sky130_fd_sc_hd__o22a_1
X_2963_ _3382_/A vssd1 vssd1 vccd1 vccd1 _3513_/A sky130_fd_sc_hd__inv_4
X_4702_ _4676_/A _4676_/B _4676_/C _4687_/Y _4677_/A vssd1 vssd1 vccd1 vccd1 _4703_/C
+ sky130_fd_sc_hd__a311o_1
X_5682_ _5682_/A _5682_/B _5682_/C vssd1 vssd1 vccd1 vccd1 _5682_/X sky130_fd_sc_hd__or3_1
X_4633_ hold454/X _4612_/B _4632_/X _4474_/X vssd1 vssd1 vccd1 vccd1 _4633_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_44_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold602 _5488_/X vssd1 vssd1 vccd1 vccd1 _6179_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__6040__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4564_ _4061_/A _6059_/Q _4564_/S vssd1 vssd1 vccd1 vccd1 _4564_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold635 _6159_/Q vssd1 vssd1 vccd1 vccd1 hold635/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold624 _5309_/X vssd1 vssd1 vccd1 vccd1 _6157_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3515_ _6164_/Q _3514_/Y _3508_/A vssd1 vssd1 vccd1 vccd1 _3515_/X sky130_fd_sc_hd__a21o_1
Xhold613 _3519_/X vssd1 vssd1 vccd1 vccd1 _6170_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6234_ _6235_/CLK _6234_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6234_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5479__A0 _6179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold646 _5227_/X vssd1 vssd1 vccd1 vccd1 _6125_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 _6168_/Q vssd1 vssd1 vccd1 vccd1 hold657/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4495_ hold149/X _5997_/Q hold90/X _5958_/Q _4272_/B _5076_/A0 vssd1 vssd1 vccd1
+ vccd1 _4495_/X sky130_fd_sc_hd__mux4_1
X_3446_ _3446_/A _4043_/C vssd1 vssd1 vccd1 vccd1 _4046_/B sky130_fd_sc_hd__nand2_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6165_ _6171_/CLK _6165_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6165_/Q sky130_fd_sc_hd__dfrtp_4
X_3377_ _4497_/S _6163_/Q _6164_/Q _4725_/B vssd1 vssd1 vccd1 vccd1 _3377_/X sky130_fd_sc_hd__o31a_2
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _5116_/A _5116_/B _5116_/C vssd1 vssd1 vccd1 vccd1 _5116_/X sky130_fd_sc_hd__and3_1
X_6096_ _6102_/CLK _6096_/D vssd1 vssd1 vccd1 vccd1 _6096_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5047_ _3648_/Y _5045_/X _5046_/X _5026_/Y _5044_/X vssd1 vssd1 vccd1 vccd1 _5047_/X
+ sky130_fd_sc_hd__o311a_1
Xclkbuf_leaf_34_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6247_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3257__A2 _4759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4454__A1 _6048_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5597__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5949_ _6033_/CLK _5949_/D vssd1 vssd1 vccd1 vccd1 _5949_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6128__RESET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5167__C1 _3594_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2985__A _6157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4693__A1 _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5361__A _5363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3879__S0 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4540__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3653__C1 _4391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5300__S _5305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5158__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3300_ _4765_/A _4390_/A vssd1 vssd1 vccd1 vccd1 _3301_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4280_ hold72/X _4226_/X _4282_/S vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__mux2_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3439_/B _3221_/X _3215_/Y vssd1 vssd1 vccd1 vccd1 _3231_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_39_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _4070_/B _4036_/B vssd1 vssd1 vccd1 vccd1 _3622_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_55_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3503__B _6047_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4436__B2 _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3093_ _3112_/A _4094_/D _3125_/C vssd1 vssd1 vccd1 vccd1 _5424_/A sky130_fd_sc_hd__or3_4
XFILLER_0_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5803_ _6238_/Q _5352_/A _5457_/A hold437/X vssd1 vssd1 vccd1 vccd1 _5803_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_64_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_196 vssd1 vssd1 vccd1 vccd1 ci2406_z80_196/HI io_oeb[11] sky130_fd_sc_hd__conb_1
Xci2406_z80_185 vssd1 vssd1 vccd1 vccd1 ci2406_z80_185/HI io_oeb[0] sky130_fd_sc_hd__conb_1
X_3995_ _5046_/A _3995_/B vssd1 vssd1 vccd1 vccd1 _3998_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_9_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5734_ _4116_/Y _4865_/B _4579_/Y _5762_/C vssd1 vssd1 vccd1 vccd1 _5734_/X sky130_fd_sc_hd__o22a_1
X_2946_ _4077_/A vssd1 vssd1 vccd1 vccd1 _5220_/A sky130_fd_sc_hd__inv_2
X_5665_ _6184_/Q _6200_/Q _5701_/S vssd1 vssd1 vccd1 vccd1 _5665_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4616_ _4772_/D _4616_/B vssd1 vssd1 vccd1 vccd1 _4617_/D sky130_fd_sc_hd__nor2_1
Xhold410 _6116_/Q vssd1 vssd1 vccd1 vccd1 _2978_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5596_ _4119_/B _5595_/X _4865_/Y vssd1 vssd1 vccd1 vccd1 _5596_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_4_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold443 _6233_/Q vssd1 vssd1 vccd1 vccd1 hold443/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold454 _6063_/Q vssd1 vssd1 vccd1 vccd1 hold454/X sky130_fd_sc_hd__clkbuf_2
Xhold421 _6193_/Q vssd1 vssd1 vccd1 vccd1 hold421/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold432 _5574_/X vssd1 vssd1 vccd1 vccd1 _6192_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4547_ _4547_/A _4547_/B vssd1 vssd1 vccd1 vccd1 _4547_/Y sky130_fd_sc_hd__xnor2_2
Xhold476 _6225_/Q vssd1 vssd1 vccd1 vccd1 hold476/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold465 _5760_/X vssd1 vssd1 vccd1 vccd1 _6217_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 _5745_/X vssd1 vssd1 vccd1 vccd1 _6212_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4478_ _4478_/A hold46/X vssd1 vssd1 vccd1 vccd1 _4479_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6217_ _6218_/CLK _6217_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6217_/Q sky130_fd_sc_hd__dfstp_2
Xhold498 _5234_/X vssd1 vssd1 vccd1 vccd1 _6128_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4496__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3429_ _3154_/B _3428_/Y _5489_/D vssd1 vssd1 vccd1 vccd1 _3429_/Y sky130_fd_sc_hd__o21ai_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6148_ _6148_/CLK _6148_/D vssd1 vssd1 vccd1 vccd1 _6148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5624__B1 _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6079_ _6170_/CLK _6079_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6079_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5155__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4666__A1 _4522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4210__S0 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3604__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4435__A _5424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5091__B2 _4433_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3780_ _3650_/X _5387_/A _3779_/X _6115_/Q vssd1 vssd1 vccd1 vccd1 _3780_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_6_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5450_ _5033_/A _3840_/B _5026_/A _6176_/Q vssd1 vssd1 vccd1 vccd1 _5450_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_54_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5146__A2 _5105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4401_ _3527_/A _4400_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _6040_/D sky130_fd_sc_hd__mux2_1
X_5381_ _2958_/Y _6046_/Q _6073_/Q vssd1 vssd1 vccd1 vccd1 _5381_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4332_ _3836_/X hold194/X _4336_/S vssd1 vssd1 vccd1 vccd1 _4332_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4263_ _4263_/A _4364_/B vssd1 vssd1 vccd1 vccd1 _4271_/S sky130_fd_sc_hd__nor2_4
XANTENNA__4657__A1 _4943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3214_ _4398_/B _4765_/A vssd1 vssd1 vccd1 vccd1 _4043_/C sky130_fd_sc_hd__or2_4
X_6002_ _6010_/CLK _6002_/D vssd1 vssd1 vccd1 vccd1 _6002_/Q sky130_fd_sc_hd__dfxtp_1
X_4194_ hold124/X _4193_/X _4262_/S vssd1 vssd1 vccd1 vccd1 _4194_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4409__A1 _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4409__B2 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3145_ _3777_/A _5356_/A _3643_/A vssd1 vssd1 vccd1 vccd1 _4085_/B sky130_fd_sc_hd__nand3b_4
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3076_ _3511_/D _3063_/X _4117_/C _3074_/Y _4118_/B vssd1 vssd1 vccd1 vccd1 _4727_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5082__B2 _4391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout161_A _5936_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ hold260/X hold284/X hold161/X hold179/X _5179_/S _3740_/S vssd1 vssd1 vccd1
+ vccd1 _3978_/X sky130_fd_sc_hd__mux4_2
X_5717_ _3664_/X _5715_/B _5715_/Y _5716_/X vssd1 vssd1 vccd1 vccd1 _5717_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_45_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5648_ _6198_/Q _5685_/B _5639_/X vssd1 vssd1 vccd1 vccd1 _5649_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5579_ _5578_/X hold421/X _5705_/S vssd1 vssd1 vccd1 vccd1 _5579_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3699__A2 _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold251 _4309_/X vssd1 vssd1 vccd1 vccd1 _5972_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 _5961_/Q vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold240 _5894_/Q vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3127__C _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold295 _4354_/X vssd1 vssd1 vccd1 vccd1 _6019_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _5979_/Q vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold284 _5912_/Q vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_hold373_A _6117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout74_A _4239_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3143__B _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4820__A1 _4819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3084__B1 _4486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 io_in[31] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4864__S _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_0__f_wb_clk_i clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _5978_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4950_ _4966_/B _4950_/B vssd1 vssd1 vccd1 vccd1 _4950_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_59_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4881_ _4879_/B _4880_/X _4963_/A vssd1 vssd1 vccd1 vccd1 _4881_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3901_ _3900_/A _3900_/B _3848_/B vssd1 vssd1 vccd1 vccd1 _3901_/X sky130_fd_sc_hd__o21a_1
X_3832_ _3832_/A vssd1 vssd1 vccd1 vccd1 _3832_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3378__A1 _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4612__B _4612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3763_ _5024_/A _3765_/A vssd1 vssd1 vccd1 vccd1 _3763_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__3509__A _3517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5502_ _5502_/A _5502_/B _5502_/C _5502_/D vssd1 vssd1 vccd1 vccd1 _5502_/X sky130_fd_sc_hd__or4_1
X_3694_ _3777_/A _4735_/A _3694_/C vssd1 vssd1 vccd1 vccd1 _3695_/B sky130_fd_sc_hd__and3_1
X_5433_ _5457_/A _5433_/B _5433_/C vssd1 vssd1 vccd1 vccd1 _5433_/X sky130_fd_sc_hd__or3_1
X_5364_ _5033_/A _5448_/B _5025_/A _6173_/Q vssd1 vssd1 vccd1 vccd1 _5364_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_2_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4878__A1 _4877_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4315_ _3880_/X hold205/X _4318_/S vssd1 vssd1 vccd1 vccd1 _5984_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5295_ hold48/X _5294_/X _5875_/A vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__mux2_1
X_4246_ _5944_/Q _3611_/X _3613_/X _5935_/Q _4245_/X vssd1 vssd1 vccd1 vccd1 _4249_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4177_ _4223_/A _5055_/A vssd1 vssd1 vccd1 vccd1 _4177_/Y sky130_fd_sc_hd__nor2_1
X_3128_ _3210_/A _3203_/B _4485_/A _3777_/A vssd1 vssd1 vccd1 vccd1 _3128_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_96_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_42_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3059_ _3556_/A _4061_/A vssd1 vssd1 vccd1 vccd1 _4406_/A sky130_fd_sc_hd__nand2_2
XANTENNA__4802__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4522__B _4522_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold588_A _5918_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3601__B _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3329__A _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3780__B2 _6115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5080_ _5502_/A _5080_/B vssd1 vssd1 vccd1 vccd1 _5080_/Y sky130_fd_sc_hd__nor2_1
X_4100_ _4061_/A _4124_/B _3143_/Y _4044_/B _3097_/Y vssd1 vssd1 vccd1 vccd1 _4100_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5285__A1 _6160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5285__B2 _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4031_ _3597_/X _4030_/A _3539_/Y vssd1 vssd1 vccd1 vccd1 _4031_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__3999__A _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3296__B1 _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3511__B _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5982_ _6010_/CLK _5982_/D vssd1 vssd1 vccd1 vccd1 _5982_/Q sky130_fd_sc_hd__dfxtp_1
X_4933_ _6064_/Q _4948_/C vssd1 vssd1 vccd1 vccd1 _4933_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4548__A0 _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_13 _6121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4864_ hold347/X _4863_/X _4927_/S vssd1 vssd1 vccd1 vccd1 _4864_/X sky130_fd_sc_hd__mux2_1
X_3815_ _5024_/A _6138_/Q _6116_/Q _3848_/B _3814_/X vssd1 vssd1 vccd1 vccd1 _5375_/B
+ sky130_fd_sc_hd__o41a_2
X_4795_ _6054_/Q _5013_/S _6055_/Q vssd1 vssd1 vccd1 vccd1 _4796_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_35 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_24 _6094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout124_A _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3746_ _3620_/X _3732_/B _3730_/X vssd1 vssd1 vccd1 vccd1 _3759_/A sky130_fd_sc_hd__a21o_1
X_5416_ _6161_/Q _6160_/Q vssd1 vssd1 vccd1 vccd1 _5417_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3673__S _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3677_ _5209_/A _3677_/B _3677_/C vssd1 vssd1 vccd1 vccd1 _3677_/X sky130_fd_sc_hd__or3_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_100_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4720__B1 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5347_ _6172_/Q _5342_/Y _5346_/X _3377_/X vssd1 vssd1 vccd1 vccd1 _5347_/X sky130_fd_sc_hd__o22a_1
X_5278_ _5245_/A hold416/X _5245_/Y _5277_/X vssd1 vssd1 vccd1 vccd1 _5278_/X sky130_fd_sc_hd__a22o_1
X_4229_ hold64/X _3611_/X _3613_/X hold80/X _4228_/X vssd1 vssd1 vccd1 vccd1 _4232_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3149__A _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2988__A _6160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3514__A1 _3252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3817__A2 _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5303__S _5305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5019__A1 _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4490__A2 _4598_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4778__A0 _6188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput11 io_in[34] vssd1 vssd1 vccd1 vccd1 _3383_/B sky130_fd_sc_hd__buf_4
XFILLER_0_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4625__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4580_ hold552/X _4612_/B _4579_/Y _4474_/X vssd1 vssd1 vccd1 vccd1 _4580_/X sky130_fd_sc_hd__a22o_1
X_3600_ _3968_/A _3983_/S _3982_/S vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__or3_1
XANTENNA__3059__A _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3531_ _6073_/Q _5460_/S vssd1 vssd1 vccd1 vccd1 _3531_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_52_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3493__S _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6250_ _6251_/CLK _6250_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6250_/Q sky130_fd_sc_hd__dfrtp_1
X_3462_ _4478_/A _3525_/C _3715_/B vssd1 vssd1 vccd1 vccd1 _3462_/Y sky130_fd_sc_hd__o21ai_1
X_6181_ _6238_/CLK _6181_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6181_/Q sky130_fd_sc_hd__dfrtp_1
X_5201_ _5201_/A _5201_/B vssd1 vssd1 vccd1 vccd1 _5201_/X sky130_fd_sc_hd__or2_1
XANTENNA__3506__B _3517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3505__A1 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3393_ _3389_/B _4457_/B _3392_/Y _3388_/B vssd1 vssd1 vccd1 vccd1 _3393_/X sky130_fd_sc_hd__a22o_1
X_5132_ _6013_/Q _5200_/A2 _5200_/B1 _5946_/Q _4256_/S vssd1 vssd1 vccd1 vccd1 _5134_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5258__B2 _5257_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5258__A1 _5245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5063_ hold13/X _3875_/B _5073_/S vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__mux2_1
XFILLER_0_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4014_ _4014_/A _4014_/B vssd1 vssd1 vccd1 vccd1 _4014_/X sky130_fd_sc_hd__or2_1
XFILLER_0_90_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5965_ _6110_/CLK _5965_/D vssd1 vssd1 vccd1 vccd1 _5965_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4916_ _4104_/B _4914_/X _4915_/X _4999_/A1 vssd1 vssd1 vccd1 vccd1 _4916_/X sky130_fd_sc_hd__o211a_1
X_5896_ _6029_/CLK _5896_/D vssd1 vssd1 vccd1 vccd1 _5896_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4847_ _4119_/B _4846_/X _4836_/Y vssd1 vssd1 vccd1 vccd1 _4847_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_7_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4778_ _6188_/Q _6054_/Q _5216_/A vssd1 vssd1 vccd1 vccd1 _4778_/X sky130_fd_sc_hd__mux2_1
X_3729_ _5259_/A vssd1 vssd1 vccd1 vccd1 _3729_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_100_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4962__S _5216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4224__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_wb_clk_i _5978_/CLK vssd1 vssd1 vccd1 vccd1 _6146_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_0_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4448__C1 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3996__B _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4215__A2 _3588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5750_ _3785_/Y _5771_/S _5742_/Y _5749_/X vssd1 vssd1 vccd1 vccd1 _5750_/X sky130_fd_sc_hd__o22a_1
X_2962_ _3461_/A vssd1 vssd1 vccd1 vccd1 _5362_/A sky130_fd_sc_hd__inv_2
X_5681_ _5682_/A _5682_/B _5682_/C vssd1 vssd1 vccd1 vccd1 _5681_/Y sky130_fd_sc_hd__o21ai_1
X_4701_ _4716_/A _4701_/B vssd1 vssd1 vccd1 vccd1 _4705_/A sky130_fd_sc_hd__nand2_1
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4632_ _4632_/A _4632_/B vssd1 vssd1 vccd1 vccd1 _4632_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold603 _6237_/Q vssd1 vssd1 vccd1 vccd1 hold603/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4563_ _4563_/A _4563_/B vssd1 vssd1 vccd1 vccd1 _4563_/Y sky130_fd_sc_hd__xnor2_1
Xhold636 _6161_/Q vssd1 vssd1 vccd1 vccd1 hold636/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__4112__S _4115_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold625 _6255_/Q vssd1 vssd1 vccd1 vccd1 hold625/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3514_ _3252_/B _3508_/C _3513_/C vssd1 vssd1 vccd1 vccd1 _3514_/Y sky130_fd_sc_hd__o21ai_1
Xhold614 _6073_/Q vssd1 vssd1 vccd1 vccd1 hold614/X sky130_fd_sc_hd__dlygate4sd3_1
X_4494_ hold132/X hold191/X hold91/X hold208/X _4272_/B _5076_/A0 vssd1 vssd1 vccd1
+ vccd1 _4494_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_100_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6233_ _6233_/CLK _6233_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6233_/Q sky130_fd_sc_hd__dfstp_1
X_3445_ _3298_/A _3296_/X _5838_/C _3228_/B _3444_/X vssd1 vssd1 vccd1 vccd1 _3445_/X
+ sky130_fd_sc_hd__a221o_1
Xhold647 _5936_/Q vssd1 vssd1 vccd1 vccd1 hold647/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold658 _6005_/Q vssd1 vssd1 vccd1 vccd1 hold658/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3951__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3376_/A _3376_/B _3376_/C hold34/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__or4_1
X_6164_ _6171_/CLK _6164_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6164_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3252__A _6050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5115_ _3595_/X _5209_/A _5185_/S _5114_/X vssd1 vssd1 vccd1 vccd1 _5115_/X sky130_fd_sc_hd__a211o_1
X_6095_ _6256_/CLK _6095_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6095_/Q sky130_fd_sc_hd__dfrtp_1
X_5046_ _5046_/A _6139_/Q _6140_/Q _6141_/Q vssd1 vssd1 vccd1 vccd1 _5046_/X sky130_fd_sc_hd__or4_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4454__A2 _3517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5948_ _6035_/CLK _5948_/D vssd1 vssd1 vccd1 vccd1 _5948_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3414__B1 _5424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5879_ _3112_/A _5875_/X _5876_/Y _5878_/X vssd1 vssd1 vccd1 vccd1 _5879_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5167__B1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5626__B _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4914__A0 _6197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3717__A1 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4693__A2 _4620_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3162__A _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3879__S1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3653__B1 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5158__B1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3708__A1 _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4867__S _5216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _3200_/X _3220_/X _3229_/X _3164_/Y vssd1 vssd1 vccd1 vccd1 _3234_/C sky130_fd_sc_hd__a31o_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _4413_/A _3160_/X _4415_/A vssd1 vssd1 vccd1 vccd1 _3234_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__3503__C _3503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5633__A1 _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3092_ _4417_/B _3125_/C vssd1 vssd1 vccd1 vccd1 _4446_/A sky130_fd_sc_hd__or2_2
XANTENNA__3800__A _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5802_ hold603/X _5801_/X _5832_/S vssd1 vssd1 vccd1 vccd1 _6237_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_71_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_197 vssd1 vssd1 vccd1 vccd1 ci2406_z80_197/HI io_oeb[12] sky130_fd_sc_hd__conb_1
Xci2406_z80_186 vssd1 vssd1 vccd1 vccd1 ci2406_z80_186/HI io_oeb[1] sky130_fd_sc_hd__conb_1
XFILLER_0_57_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3994_ _3935_/Y _3936_/X _3939_/B vssd1 vssd1 vccd1 vccd1 _3995_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5733_ hold569/X _5714_/Y _5732_/X _5023_/A vssd1 vssd1 vccd1 vccd1 _5733_/X sky130_fd_sc_hd__o22a_1
X_5664_ _5664_/A _5664_/B vssd1 vssd1 vccd1 vccd1 _5664_/Y sky130_fd_sc_hd__xnor2_1
X_5595_ _5594_/X _6060_/Q _5595_/S vssd1 vssd1 vccd1 vccd1 _5595_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4615_ _4728_/C _4615_/B _4727_/B _4615_/D vssd1 vssd1 vccd1 vccd1 _4616_/B sky130_fd_sc_hd__or4_1
Xhold411 _5164_/X vssd1 vssd1 vccd1 vccd1 _6116_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold400 _6138_/Q vssd1 vssd1 vccd1 vccd1 hold400/X sky130_fd_sc_hd__dlygate4sd3_1
X_4546_ _4529_/B _4531_/B _4529_/A vssd1 vssd1 vccd1 vccd1 _4547_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3247__A _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold444 _5787_/X vssd1 vssd1 vccd1 vccd1 _6233_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold433 _6234_/Q vssd1 vssd1 vccd1 vccd1 hold433/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 _5587_/X vssd1 vssd1 vccd1 vccd1 _6193_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 _6200_/Q vssd1 vssd1 vccd1 vccd1 _5658_/A sky130_fd_sc_hd__buf_1
Xhold477 _5779_/X vssd1 vssd1 vccd1 vccd1 _6225_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold455 _4637_/X vssd1 vssd1 vccd1 vccd1 _6063_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4477_ _4478_/A hold300/X _5498_/A _3252_/B vssd1 vssd1 vccd1 vccd1 _5872_/B sky130_fd_sc_hd__a211o_1
Xhold488 _6223_/Q vssd1 vssd1 vccd1 vccd1 hold488/X sky130_fd_sc_hd__dlygate4sd3_1
X_6216_ _6218_/CLK _6216_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6216_/Q sky130_fd_sc_hd__dfstp_1
Xhold499 _6162_/Q vssd1 vssd1 vccd1 vccd1 _5319_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3428_ _4021_/B _3428_/B vssd1 vssd1 vccd1 vccd1 _3428_/Y sky130_fd_sc_hd__nor2_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _5220_/A _3370_/B _3370_/C vssd1 vssd1 vccd1 vccd1 _3368_/C sky130_fd_sc_hd__and3_1
X_6147_ _6152_/CLK hold75/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__3883__B1 _3615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5624__A1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6078_ _6086_/CLK _6078_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6078_/Q sky130_fd_sc_hd__dfrtp_1
X_5029_ _5373_/A _5373_/B _5029_/C vssd1 vssd1 vccd1 vccd1 _5029_/X sky130_fd_sc_hd__or3_1
XANTENNA__6293__A _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5356__B _6165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5312__A0 input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4666__A2 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5863__B2 _5245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4210__S1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3604__B _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5311__S _5313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4400_ _5259_/B _4410_/B _5317_/A vssd1 vssd1 vccd1 vccd1 _4400_/X sky130_fd_sc_hd__o21a_1
X_5380_ _3647_/C _5371_/Y _5378_/Y _5379_/X vssd1 vssd1 vccd1 vccd1 _5380_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4597__S _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4331_ _3789_/X hold185/X _4336_/S vssd1 vssd1 vccd1 vccd1 _5998_/D sky130_fd_sc_hd__mux2_1
X_4262_ hold211/X _4261_/X _4262_/S vssd1 vssd1 vccd1 vccd1 _4262_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5854__A1 _3832_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6001_ _6006_/CLK _6001_/D vssd1 vssd1 vccd1 vccd1 _6001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3213_ _4398_/B _4765_/A vssd1 vssd1 vccd1 vccd1 _4759_/A sky130_fd_sc_hd__nor2_4
X_4193_ _4191_/X _4192_/X _4242_/S vssd1 vssd1 vccd1 vccd1 _4193_/X sky130_fd_sc_hd__mux2_2
X_3144_ _3694_/C _4061_/C vssd1 vssd1 vccd1 vccd1 _4036_/B sky130_fd_sc_hd__nor2_8
X_3075_ _4117_/B _4117_/C vssd1 vssd1 vccd1 vccd1 _4118_/B sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_32_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_82_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3977_ hold1/X _4253_/A2 _3960_/Y _3976_/Y vssd1 vssd1 vccd1 vccd1 _3977_/X sky130_fd_sc_hd__o22a_1
X_5716_ _4119_/A _4779_/B _4473_/Y _5762_/C vssd1 vssd1 vccd1 vccd1 _5716_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_45_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5647_ _5647_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5660_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5578_ _5577_/X _6059_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _5578_/X sky130_fd_sc_hd__mux2_1
Xhold230 _6017_/Q vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _6029_/Q vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
X_4529_ _4529_/A _4529_/B vssd1 vssd1 vccd1 vccd1 _4531_/A sky130_fd_sc_hd__nand2_1
Xhold241 _5964_/Q vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 _3371_/X vssd1 vssd1 vccd1 vccd1 _5979_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 _5957_/Q vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4300__S _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold285 _6010_/Q vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 _6003_/Q vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout67_A _4926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5781__A0 _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5306__S _5313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3615__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5022__B1_N _5052_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput9 io_in[32] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__3350__A _5314_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4880__S _5216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4880_ _6195_/Q _6061_/Q _5216_/A vssd1 vssd1 vccd1 vccd1 _4880_/X sky130_fd_sc_hd__mux2_1
X_3900_ _3900_/A _3900_/B vssd1 vssd1 vccd1 vccd1 _3900_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_86_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3831_ _3830_/X _3805_/B _3958_/S vssd1 vssd1 vccd1 vccd1 _3832_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_52_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3762_ _3764_/B _3764_/C _6137_/Q vssd1 vssd1 vccd1 vccd1 _3765_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3509__B _3517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5501_ _2957_/Y _4618_/A _4043_/C _4460_/A vssd1 vssd1 vccd1 vccd1 _5501_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_42_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3693_ _3648_/A _5404_/B _5395_/B _3920_/A vssd1 vssd1 vccd1 vccd1 _3693_/X sky130_fd_sc_hd__a22o_1
X_5432_ _6175_/Q _5352_/Y _5354_/B _2989_/Y vssd1 vssd1 vccd1 vccd1 _5433_/C sky130_fd_sc_hd__o211a_1
XFILLER_0_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5363_ _5487_/S _5363_/B _5363_/C vssd1 vssd1 vccd1 vccd1 _5363_/X sky130_fd_sc_hd__and3_1
X_4314_ _3836_/X hold237/X _4318_/S vssd1 vssd1 vccd1 vccd1 _5983_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_10_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3525__A _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5294_ _3275_/B _5250_/B _5250_/A vssd1 vssd1 vccd1 vccd1 _5294_/X sky130_fd_sc_hd__a21o_1
X_4245_ _6027_/Q _3599_/X _3601_/X _5972_/Q vssd1 vssd1 vccd1 vccd1 _4245_/X sky130_fd_sc_hd__a22o_1
X_4176_ _4195_/A _4176_/B vssd1 vssd1 vccd1 vccd1 _5055_/A sky130_fd_sc_hd__xnor2_1
X_3127_ _6252_/Q _3127_/B _3277_/A _3178_/C vssd1 vssd1 vccd1 vccd1 _3154_/A sky130_fd_sc_hd__and4_1
XFILLER_0_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3058_ _4735_/A _3694_/C vssd1 vssd1 vccd1 vccd1 _4391_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4566__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5294__A2 _5250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3170__A _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5809__A1 _6239_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5809__B2 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4030_ _4030_/A vssd1 vssd1 vccd1 vccd1 _4030_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3999__B _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3296__A1 _4451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3048__A1 _3193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5981_ _6144_/CLK _5981_/D vssd1 vssd1 vccd1 vccd1 _5981_/Q sky130_fd_sc_hd__dfxtp_1
X_4932_ _4928_/B _4931_/X _4963_/A vssd1 vssd1 vccd1 vccd1 _4932_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_14 _6121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4863_ _4862_/X _6059_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _4863_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4115__S _4115_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_25 _6089_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3814_ _3811_/X _3812_/Y _3813_/X vssd1 vssd1 vccd1 vccd1 _3814_/X sky130_fd_sc_hd__a21o_1
X_4794_ _6054_/Q _6055_/Q _5013_/S vssd1 vssd1 vccd1 vccd1 _4823_/C sky130_fd_sc_hd__and3_1
XFILLER_0_15_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3745_ _5116_/A _3741_/X _3744_/X vssd1 vssd1 vccd1 vccd1 _3745_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3220__A1 _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5415_ _6157_/Q _6156_/Q vssd1 vssd1 vccd1 vccd1 _5417_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout117_A _5360_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3676_ _5997_/Q _3591_/A _3740_/S _5958_/Q _4256_/S vssd1 vssd1 vccd1 vccd1 _3677_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_100_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_28_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6238_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5346_ _5705_/S _5344_/X _5345_/Y _5340_/Y hold456/X vssd1 vssd1 vccd1 vccd1 _5346_/X
+ sky130_fd_sc_hd__o32a_1
X_5277_ _5248_/Y _5274_/X _5276_/X vssd1 vssd1 vccd1 vccd1 _5277_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4228_ _6026_/Q _3599_/X _3601_/X _5971_/Q vssd1 vssd1 vccd1 vccd1 _4228_/X sky130_fd_sc_hd__a22o_1
X_4159_ _4219_/A _4159_/B vssd1 vssd1 vccd1 vccd1 _4174_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5629__B _5629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5200__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3149__B _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3817__A3 _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3612__B _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4490__A3 _4612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 io_in[35] vssd1 vssd1 vccd1 vccd1 _3001_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__4625__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3059__B _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3530_ _6072_/Q _6070_/Q _5333_/B vssd1 vssd1 vccd1 vccd1 _5460_/S sky130_fd_sc_hd__nand3_4
XFILLER_0_52_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3461_ _3461_/A _3503_/C vssd1 vssd1 vccd1 vccd1 _3525_/C sky130_fd_sc_hd__nor2_1
X_6180_ _6238_/CLK _6180_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6180_/Q sky130_fd_sc_hd__dfrtp_1
X_5200_ _5926_/Q _5200_/A2 _5200_/B1 _6034_/Q _5182_/S vssd1 vssd1 vccd1 vccd1 _5201_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4163__C1 _3671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3392_ _3392_/A _4457_/B vssd1 vssd1 vccd1 vccd1 _3392_/Y sky130_fd_sc_hd__nor2_1
X_5131_ _6205_/Q _5106_/Y _5122_/Y _6189_/Q _5130_/X vssd1 vssd1 vccd1 vccd1 _5139_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_58_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5062_ hold19/X _3800_/B _5073_/S vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__mux2_1
XANTENNA__3803__A _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4013_ _4013_/A _4014_/B vssd1 vssd1 vccd1 vccd1 _5390_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4618__B _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3241__C _6174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3949__S _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5430__A2 _5352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5964_ _6152_/CLK _5964_/D vssd1 vssd1 vccd1 vccd1 _5964_/Q sky130_fd_sc_hd__dfxtp_1
X_4915_ _4963_/A _4915_/B vssd1 vssd1 vccd1 vccd1 _4915_/X sky130_fd_sc_hd__or2_1
XFILLER_0_74_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5895_ _6152_/CLK _5895_/D vssd1 vssd1 vccd1 vccd1 _5895_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3441__A1 _5838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4846_ _6058_/Q _5702_/A2 _5607_/B1 _4845_/X vssd1 vssd1 vccd1 vccd1 _4846_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_47_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5194__A1 _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4777_ _6054_/Q _5013_/S vssd1 vssd1 vccd1 vccd1 _4777_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3728_ _3730_/B _3730_/C vssd1 vssd1 vccd1 vccd1 _5259_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3659_ _3657_/A _3645_/X _3648_/A _5404_/A vssd1 vssd1 vccd1 vccd1 _3659_/X sky130_fd_sc_hd__a22o_1
X_5329_ _6074_/Q _3496_/X _3646_/X vssd1 vssd1 vccd1 vccd1 _5365_/S sky130_fd_sc_hd__a21o_2
XANTENNA__6296__A _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3713__A _3713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold181_A _6166_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4393__C1 _4737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3499__A1 _6127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3623__A _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4999__B2 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4999__A1 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2961_ _6127_/Q vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__inv_2
XANTENNA__3423__B2 _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3423__A1 _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4620__B1 _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5680_ _5664_/A _5664_/B _5659_/A vssd1 vssd1 vccd1 vccd1 _5682_/C sky130_fd_sc_hd__o21a_1
X_4700_ _4715_/A _4700_/B vssd1 vssd1 vccd1 vccd1 _4701_/B sky130_fd_sc_hd__or2_1
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4631_ _4647_/A _4631_/B vssd1 vssd1 vccd1 vccd1 _4632_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_71_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4562_ _4545_/B _4547_/B _4545_/A vssd1 vssd1 vccd1 vccd1 _4563_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3726__A2 _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4493_ _4589_/S _4493_/B vssd1 vssd1 vccd1 vccd1 _4498_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_52_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold626 _5883_/X vssd1 vssd1 vccd1 vccd1 _6255_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold604 _6127_/Q vssd1 vssd1 vccd1 vccd1 hold604/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3517__B _3517_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3513_ _3513_/A _6170_/Q _3513_/C vssd1 vssd1 vccd1 vccd1 _3516_/C sky130_fd_sc_hd__or3_1
Xhold615 _4748_/X vssd1 vssd1 vccd1 vccd1 _6073_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold637 _6154_/Q vssd1 vssd1 vccd1 vccd1 hold637/X sky130_fd_sc_hd__dlygate4sd3_1
X_6232_ _6247_/CLK _6232_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6232_/Q sky130_fd_sc_hd__dfstp_1
XFILLER_0_69_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3444_ _4045_/A _3713_/B _3408_/X _4451_/C vssd1 vssd1 vccd1 vccd1 _3444_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold648 _6112_/Q vssd1 vssd1 vccd1 vccd1 hold648/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold659 _3678_/X vssd1 vssd1 vccd1 vccd1 hold659/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ hold42/A hold56/A hold33/X _5979_/Q _3353_/X vssd1 vssd1 vccd1 vccd1 hold34/A
+ sky130_fd_sc_hd__o41a_1
X_6163_ _6171_/CLK _6163_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6163_/Q sky130_fd_sc_hd__dfrtp_1
X_6094_ _6206_/CLK _6094_/D vssd1 vssd1 vccd1 vccd1 _6094_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5116_/A _5114_/B _5114_/C vssd1 vssd1 vccd1 vccd1 _5114_/X sky130_fd_sc_hd__and3_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5404_/A _5404_/B _5403_/A _5403_/B vssd1 vssd1 vccd1 vccd1 _5045_/X sky130_fd_sc_hd__or4_1
XANTENNA__3252__B _3252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5100__A1 _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5651__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout184_A input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5947_ _6014_/CLK _5947_/D vssd1 vssd1 vccd1 vccd1 _5947_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3965__A2 _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5878_ input2/X _5890_/B vssd1 vssd1 vccd1 vccd1 _5878_/X sky130_fd_sc_hd__and2_1
X_4829_ _4829_/A _4829_/B _4829_/C vssd1 vssd1 vccd1 vccd1 _4829_/X sky130_fd_sc_hd__or3_1
XFILLER_0_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_43_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6123_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4303__S _4309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold396_A _6088_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3162__B _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5642__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5309__S _5313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4905__A1 _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3708__A2 _3707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3353__A _5216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _3127_/B _4729_/B _4413_/C _3158_/X _3159_/X vssd1 vssd1 vccd1 vccd1 _3160_/X
+ sky130_fd_sc_hd__a2111o_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3072__B _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3091_ _4051_/B _3125_/C vssd1 vssd1 vccd1 vccd1 _5362_/B sky130_fd_sc_hd__or2_2
XANTENNA_clkbuf_leaf_22_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__5094__B1 _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5801_ _5800_/X _3707_/X _5831_/S vssd1 vssd1 vccd1 vccd1 _5801_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_76_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xci2406_z80_187 vssd1 vssd1 vccd1 vccd1 ci2406_z80_187/HI io_oeb[2] sky130_fd_sc_hd__conb_1
XFILLER_0_91_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5732_ _3926_/X _5715_/B _5715_/Y _5731_/X vssd1 vssd1 vccd1 vccd1 _5732_/X sky130_fd_sc_hd__o22a_1
X_3993_ _4223_/A _5054_/A vssd1 vssd1 vccd1 vccd1 _3993_/Y sky130_fd_sc_hd__nor2_1
Xci2406_z80_198 vssd1 vssd1 vccd1 vccd1 ci2406_z80_198/HI io_oeb[13] sky130_fd_sc_hd__conb_1
XANTENNA__4912__A _6237_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5663_ _5615_/X _5661_/X _5662_/X vssd1 vssd1 vccd1 vccd1 _5664_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__5149__A1 _6238_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5594_ _6194_/Q _5606_/S _4866_/X vssd1 vssd1 vccd1 vccd1 _5594_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4614_ _5502_/B _4614_/B _4614_/C _4614_/D vssd1 vssd1 vccd1 vccd1 _4615_/D sky130_fd_sc_hd__or4_1
Xhold401 _5273_/X vssd1 vssd1 vccd1 vccd1 _6138_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4545_ _4545_/A _4545_/B vssd1 vssd1 vccd1 vccd1 _4547_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3247__B _5093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold412 _6181_/Q vssd1 vssd1 vccd1 vccd1 hold412/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 _6068_/Q vssd1 vssd1 vccd1 vccd1 hold423/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold434 _5788_/X vssd1 vssd1 vccd1 vccd1 _6234_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3580__B1 _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold445 _6169_/Q vssd1 vssd1 vccd1 vccd1 _3508_/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold467 _5672_/X vssd1 vssd1 vccd1 vccd1 _6200_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold478 _6229_/Q vssd1 vssd1 vccd1 vccd1 hold478/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold456 _6228_/Q vssd1 vssd1 vccd1 vccd1 hold456/X sky130_fd_sc_hd__dlygate4sd3_1
X_4476_ _5872_/A _4565_/S vssd1 vssd1 vccd1 vccd1 _4611_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold489 _5777_/X vssd1 vssd1 vccd1 vccd1 _6223_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6215_ _6218_/CLK _6215_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6215_/Q sky130_fd_sc_hd__dfstp_1
X_3427_ _4094_/B _4070_/B _3827_/B _3154_/B vssd1 vssd1 vccd1 vccd1 _3427_/X sky130_fd_sc_hd__a31o_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ hold42/X _3353_/X _3376_/A vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__a21o_1
X_6146_ _6146_/CLK _6146_/D vssd1 vssd1 vccd1 vccd1 _6146_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4793__S _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3289_ _3289_/A vssd1 vssd1 vccd1 vccd1 _3289_/Y sky130_fd_sc_hd__inv_2
X_6077_ _6129_/CLK _6077_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6077_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4832__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5028_ _5028_/A _5375_/B _5375_/A vssd1 vssd1 vccd1 vccd1 _5029_/C sky130_fd_sc_hd__or3b_1
XFILLER_0_95_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4060__A1 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4899__A0 _4895_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5863__A2 _5836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5076__A0 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3348__A _3513_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4878__S _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6059__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4330_ _3737_/X hold305/X _4336_/S vssd1 vssd1 vccd1 vccd1 _4330_/X sky130_fd_sc_hd__mux2_1
X_4261_ _4252_/Y _4253_/X _4260_/X _4242_/S vssd1 vssd1 vccd1 vccd1 _4261_/X sky130_fd_sc_hd__a22o_2
X_6000_ _6029_/CLK _6000_/D vssd1 vssd1 vccd1 vccd1 _6000_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3314__B1 _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3212_ _3713_/A _3543_/B _3422_/B _3540_/A _3554_/A vssd1 vssd1 vccd1 vccd1 _3212_/X
+ sky130_fd_sc_hd__o221a_1
X_4192_ hold248/X hold159/X hold286/X hold82/X _5182_/S _4255_/S vssd1 vssd1 vccd1
+ vccd1 _4192_/X sky130_fd_sc_hd__mux4_1
X_3143_ _4417_/B _3210_/C vssd1 vssd1 vccd1 vccd1 _3143_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_89_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3074_ _3654_/S _3116_/A vssd1 vssd1 vccd1 vccd1 _3074_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_89_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3976_ _4223_/A _5053_/C vssd1 vssd1 vccd1 vccd1 _3976_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_fanout147_A _3302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5715_ _5764_/B _5715_/B vssd1 vssd1 vccd1 vccd1 _5715_/Y sky130_fd_sc_hd__nand2_2
X_5646_ _5672_/S _5645_/X _5624_/X _5636_/A vssd1 vssd1 vccd1 vccd1 _5646_/X sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5473__A _6157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5577_ _4119_/B _5576_/X _4850_/Y vssd1 vssd1 vccd1 vccd1 _5577_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__3692__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4788__S _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 _5963_/Q vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 _5970_/Q vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold231 _4352_/X vssd1 vssd1 vccd1 vccd1 _6017_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 _6035_/Q vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
X_4528_ _4575_/A _4527_/B _4527_/C vssd1 vssd1 vccd1 vccd1 _4529_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_13_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold286 _6023_/Q vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold275 _5948_/Q vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 _6000_/Q vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
X_4459_ _4391_/B _3388_/B _3386_/X _4457_/X _3272_/A vssd1 vssd1 vccd1 vccd1 _4459_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3305__B1 _5838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold297 _4293_/X vssd1 vssd1 vccd1 vccd1 _5957_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_6129_ _6129_/CLK _6129_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6129_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3792__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5383__A _6135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3615__B _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4446__B _4446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3350__B _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3830_ _4522_/B _3829_/Y _6074_/Q vssd1 vssd1 vccd1 vccd1 _3830_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4024__B2 _6172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4024__A1 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3761_ _5333_/B _3761_/B vssd1 vssd1 vccd1 vccd1 _3764_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3783__A0 _4507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5500_ _5872_/A _5313_/S _5499_/X _3405_/B vssd1 vssd1 vccd1 vccd1 _5707_/S sky130_fd_sc_hd__a211oi_4
X_3692_ _6135_/Q _6137_/Q _5868_/S vssd1 vssd1 vccd1 vccd1 _5395_/B sky130_fd_sc_hd__mux2_1
X_5431_ _2989_/Y _5317_/A _5430_/Y vssd1 vssd1 vccd1 vccd1 _5433_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4401__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5362_ _5362_/A _5362_/B _5424_/B _5424_/C vssd1 vssd1 vccd1 vccd1 _5363_/C sky130_fd_sc_hd__or4_4
XFILLER_0_50_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3525__B _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4313_ _3789_/X hold128/X _4318_/S vssd1 vssd1 vccd1 vccd1 _4313_/X sky130_fd_sc_hd__mux2_1
X_5293_ _5245_/A _5046_/A _5245_/Y _5292_/X vssd1 vssd1 vccd1 vccd1 _5293_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4244_ _4234_/A _4233_/Y _4238_/A vssd1 vssd1 vccd1 vccd1 _4251_/A sky130_fd_sc_hd__a21o_1
X_4175_ _4219_/A _4143_/Y _4174_/X _4145_/B _4158_/Y vssd1 vssd1 vccd1 vccd1 _4176_/B
+ sky130_fd_sc_hd__a221o_1
X_3126_ _3148_/C _3426_/A _3511_/C _3101_/Y vssd1 vssd1 vccd1 vccd1 _3126_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3260__B _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5460__A0 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3057_ _4426_/A _3483_/A _3057_/C _4727_/A vssd1 vssd1 vccd1 vccd1 _3086_/A sky130_fd_sc_hd__or4_1
XFILLER_0_18_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3959_ _3959_/A vssd1 vssd1 vccd1 vccd1 _3959_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3774__A0 _6115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5629_ _5629_/A _5629_/B vssd1 vssd1 vccd1 vccd1 _5629_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6299__A _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5515__A1 _6188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4311__S _4318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5754__B2 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3296__A2 _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5442__B1 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5980_ _6151_/CLK _5980_/D vssd1 vssd1 vccd1 vccd1 _5980_/Q sky130_fd_sc_hd__dfxtp_1
X_4931_ _6198_/Q _6064_/Q _6038_/Q vssd1 vssd1 vccd1 vccd1 _4931_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3453__C1 _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4862_ _4119_/B _4861_/X _4850_/Y vssd1 vssd1 vccd1 vccd1 _4862_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_74_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3813_ _5024_/B _3807_/X _3811_/A _3639_/X vssd1 vssd1 vccd1 vccd1 _3813_/X sky130_fd_sc_hd__a22o_1
XANTENNA_15 _6121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5745__B2 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_26 _4787_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4793_ _4789_/B _4792_/X _4963_/A vssd1 vssd1 vccd1 vccd1 _4793_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5823__A2_N _5352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3744_ _5209_/A _3744_/B _3744_/C vssd1 vssd1 vccd1 vccd1 _3744_/X sky130_fd_sc_hd__or3_1
XFILLER_0_15_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3675_ _5893_/Q _3591_/A _3740_/S hold658/X _5179_/S vssd1 vssd1 vccd1 vccd1 _3677_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5414_ _5475_/S _5414_/B vssd1 vssd1 vccd1 vccd1 _5414_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3536__A _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4720__A2 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5345_ _2959_/Y _5343_/X _5340_/Y vssd1 vssd1 vccd1 vccd1 _5345_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5276_ _6208_/Q _5251_/Y _5252_/Y _6216_/Q _5275_/X vssd1 vssd1 vccd1 vccd1 _5276_/X
+ sky130_fd_sc_hd__a221o_1
X_4227_ hold137/X _4226_/X _4262_/S vssd1 vssd1 vccd1 vccd1 _4227_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4158_ _4250_/A _4159_/B vssd1 vssd1 vccd1 vccd1 _4158_/Y sky130_fd_sc_hd__nor2_1
X_3109_ _3249_/A _3210_/C vssd1 vssd1 vccd1 vccd1 _4433_/B sky130_fd_sc_hd__nor2_2
X_4089_ _3097_/Y _3543_/B _4088_/X _3556_/A _4058_/X vssd1 vssd1 vccd1 vccd1 _4089_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3444__C1 _4451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4306__S _4309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5736__B2 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5197__C1 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3446__A _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold593_A _6238_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3165__B _4486_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3880__S _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5600__S _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3450__A2 _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5727__B2 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5836__A _5836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput13 rst_n vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3356__A _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3460_ _3556_/A _3459_/X _4377_/B vssd1 vssd1 vccd1 vccd1 _3460_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__3790__S _4035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3505__A3 _3383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3391_ _4460_/A _3384_/X hold581/X vssd1 vssd1 vccd1 vccd1 _3391_/X sky130_fd_sc_hd__a21o_1
X_5130_ _6237_/Q _5108_/Y _5129_/Y _6213_/Q vssd1 vssd1 vccd1 vccd1 _5130_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5112__C1 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5061_ hold7/X _3755_/Y _5296_/S vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__mux2_1
X_4012_ _4012_/A _4012_/B vssd1 vssd1 vccd1 vccd1 _4014_/B sky130_fd_sc_hd__nor2_1
XANTENNA__4618__C _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4915__A _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5963_ _6010_/CLK _5963_/D vssd1 vssd1 vccd1 vccd1 _5963_/Q sky130_fd_sc_hd__dfxtp_1
X_4914_ _6197_/Q _6063_/Q _5216_/A vssd1 vssd1 vccd1 vccd1 _4914_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5894_ _6006_/CLK _5894_/D vssd1 vssd1 vccd1 vccd1 _5894_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5718__B2 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4845_ _6058_/Q _4844_/X _5606_/S vssd1 vssd1 vccd1 vccd1 _4845_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4776_ _5013_/S vssd1 vssd1 vccd1 vccd1 _4776_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3727_ _3616_/B _3724_/X _3726_/Y _3968_/A vssd1 vssd1 vccd1 vccd1 _3730_/C sky130_fd_sc_hd__a211o_1
XFILLER_0_43_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3658_ _3657_/A _3646_/X _3657_/Y _3645_/X vssd1 vssd1 vccd1 vccd1 _3658_/X sky130_fd_sc_hd__a211o_1
X_3589_ _3988_/A _3616_/B _3982_/S vssd1 vssd1 vccd1 vccd1 _4132_/A sky130_fd_sc_hd__or3_4
X_5328_ _6074_/Q _3496_/X _3646_/X vssd1 vssd1 vccd1 vccd1 _5330_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5259_ _5259_/A _5259_/B vssd1 vssd1 vccd1 vccd1 _5259_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold606_A _6178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_12_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__4735__A _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4620__A1 _4617_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2960_ _6178_/Q vssd1 vssd1 vccd1 vccd1 _2960_/Y sky130_fd_sc_hd__inv_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4630_ _4628_/Y _4630_/B vssd1 vssd1 vccd1 vccd1 _4632_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4561_ _4561_/A _4561_/B vssd1 vssd1 vccd1 vccd1 _4563_/A sky130_fd_sc_hd__nand2_1
Xhold616 _6176_/Q vssd1 vssd1 vccd1 vccd1 hold616/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold627 _6164_/Q vssd1 vssd1 vccd1 vccd1 _3383_/A sky130_fd_sc_hd__buf_2
XFILLER_0_4_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold605 _5232_/X vssd1 vssd1 vccd1 vccd1 _6127_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3517__C _3517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4492_ _4618_/B _3714_/X _3716_/X _3712_/Y _4497_/S vssd1 vssd1 vccd1 vccd1 _4575_/A
+ sky130_fd_sc_hd__a311o_4
X_3512_ _3554_/A _5424_/B _5424_/C vssd1 vssd1 vccd1 vccd1 _3513_/C sky130_fd_sc_hd__or3_2
XFILLER_0_100_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6231_ _6235_/CLK _6231_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6231_/Q sky130_fd_sc_hd__dfstp_1
Xhold649 _6172_/Q vssd1 vssd1 vccd1 vccd1 hold649/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4136__B1 _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3443_ _3196_/B _3442_/X _4054_/C vssd1 vssd1 vccd1 vccd1 _3443_/X sky130_fd_sc_hd__o21a_1
Xhold638 _6254_/Q vssd1 vssd1 vccd1 vccd1 hold638/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ _6171_/CLK _6162_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6162_/Q sky130_fd_sc_hd__dfstp_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5113_ _6028_/Q _5200_/A2 _5200_/B1 _5920_/Q _4256_/S vssd1 vssd1 vccd1 vccd1 _5116_/C
+ sky130_fd_sc_hd__a221o_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ hold50/X _3366_/X _3376_/C _3373_/X _3364_/Y vssd1 vssd1 vccd1 vccd1 hold51/A
+ sky130_fd_sc_hd__a2111o_1
X_6093_ _6227_/CLK _6093_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6093_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ _5044_/A _5044_/B _5044_/C _3646_/X vssd1 vssd1 vccd1 vccd1 _5044_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_79_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout177_A fanout184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5946_ _6034_/CLK _5946_/D vssd1 vssd1 vccd1 vccd1 _5946_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5877_ hold353/X _5875_/X _5876_/Y _5873_/X vssd1 vssd1 vccd1 vccd1 _5877_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4828_ _6157_/Q _5008_/B _4826_/X _4999_/A1 vssd1 vssd1 vccd1 vccd1 _4829_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_47_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5167__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4759_ _4759_/A _4759_/B _4759_/C vssd1 vssd1 vccd1 vccd1 _4760_/D sky130_fd_sc_hd__and3_1
XFILLER_0_31_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4127__B1 _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4678__B2 _4474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6034_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_hold556_A _6165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3653__A2 _6172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5158__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4905__A2 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5315__C1 _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
X_3090_ _4051_/B _3125_/C vssd1 vssd1 vccd1 vccd1 _3090_/Y sky130_fd_sc_hd__nor2_1
X_5800_ hold412/X _5794_/Y _5799_/X _5794_/B vssd1 vssd1 vccd1 vccd1 _5800_/X sky130_fd_sc_hd__a22o_1
X_3992_ _4134_/B _3992_/B vssd1 vssd1 vccd1 vccd1 _5054_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xci2406_z80_188 vssd1 vssd1 vccd1 vccd1 ci2406_z80_188/HI io_oeb[3] sky130_fd_sc_hd__conb_1
XFILLER_0_29_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5731_ _4119_/A _4850_/B _4563_/Y _5762_/C vssd1 vssd1 vccd1 vccd1 _5731_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_9_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_199 vssd1 vssd1 vccd1 vccd1 ci2406_z80_199/HI io_oeb[14] sky130_fd_sc_hd__conb_1
XFILLER_0_84_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4912__B _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5662_ _6196_/Q _6197_/Q _6198_/Q _6199_/Q _5685_/B vssd1 vssd1 vccd1 vccd1 _5662_/X
+ sky130_fd_sc_hd__o41a_1
X_5593_ _5604_/B _5593_/B vssd1 vssd1 vccd1 vccd1 _5593_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4613_ _4613_/A _4613_/B _4613_/C vssd1 vssd1 vccd1 vccd1 _4760_/B sky130_fd_sc_hd__nor3_1
X_4544_ _4575_/A _4543_/B _4543_/C vssd1 vssd1 vccd1 vccd1 _4545_/B sky130_fd_sc_hd__a21o_1
Xhold402 _6171_/Q vssd1 vssd1 vccd1 vccd1 _5498_/A sky130_fd_sc_hd__buf_1
XFILLER_0_13_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold413 _5491_/X vssd1 vssd1 vccd1 vccd1 _6181_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold424 _4710_/X vssd1 vssd1 vccd1 vccd1 _6068_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 _6115_/Q vssd1 vssd1 vccd1 vccd1 _2977_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xhold468 _6227_/Q vssd1 vssd1 vccd1 vccd1 hold468/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6214_ _6218_/CLK _6214_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6214_/Q sky130_fd_sc_hd__dfstp_1
Xhold457 _5782_/X vssd1 vssd1 vccd1 vccd1 _6228_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5857__A0 _6117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4475_ _6129_/Q _4497_/S vssd1 vssd1 vccd1 vccd1 _4565_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_13_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold446 _3515_/X vssd1 vssd1 vccd1 vccd1 _3516_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold479 _5783_/X vssd1 vssd1 vccd1 vccd1 _6229_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3426_ _3426_/A _5356_/A _3694_/C vssd1 vssd1 vccd1 vccd1 _3827_/B sky130_fd_sc_hd__and3_1
XFILLER_0_96_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _3370_/B _3356_/X _3353_/X vssd1 vssd1 vccd1 vccd1 _3376_/A sky130_fd_sc_hd__a21oi_1
X_6145_ _6151_/CLK hold85/X vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_99_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3883__A2 _3588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ _6129_/CLK hold35/X fanout170/X vssd1 vssd1 vccd1 vccd1 _6076_/Q sky130_fd_sc_hd__dfrtp_1
X_3288_ _3446_/A _3288_/B vssd1 vssd1 vccd1 vccd1 _3289_/A sky130_fd_sc_hd__and2_1
X_5027_ _2960_/Y _6045_/Q _5374_/A _5374_/B vssd1 vssd1 vccd1 vccd1 _5028_/A sky130_fd_sc_hd__a211o_1
XANTENNA__4094__B _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5929_ _6034_/CLK hold79/X vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_0_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4314__S _4318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5356__D _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3571__A1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5848__A0 _6119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3454__A _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4520__A0 _6156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3629__A _6135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4451__C _4451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3348__B _3383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3364__A _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4260_ _5116_/A _4256_/X _4259_/X vssd1 vssd1 vccd1 vccd1 _4260_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4191_ hold9/X _4253_/A2 _3833_/Y _4190_/Y vssd1 vssd1 vccd1 vccd1 _4191_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3314__B2 _3488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4894__S _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3211_ _3554_/A _3439_/B _3306_/C _3422_/B vssd1 vssd1 vccd1 vccd1 _3211_/Y sky130_fd_sc_hd__nand4_2
X_3142_ _3148_/B _5356_/A _3141_/X _3112_/A vssd1 vssd1 vccd1 vccd1 _3142_/Y sky130_fd_sc_hd__o211ai_1
X_3073_ _4486_/A _3208_/A vssd1 vssd1 vccd1 vccd1 _4117_/C sky130_fd_sc_hd__nor2_2
XFILLER_0_89_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3975_ _3975_/A _3975_/B vssd1 vssd1 vccd1 vccd1 _5053_/C sky130_fd_sc_hd__or2_1
X_5714_ _5715_/B _5713_/A _5767_/A vssd1 vssd1 vccd1 vccd1 _5714_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5645_ _4940_/Y _5629_/Y _5644_/X _5640_/X _5511_/X vssd1 vssd1 vccd1 vccd1 _5645_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5473__B _6156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold210 _4166_/X vssd1 vssd1 vccd1 vccd1 _5921_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_60_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5576_ _5575_/X _6059_/Q _5595_/S vssd1 vssd1 vccd1 vccd1 _5576_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3553__A1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3002__B1 _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold243 _4372_/X vssd1 vssd1 vccd1 vccd1 _6035_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 _5897_/Q vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
X_4527_ _4575_/A _4527_/B _4527_/C vssd1 vssd1 vccd1 vccd1 _4529_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_13_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3274__A _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold221 _4299_/X vssd1 vssd1 vccd1 vccd1 _5963_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _4287_/X vssd1 vssd1 vccd1 vccd1 _5948_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold265 _5949_/Q vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold254 _5971_/Q vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4458_ _3694_/C _3388_/B _3386_/X _4457_/X _3272_/B vssd1 vssd1 vccd1 vccd1 _4458_/X
+ sky130_fd_sc_hd__a32o_1
Xhold287 _6133_/Q vssd1 vssd1 vccd1 vccd1 _3517_/A sky130_fd_sc_hd__buf_1
X_3409_ _6048_/Q _3395_/B _3488_/B _3408_/X _4728_/B vssd1 vssd1 vccd1 vccd1 _3409_/X
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__3305__A1 _4433_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold298 _6123_/Q vssd1 vssd1 vccd1 vccd1 _3523_/A sky130_fd_sc_hd__dlygate4sd3_1
X_6128_ _6130_/CLK _6128_/D fanout171/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__dfrtp_2
X_4389_ _4398_/A _5360_/D _3337_/D _4445_/B vssd1 vssd1 vccd1 vccd1 _4389_/X sky130_fd_sc_hd__o211a_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5058__A1 _5249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4309__S _4309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6059_ _6060_/CLK _6059_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6059_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5230__A1 _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4979__S _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6192__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5049__B2 _2960_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4257__C1 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3350__C _3503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4655__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3760_ _5024_/A _6115_/Q vssd1 vssd1 vccd1 vccd1 _3764_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3359__A _5220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4980__A0 _4976_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5430_ _6175_/Q _5352_/A _5354_/Y vssd1 vssd1 vccd1 vccd1 _5430_/Y sky130_fd_sc_hd__a21oi_1
X_3691_ _6114_/Q _6118_/Q _6070_/Q vssd1 vssd1 vccd1 vccd1 _5404_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5361_ _5363_/B vssd1 vssd1 vccd1 vccd1 _5475_/S sky130_fd_sc_hd__inv_2
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3094__A _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5292_ _5248_/Y _5289_/X _5291_/X vssd1 vssd1 vccd1 vccd1 _5292_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4312_ _3737_/X hold149/X _4318_/S vssd1 vssd1 vccd1 vccd1 _4312_/X sky130_fd_sc_hd__mux2_1
X_4243_ hold157/X _4242_/X _4262_/S vssd1 vssd1 vccd1 vccd1 _4243_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5288__A1 _5245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4174_ _4146_/B _4174_/B vssd1 vssd1 vccd1 vccd1 _4174_/X sky130_fd_sc_hd__and2b_1
X_3125_ _3426_/A _4739_/A _3125_/C _4056_/B vssd1 vssd1 vccd1 vccd1 _3125_/X sky130_fd_sc_hd__or4_1
XFILLER_0_96_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3056_ _3396_/A _3056_/B vssd1 vssd1 vccd1 vccd1 _4727_/A sky130_fd_sc_hd__or2_1
XFILLER_0_77_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5212__A1 _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3958_ _3957_/X _2980_/Y _3958_/S vssd1 vssd1 vccd1 vccd1 _3959_/A sky130_fd_sc_hd__mux2_4
XANTENNA__3774__A1 _6119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3889_ _4234_/A _3890_/B vssd1 vssd1 vccd1 vccd1 _3974_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5628_ _5661_/A _5628_/B vssd1 vssd1 vccd1 vccd1 _5628_/Y sky130_fd_sc_hd__xnor2_1
X_5559_ _5559_/A _5571_/B vssd1 vssd1 vccd1 vccd1 _5559_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout72_A _3582_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold636_A _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3462__B1 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3626__B _6113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4930_ _6214_/Q _5009_/A2 _4769_/Y _4928_/B _4929_/X vssd1 vssd1 vccd1 vccd1 _4930_/X
+ sky130_fd_sc_hd__a221o_1
X_4861_ _4860_/X _6059_/Q _5595_/S vssd1 vssd1 vccd1 vccd1 _4861_/X sky130_fd_sc_hd__mux2_1
X_3812_ _3811_/A _3811_/B _3647_/C vssd1 vssd1 vccd1 vccd1 _3812_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_16 _6121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 _4819_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4792_ _6189_/Q _6055_/Q _6038_/Q vssd1 vssd1 vccd1 vccd1 _4792_/X sky130_fd_sc_hd__mux2_1
X_3743_ _5998_/Q _3591_/A _3739_/S _5959_/Q _4256_/S vssd1 vssd1 vccd1 vccd1 _3744_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3674_ _3672_/X _3673_/X _4256_/S vssd1 vssd1 vccd1 vccd1 _3674_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5413_ _5365_/S _5369_/X _5382_/X _5412_/Y vssd1 vssd1 vccd1 vccd1 _5414_/B sky130_fd_sc_hd__o22a_1
XANTENNA__3536__B _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5344_ _5507_/A _3193_/C _4614_/B _5343_/X _2959_/Y vssd1 vssd1 vccd1 vccd1 _5344_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__6043__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5275_ _6158_/Q _5253_/Y _5254_/Y _6240_/Q vssd1 vssd1 vccd1 vccd1 _5275_/X sky130_fd_sc_hd__a22o_1
X_4226_ _4224_/X _4225_/X _4242_/S vssd1 vssd1 vccd1 vccd1 _4226_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4157_ _4159_/B vssd1 vssd1 vccd1 vccd1 _4157_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3692__A0 _6135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3108_ _4061_/A _3208_/B vssd1 vssd1 vccd1 vccd1 _3306_/A sky130_fd_sc_hd__or2_1
X_4088_ _4124_/B _3143_/Y _4087_/X _3694_/C vssd1 vssd1 vccd1 vccd1 _4088_/X sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_37_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6175_/CLK
+ sky130_fd_sc_hd__clkbuf_16
X_3039_ _3777_/A _5356_/A vssd1 vssd1 vccd1 vccd1 _5489_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_65_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5197__B1 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4322__S _4327_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3446__B _4043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3199__C1 _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3356__B _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3390_ _3208_/A _3388_/B _3386_/X _3389_/X vssd1 vssd1 vccd1 vccd1 _3390_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5063__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5112__B1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5060_ hold11/X _3729_/Y _5296_/S vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__mux2_1
X_4011_ _4011_/A _4011_/B vssd1 vssd1 vccd1 vccd1 _4013_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4871__C1 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4915__B _4915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5962_ _6029_/CLK _5962_/D vssd1 vssd1 vccd1 vccd1 _5962_/Q sky130_fd_sc_hd__dfxtp_1
X_4913_ _6213_/Q _5009_/A2 _4769_/Y _4915_/B _4912_/X vssd1 vssd1 vccd1 vccd1 _4913_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5893_ _6146_/CLK _5893_/D vssd1 vssd1 vccd1 vccd1 _5893_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4844_ _6192_/Q _4767_/X _4842_/X _4843_/X vssd1 vssd1 vccd1 vccd1 _4844_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_7_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4775_ _3399_/B _4774_/Y _5838_/C vssd1 vssd1 vccd1 vccd1 _5013_/S sky130_fd_sc_hd__o21a_4
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3726_ _2972_/Y _3724_/S _3725_/X _3616_/B vssd1 vssd1 vccd1 vccd1 _3726_/Y sky130_fd_sc_hd__a211oi_1
XFILLER_0_43_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5762__A _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3657_ _3657_/A _3950_/B vssd1 vssd1 vccd1 vccd1 _3657_/Y sky130_fd_sc_hd__nor2_1
X_3588_ _3968_/A _3983_/S _3724_/S vssd1 vssd1 vccd1 vccd1 _3588_/X sky130_fd_sc_hd__and3_4
X_5327_ _5790_/D _5327_/B _5790_/B _5790_/C vssd1 vssd1 vccd1 vccd1 _5487_/S sky130_fd_sc_hd__nand4b_4
XANTENNA__4809__C _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5258_ _5245_/A hold508/X _5245_/Y _5257_/X vssd1 vssd1 vccd1 vccd1 _5258_/X sky130_fd_sc_hd__a22o_1
X_4209_ hold29/X _4253_/A2 _3865_/Y _4208_/Y vssd1 vssd1 vccd1 vccd1 _4209_/X sky130_fd_sc_hd__o22a_1
X_5189_ _6193_/Q _5122_/Y _5186_/X _5109_/Y vssd1 vssd1 vccd1 vccd1 _5189_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4209__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4317__S _4318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire93 wire93/A vssd1 vssd1 vccd1 vccd1 wire93/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4393__A1 _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3457__A _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout180 fanout183/X vssd1 vssd1 vccd1 vccd1 fanout180/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__6207__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5611__S _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4735__B _4759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3408__B1 _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4081__B1 _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _4575_/A _4559_/B _4559_/C vssd1 vssd1 vccd1 vccd1 _4561_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_25_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold617 _5453_/X vssd1 vssd1 vccd1 vccd1 _6176_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold606 _6178_/Q vssd1 vssd1 vccd1 vccd1 hold606/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4491_ _5296_/S _4482_/X _4490_/X hold527/X vssd1 vssd1 vccd1 vccd1 _4491_/X sky130_fd_sc_hd__a22o_1
X_3511_ _4118_/A _4497_/S _3511_/C _3511_/D vssd1 vssd1 vccd1 vccd1 _3511_/X sky130_fd_sc_hd__and4_1
XFILLER_0_100_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6230_ _6247_/CLK _6230_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6230_/Q sky130_fd_sc_hd__dfstp_1
Xhold628 _6074_/Q vssd1 vssd1 vccd1 vccd1 hold628/X sky130_fd_sc_hd__dlygate4sd3_1
X_3442_ _4398_/A _5502_/D _3396_/A vssd1 vssd1 vccd1 vccd1 _3442_/X sky130_fd_sc_hd__a21o_1
Xhold639 _5881_/X vssd1 vssd1 vccd1 vccd1 _6254_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6161_ _6242_/CLK _6161_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6161_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ hold44/X _5977_/Q hold33/X _5979_/Q _3353_/X vssd1 vssd1 vccd1 vccd1 _3373_/X
+ sky130_fd_sc_hd__o41a_1
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5945_/Q _5200_/A2 _5200_/B1 _6012_/Q _5182_/S vssd1 vssd1 vccd1 vccd1 _5116_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6092_ _6227_/CLK _6092_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6092_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _6117_/Q _3238_/Y _3778_/B _6115_/Q _5042_/X vssd1 vssd1 vccd1 vccd1 _5044_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5521__S _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5945_ _6110_/CLK _5945_/D vssd1 vssd1 vccd1 vccd1 _5945_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4072__B1 _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5876_ _5341_/A _4479_/C _5875_/X vssd1 vssd1 vccd1 vccd1 _5876_/Y sky130_fd_sc_hd__o21ai_4
X_4827_ _6207_/Q _4768_/Y _4769_/Y _4821_/B _4815_/B vssd1 vssd1 vccd1 vccd1 _4829_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3277__A _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4758_ _4735_/A _4614_/B _4728_/C _5502_/A vssd1 vssd1 vccd1 vccd1 _4760_/C sky130_fd_sc_hd__a211oi_1
X_4689_ _4687_/Y _4703_/B vssd1 vssd1 vccd1 vccd1 _4691_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3709_ _4737_/A _3709_/B vssd1 vssd1 vccd1 vccd1 _3709_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4678__A2 _4612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5627__A1 _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4836__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5563__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5606__S _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4510__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5866__A1 _3959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3650__A _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3991_ _4234_/A _3970_/B _3975_/A vssd1 vssd1 vccd1 vccd1 _3992_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5730_ hold563/X _5714_/Y _5729_/X _5023_/A vssd1 vssd1 vccd1 vccd1 _5730_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xci2406_z80_189 vssd1 vssd1 vccd1 vccd1 ci2406_z80_189/HI io_oeb[4] sky130_fd_sc_hd__conb_1
XFILLER_0_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5661_ _5661_/A _5661_/B vssd1 vssd1 vccd1 vccd1 _5661_/X sky130_fd_sc_hd__and2_1
X_4612_ _5762_/A _4612_/B vssd1 vssd1 vccd1 vccd1 _4612_/X sky130_fd_sc_hd__or2_1
X_5592_ _5592_/A _5592_/B _5590_/Y vssd1 vssd1 vccd1 vccd1 _5593_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4543_ _4575_/A _4543_/B _4543_/C vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3565__C1 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5306__A0 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold436 _5151_/X vssd1 vssd1 vccd1 vccd1 _6115_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold414 _6194_/Q vssd1 vssd1 vccd1 vccd1 _2996_/A sky130_fd_sc_hd__buf_1
XFILLER_0_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold425 _6191_/Q vssd1 vssd1 vccd1 vccd1 _2993_/A sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold403 _3522_/X vssd1 vssd1 vccd1 vccd1 _6171_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3580__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold469 _5781_/X vssd1 vssd1 vccd1 vccd1 _6227_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 _6069_/Q vssd1 vssd1 vccd1 vccd1 hold458/X sky130_fd_sc_hd__dlygate4sd3_1
X_6213_ _6218_/CLK _6213_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6213_/Q sky130_fd_sc_hd__dfstp_1
X_4474_ _4474_/A _4497_/S vssd1 vssd1 vccd1 vccd1 _4474_/X sky130_fd_sc_hd__and2_4
Xhold447 _3516_/X vssd1 vssd1 vccd1 vccd1 _6169_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3425_ _5875_/A _3423_/X hold378/X vssd1 vssd1 vccd1 vccd1 _3425_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _4077_/A _4124_/A _4765_/A _3363_/B vssd1 vssd1 vccd1 vccd1 _3356_/X sky130_fd_sc_hd__or4_1
X_6144_ _6144_/CLK hold24/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfxtp_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _4043_/C _5498_/B vssd1 vssd1 vccd1 vccd1 _3288_/B sky130_fd_sc_hd__nand2_1
X_6075_ _6129_/CLK hold51/X fanout170/X vssd1 vssd1 vccd1 vccd1 _6075_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5026_ _5026_/A vssd1 vssd1 vccd1 vccd1 _5026_/Y sky130_fd_sc_hd__inv_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4596__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5928_ _6149_/CLK _5928_/D vssd1 vssd1 vccd1 vccd1 _5928_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4391__A _6127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5859_ hold334/X _5836_/A _5858_/X _5245_/A vssd1 vssd1 vccd1 vccd1 _5859_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_63_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5545__B1 _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4330__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5848__A1 _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3454__B _5424_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5784__A0 _6174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4505__S _4598_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4451__D _5917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5000__A2 _4766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4190_ _4223_/A _5055_/B vssd1 vssd1 vccd1 vccd1 _4190_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3210_ _3210_/A _4485_/A _3210_/C vssd1 vssd1 vccd1 vccd1 _3422_/B sky130_fd_sc_hd__or3_2
XANTENNA__4476__A _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3141_ _3148_/B _3777_/A _3643_/A _4485_/A vssd1 vssd1 vccd1 vccd1 _3141_/X sky130_fd_sc_hd__a31o_1
XANTENNA__5071__S _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3072_ _3556_/A _4061_/A vssd1 vssd1 vccd1 vccd1 _3208_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_89_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4027__A0 _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5775__A0 _6237_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3974_ _3974_/A _3974_/B _3974_/C vssd1 vssd1 vccd1 vccd1 _3975_/B sky130_fd_sc_hd__and3_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5713_ _5713_/A vssd1 vssd1 vccd1 vccd1 _5713_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_72_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3539__B _3539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5644_ _4928_/Y _5643_/Y _5704_/S vssd1 vssd1 vccd1 vccd1 _5644_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold211 _5927_/Q vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold200 _4342_/X vssd1 vssd1 vccd1 vccd1 _6008_/D sky130_fd_sc_hd__dlygate4sd3_1
X_5575_ _6193_/Q _5606_/S _4851_/X vssd1 vssd1 vccd1 vccd1 _5575_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_53_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5473__C _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4526_ _6207_/Q _4821_/B _4589_/S vssd1 vssd1 vccd1 vccd1 _4527_/C sky130_fd_sc_hd__mux2_1
Xhold222 _5895_/Q vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 _5977_/Q vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 _6122_/Q vssd1 vssd1 vccd1 vccd1 _3532_/B sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3274__B _4104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold266 _6016_/Q vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _6030_/Q vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 _6013_/Q vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
X_4457_ _4457_/A _4457_/B vssd1 vssd1 vccd1 vccd1 _4457_/X sky130_fd_sc_hd__or2_1
XANTENNA__4502__B2 _4474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3408_ _4483_/A _4439_/B _4036_/B vssd1 vssd1 vccd1 vccd1 _3408_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold299 _3524_/X vssd1 vssd1 vccd1 vccd1 _6122_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 _4454_/X vssd1 vssd1 vccd1 vccd1 _6048_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6127_ _6130_/CLK _6127_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6127_/Q sky130_fd_sc_hd__dfrtp_4
X_4388_ _4048_/A _4384_/X _4386_/X _4387_/X _4485_/B vssd1 vssd1 vccd1 vccd1 _4388_/Y
+ sky130_fd_sc_hd__o311ai_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _5918_/Q _3320_/B _3335_/X _3338_/Y _6130_/Q vssd1 vssd1 vccd1 vccd1 _3344_/S
+ sky130_fd_sc_hd__a2111o_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ _6060_/CLK _6058_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6058_/Q sky130_fd_sc_hd__dfrtp_4
X_5009_ _6219_/Q _5009_/A2 _4769_/Y _5007_/B _5008_/X vssd1 vssd1 vccd1 vccd1 _5009_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4325__S _4327_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5766__B1 _5771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3792__A2 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3544__A2 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4655__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3359__B _3370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5509__B1 _5220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3690_ _5024_/A _6136_/Q _6114_/Q _3848_/B _3689_/X vssd1 vssd1 vccd1 vccd1 _5374_/B
+ sky130_fd_sc_hd__o41a_2
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5360_ _5360_/A _5424_/B _5566_/S _5360_/D vssd1 vssd1 vccd1 vccd1 _5363_/B sky130_fd_sc_hd__or4_4
XFILLER_0_77_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5291_ hold583/X _5251_/Y _5252_/Y hold554/X _5290_/X vssd1 vssd1 vccd1 vccd1 _5291_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4311_ _3668_/X hold217/X _4318_/S vssd1 vssd1 vccd1 vccd1 _4311_/X sky130_fd_sc_hd__mux2_1
X_4242_ _4240_/X _4241_/X _4242_/S vssd1 vssd1 vccd1 vccd1 _4242_/X sky130_fd_sc_hd__mux2_2
X_4173_ _4250_/A _4173_/B vssd1 vssd1 vccd1 vccd1 _4195_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4248__B1 _3615_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3124_ _3182_/A _3507_/D _3120_/B vssd1 vssd1 vccd1 vccd1 _3124_/Y sky130_fd_sc_hd__a21oi_1
X_3055_ _4051_/B _3182_/B _3182_/A vssd1 vssd1 vccd1 vccd1 _3056_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__4799__A1 _6189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout152_A _6112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3957_ _4570_/B _3956_/Y _6074_/Q vssd1 vssd1 vccd1 vccd1 _3957_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3223__A1 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4420__B1 _5838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3888_ _3888_/A _3888_/B _3887_/Y vssd1 vssd1 vccd1 vccd1 _3890_/B sky130_fd_sc_hd__or3b_4
X_5627_ _6196_/Q _5685_/B _5615_/X vssd1 vssd1 vccd1 vccd1 _5628_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4723__A1 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5558_ _5557_/X _2993_/A _5705_/S vssd1 vssd1 vccd1 vccd1 _5558_/X sky130_fd_sc_hd__mux2_1
X_4509_ _5982_/Q hold88/A _5998_/Q _5959_/Q _5076_/A0 _4272_/B vssd1 vssd1 vccd1 vccd1
+ _4509_/X sky130_fd_sc_hd__mux4_1
X_5489_ _6165_/Q _5489_/B _5489_/C _5489_/D vssd1 vssd1 vccd1 vccd1 _5497_/S sky130_fd_sc_hd__nand4_4
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold531_A _6188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold629_A _6158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3462__A1 _4478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3366__A_N _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_31_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_7_wb_clk_i _5978_/CLK vssd1 vssd1 vccd1 vccd1 _6192_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_47_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4650__B1 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3453__A1 _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4860_ _5606_/S _4859_/X _4851_/X vssd1 vssd1 vccd1 vccd1 _4860_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_47_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3811_ _3811_/A _3811_/B vssd1 vssd1 vccd1 vccd1 _3811_/X sky130_fd_sc_hd__or2_1
XANTENNA__4402__B1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_28 _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_17 _6121_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4791_ _4789_/B _4769_/Y _5008_/B _6155_/Q vssd1 vssd1 vccd1 vccd1 _4791_/X sky130_fd_sc_hd__a22o_1
XANTENNA__4953__A1 _6199_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3742_ _5894_/Q _3591_/A _3739_/S _6006_/Q _5179_/S vssd1 vssd1 vccd1 vccd1 _3744_/B
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3673_ hold90/A _5981_/Q _3740_/S vssd1 vssd1 vccd1 vccd1 _3673_/X sky130_fd_sc_hd__mux2_1
X_5412_ _5392_/Y _5393_/X _5411_/Y vssd1 vssd1 vccd1 vccd1 _5412_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__3536__C _4726_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5343_ _3249_/B _4061_/C _3116_/A _4760_/C _5338_/Y vssd1 vssd1 vccd1 vccd1 _5343_/X
+ sky130_fd_sc_hd__o311a_2
XANTENNA__4929__A _6238_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5274_ _3875_/B _4203_/Y _5289_/S vssd1 vssd1 vccd1 vccd1 _5274_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4225_ hold253/X hold175/X hold228/X hold72/X _5182_/S _5200_/B1 vssd1 vssd1 vccd1
+ vccd1 _4225_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5130__A1 _6237_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4156_ _4156_/A _4156_/B vssd1 vssd1 vccd1 vccd1 _4159_/B sky130_fd_sc_hd__nor2_2
XANTENNA__3692__A1 _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3107_ _3643_/A _3208_/B vssd1 vssd1 vccd1 vccd1 _5489_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3979__S _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4087_ _3221_/X _3439_/Y _3469_/Y vssd1 vssd1 vccd1 vccd1 _4087_/X sky130_fd_sc_hd__a21o_1
X_3038_ _4051_/B _3323_/C vssd1 vssd1 vccd1 vccd1 _3411_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_77_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4989_ hold339/X _4988_/X _5020_/S vssd1 vssd1 vccd1 vccd1 _4989_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_46_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4555__S0 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3435__A1 _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5188__A1 _6241_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5609__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4935__A1 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4935__B2 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3356__C _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4010_ _6141_/Q _4009_/C _5046_/A vssd1 vssd1 vccd1 vccd1 _4011_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__4871__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5961_ _6029_/CLK _5961_/D vssd1 vssd1 vccd1 vccd1 _5961_/Q sky130_fd_sc_hd__dfxtp_1
X_4912_ _6237_/Q _5008_/B vssd1 vssd1 vccd1 vccd1 _4912_/X sky130_fd_sc_hd__and2_1
XANTENNA__3977__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5892_ _6151_/CLK _5892_/D vssd1 vssd1 vccd1 vccd1 _5892_/Q sky130_fd_sc_hd__dfxtp_1
X_4843_ _6158_/Q _5008_/B _4838_/X _4999_/A1 _4841_/Y vssd1 vssd1 vccd1 vccd1 _4843_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5519__S _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4926__A1 _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4423__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4774_ _5338_/D _4774_/B vssd1 vssd1 vccd1 vccd1 _4774_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3725_ _3573_/C _3986_/A2 _3584_/X _3585_/X _2971_/Y vssd1 vssd1 vccd1 vccd1 _3725_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_15_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3656_ _3950_/B vssd1 vssd1 vccd1 vccd1 _3656_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4154__A2 _3588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3587_ _3573_/C _3986_/A2 _3584_/X _3585_/X vssd1 vssd1 vccd1 vccd1 _3885_/S sky130_fd_sc_hd__o31a_4
X_5326_ _5790_/D _5327_/B _5790_/B _5790_/C vssd1 vssd1 vccd1 vccd1 _5326_/X sky130_fd_sc_hd__and4b_2
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5257_ _5246_/Y _5248_/Y _5249_/Y _5256_/X vssd1 vssd1 vccd1 vccd1 _5257_/X sky130_fd_sc_hd__a31o_1
X_4208_ _4223_/A _5055_/C vssd1 vssd1 vccd1 vccd1 _4208_/Y sky130_fd_sc_hd__nor2_1
X_5188_ _6241_/Q _5108_/Y _5119_/Y _6201_/Q vssd1 vssd1 vccd1 vccd1 _5188_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3665__A1 _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4139_ hold151/X _4355_/A _4319_/B hold145/X _4138_/X vssd1 vssd1 vccd1 vccd1 _4142_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4090__B2 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4333__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3457__B _5424_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3192__B _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout181 fanout183/X vssd1 vssd1 vccd1 vccd1 fanout181/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__4853__A0 _4850_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout170 fanout171/X vssd1 vssd1 vccd1 vccd1 fanout170/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_88_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4908__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3510_ _3517_/A _3508_/X _3509_/Y vssd1 vssd1 vccd1 vccd1 _3510_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_25_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4490_ _5341_/A _4598_/S _4612_/B _5023_/A vssd1 vssd1 vccd1 vccd1 _4490_/X sky130_fd_sc_hd__a31o_1
Xhold607 _6049_/Q vssd1 vssd1 vccd1 vccd1 hold607/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold618 _6072_/Q vssd1 vssd1 vccd1 vccd1 hold618/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold629 _6158_/Q vssd1 vssd1 vccd1 vccd1 hold629/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5074__S _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3344__A0 _3539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3441_ _5838_/B _5838_/C _3437_/Y _3440_/X vssd1 vssd1 vccd1 vccd1 _3441_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4479__A _5875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6160_ _6238_/CLK _6160_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6160_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3372_/A _3372_/B vssd1 vssd1 vccd1 vccd1 _3376_/C sky130_fd_sc_hd__or2_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5111_ _6004_/Q _3591_/A _3740_/S _5892_/Q _4256_/S vssd1 vssd1 vccd1 vccd1 _5114_/C
+ sky130_fd_sc_hd__a221o_1
X_6091_ _6227_/CLK _6091_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6091_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5097__B1 _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _6119_/Q _4036_/B _3921_/A _6118_/Q vssd1 vssd1 vccd1 vccd1 _5042_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3111__A3 _4433_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5103__A _5120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5944_ _6111_/CLK _5944_/D vssd1 vssd1 vccd1 vccd1 _5944_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4072__A1 _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5875_ _5875_/A _5875_/B _5875_/C vssd1 vssd1 vccd1 vccd1 _5875_/X sky130_fd_sc_hd__and3_4
XFILLER_0_90_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4826_ _4821_/B _4825_/X _4963_/A vssd1 vssd1 vccd1 vccd1 _4826_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_62_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5773__A _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4757_ _4990_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _4757_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4688_ _4699_/A _4688_/B vssd1 vssd1 vccd1 vccd1 _4703_/B sky130_fd_sc_hd__nand2_1
X_3708_ _4223_/A _3707_/X _3573_/B vssd1 vssd1 vccd1 vccd1 _3708_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_31_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4780__C1 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5324__B2 _3539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3639_ _6072_/Q _6070_/Q _5024_/A vssd1 vssd1 vccd1 vccd1 _3639_/X sky130_fd_sc_hd__and3_2
XFILLER_0_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3335__B1 _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5309_ input4/X hold623/X _5313_/S vssd1 vssd1 vccd1 vccd1 _5309_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3886__A1 _3582_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5627__A2 _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4836__B _4836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6218_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4063__A1 _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold611_A _6170_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4998__S _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5622__S _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5618__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3990_ _4250_/A _3990_/B vssd1 vssd1 vccd1 vccd1 _4134_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4762__A _6048_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5660_ _5660_/A _5660_/B vssd1 vssd1 vccd1 vccd1 _5661_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5069__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4611_ _4611_/A _4631_/B _4611_/C vssd1 vssd1 vccd1 vccd1 _4611_/X sky130_fd_sc_hd__and3_1
XFILLER_0_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5591_ _5592_/A _5592_/B _5590_/Y vssd1 vssd1 vccd1 vccd1 _5604_/B sky130_fd_sc_hd__o21ba_1
X_4542_ _6208_/Q _4836_/B _4589_/S vssd1 vssd1 vccd1 vccd1 _4543_/C sky130_fd_sc_hd__mux2_1
Xhold404 _6175_/Q vssd1 vssd1 vccd1 vccd1 hold404/X sky130_fd_sc_hd__dlymetal6s2s_1
Xhold415 _5600_/X vssd1 vssd1 vccd1 vccd1 _6194_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4473_ _4589_/S _4472_/Y _4501_/A vssd1 vssd1 vccd1 vccd1 _4473_/Y sky130_fd_sc_hd__a21oi_1
Xhold426 _5561_/X vssd1 vssd1 vccd1 vccd1 _6191_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold448 _6224_/Q vssd1 vssd1 vccd1 vccd1 hold448/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 _6222_/Q vssd1 vssd1 vccd1 vccd1 hold437/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold459 _4723_/X vssd1 vssd1 vccd1 vccd1 _6069_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6212_ _6218_/CLK _6212_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6212_/Q sky130_fd_sc_hd__dfstp_1
X_3424_ _3277_/A _4070_/B _3434_/D hold377/X _3405_/B vssd1 vssd1 vccd1 vccd1 _3424_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _3363_/B vssd1 vssd1 vccd1 vccd1 _3368_/B sky130_fd_sc_hd__inv_2
X_6143_ _6190_/CLK hold49/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__5532__S _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ _6256_/CLK _6074_/D fanout175/X vssd1 vssd1 vccd1 vccd1 _6074_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3540_/A _4618_/C vssd1 vssd1 vccd1 vccd1 _3286_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5025_ _5025_/A _5448_/B vssd1 vssd1 vccd1 vccd1 _5026_/A sky130_fd_sc_hd__nor2_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout182_A fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5490__A0 _6236_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5793__A1 _6236_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5927_ _6035_/CLK _5927_/D vssd1 vssd1 vccd1 vccd1 _5927_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4391__B _4391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5793__B2 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3288__A _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5858_ _3864_/Y _5834_/X _5837_/X _5857_/X vssd1 vssd1 vccd1 vccd1 _5858_/X sky130_fd_sc_hd__o22a_1
XANTENNA__5707__S _5707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5789_ _6179_/Q hold474/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5789_/X sky130_fd_sc_hd__mux2_1
X_4809_ _4839_/C _4809_/B _4824_/B vssd1 vssd1 vccd1 vccd1 _4814_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5008__A _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold561_A _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5839__A2 _6117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4757__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3140_ _3140_/A _3478_/A _3477_/A _4772_/C vssd1 vssd1 vccd1 vccd1 _4413_/C sky130_fd_sc_hd__or4_1
X_3071_ _3556_/A _3694_/C vssd1 vssd1 vccd1 vccd1 _3127_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_82_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5712_ _4116_/Y _5711_/X _5762_/A vssd1 vssd1 vccd1 vccd1 _5713_/A sky130_fd_sc_hd__a21o_2
X_3973_ _3974_/A _3974_/C _3974_/B vssd1 vssd1 vccd1 vccd1 _3975_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__3786__B1 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3539__C _4726_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5643_ _5694_/A _5643_/B vssd1 vssd1 vccd1 vccd1 _5643_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5574_ hold431/X _5573_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _5574_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold201 _6021_/Q vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
X_4525_ _4524_/X _4523_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4821_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_25_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5473__D _6160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold212 _4262_/X vssd1 vssd1 vccd1 vccd1 _5927_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _5969_/Q vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 _3837_/X vssd1 vssd1 vccd1 vccd1 _5895_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _5952_/Q vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 _6218_/Q vssd1 vssd1 vccd1 vccd1 _5767_/B sky130_fd_sc_hd__buf_1
Xhold267 _6012_/Q vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold245 _3402_/B vssd1 vssd1 vccd1 vccd1 _5977_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4456_ _4478_/A _3517_/C _3519_/B vssd1 vssd1 vccd1 vccd1 _4456_/X sky130_fd_sc_hd__a21bo_1
Xhold289 _6015_/Q vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4502__A2 _4612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3407_ _3196_/B _4618_/C _5093_/B _3247_/Y _3184_/A vssd1 vssd1 vccd1 vccd1 _3407_/X
+ sky130_fd_sc_hd__a32o_1
X_4387_ _3050_/C _4070_/Y _3210_/C vssd1 vssd1 vccd1 vccd1 _4387_/X sky130_fd_sc_hd__a21o_1
X_3338_ _3540_/A _3307_/B _3337_/X _3457_/A vssd1 vssd1 vccd1 vccd1 _3338_/Y sky130_fd_sc_hd__a211oi_1
X_6126_ _6130_/CLK _6126_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6126_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5463__B1 _5363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6057_ _6060_/CLK _6057_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6057_/Q sky130_fd_sc_hd__dfrtp_4
X_3269_ _4770_/C vssd1 vssd1 vccd1 vccd1 _4771_/C sky130_fd_sc_hd__inv_2
X_5008_ _6243_/Q _5008_/B vssd1 vssd1 vccd1 vccd1 _5008_/X sky130_fd_sc_hd__and2_1
XANTENNA__4018__A1 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5766__B2 _3959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4341__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_21_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3295__A_N _6127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5757__B2 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6130__RESET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5290_ hold636/X _5253_/Y _5254_/Y hold591/X vssd1 vssd1 vccd1 vccd1 _5290_/X sky130_fd_sc_hd__a22o_1
X_4310_ _5297_/A _4355_/A vssd1 vssd1 vccd1 vccd1 _4318_/S sky130_fd_sc_hd__or2_4
XFILLER_0_10_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__5142__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4241_ hold254/X hold80/X hold133/X hold64/X _5179_/S _4255_/S vssd1 vssd1 vccd1
+ vccd1 _4241_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4172_ _4219_/A _4173_/B vssd1 vssd1 vccd1 vccd1 _4172_/Y sky130_fd_sc_hd__nand2_1
X_3123_ _3210_/A _3203_/D _4056_/B _3249_/A vssd1 vssd1 vccd1 vccd1 _3123_/X sky130_fd_sc_hd__o211a_1
X_3054_ _3210_/A _4485_/A _3426_/A _3203_/B vssd1 vssd1 vccd1 vccd1 _3182_/B sky130_fd_sc_hd__or4bb_4
XANTENNA__4799__A2 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5748__B2 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3956_ _3623_/X _5372_/A _3955_/X vssd1 vssd1 vccd1 vccd1 _3956_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout145_A _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4420__B2 _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5626_ _5626_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5661_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3887_ _3795_/C _3884_/X _3886_/X vssd1 vssd1 vccd1 vccd1 _3887_/Y sky130_fd_sc_hd__o21ai_1
X_5557_ _5556_/X _6057_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _5557_/X sky130_fd_sc_hd__mux2_1
X_5488_ hold601/X _5487_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _5488_/X sky130_fd_sc_hd__mux2_1
X_4508_ hold74/A hold94/A _5894_/Q _6006_/Q _5076_/A0 _4272_/B vssd1 vssd1 vccd1 vccd1
+ _4508_/X sky130_fd_sc_hd__mux4_1
XANTENNA__5133__C1 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4439_ _4439_/A _4439_/B vssd1 vssd1 vccd1 vccd1 _4439_/X sky130_fd_sc_hd__or2_1
X_6109_ _6218_/CLK hold32/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout58_A _3270_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4336__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5739__B2 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4411__A1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4411__B2 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3054__C_N _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3810_ _3767_/A _3767_/B _3765_/A vssd1 vssd1 vccd1 vccd1 _3811_/B sky130_fd_sc_hd__a21bo_1
X_4790_ _6055_/Q _4764_/X _4763_/B vssd1 vssd1 vccd1 vccd1 _4790_/X sky130_fd_sc_hd__a21o_1
XANTENNA__4402__A1 _5250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3741_ _3739_/X _3740_/X _4256_/S vssd1 vssd1 vccd1 vccd1 _3741_/X sky130_fd_sc_hd__mux2_1
XANTENNA_29 _6048_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_18 _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4953__A2 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3610__C1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3672_ hold91/A _6146_/Q _3740_/S vssd1 vssd1 vccd1 vccd1 _3672_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5411_ _3920_/A _5402_/X _5410_/Y vssd1 vssd1 vccd1 vccd1 _5411_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5342_ _5629_/A _5773_/B vssd1 vssd1 vccd1 vccd1 _5342_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4929__B _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5273_ _5773_/A hold400/X _5245_/Y _5272_/X vssd1 vssd1 vccd1 vccd1 _5273_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4224_ hold31/X _4253_/A2 _3927_/X _4223_/Y vssd1 vssd1 vccd1 vccd1 _4224_/X sky130_fd_sc_hd__o22a_1
X_4155_ _5946_/Q _3605_/X _3615_/X _6029_/Q _4154_/X vssd1 vssd1 vccd1 vccd1 _4156_/B
+ sky130_fd_sc_hd__a221o_1
X_3106_ _3203_/A _3148_/B _3148_/C _3210_/C vssd1 vssd1 vccd1 vccd1 _3208_/B sky130_fd_sc_hd__or4_4
X_4086_ _3112_/A _3192_/B _4094_/C _3210_/C vssd1 vssd1 vccd1 vccd1 _4086_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_77_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6052__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3037_ _3193_/A _6259_/Q _6258_/Q _4739_/A vssd1 vssd1 vccd1 vccd1 _3323_/C sky130_fd_sc_hd__or4b_2
XANTENNA__5792__A1_N _6236_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5197__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4988_ _4987_/X _6159_/Q _5704_/S vssd1 vssd1 vccd1 vccd1 _4988_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3939_ _6071_/Q _3939_/B vssd1 vssd1 vccd1 vccd1 _3939_/X sky130_fd_sc_hd__or2_1
XFILLER_0_46_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5609_ _5608_/X _6061_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _5609_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_46_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6130_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_61_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4555__S1 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4396__B1 _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3934__A _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5112__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4765__A _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4871__B2 _4865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4623__A1 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5960_ _6149_/CLK _5960_/D vssd1 vssd1 vccd1 vccd1 _5960_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4911_ _4990_/A _4915_/B vssd1 vssd1 vccd1 vccd1 _4911_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_2_0__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5891_ hold621/X _5875_/X _5876_/Y _5890_/X vssd1 vssd1 vccd1 vccd1 _5891_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4842_ _6208_/Q _4768_/Y _4769_/Y _4836_/B _4815_/B vssd1 vssd1 vccd1 vccd1 _4842_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4773_ _4735_/A _4614_/B _4728_/C _3483_/X _4772_/X vssd1 vssd1 vccd1 vccd1 _4774_/B
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4387__B1 _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3724_ hold90/A _5981_/Q _3724_/S vssd1 vssd1 vccd1 vccd1 _3724_/X sky130_fd_sc_hd__mux2_1
X_3655_ _6070_/Q _3655_/B vssd1 vssd1 vccd1 vccd1 _3950_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_43_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5762__C _5762_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3586_ _3573_/C _3986_/A2 _3584_/X _3585_/X vssd1 vssd1 vccd1 vccd1 _3793_/D sky130_fd_sc_hd__o31ai_4
X_5325_ hold657/X _5320_/S _5317_/Y hold38/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__a22o_1
X_5256_ _6204_/Q _5251_/Y _5252_/Y hold486/X _5255_/X vssd1 vssd1 vccd1 vccd1 _5256_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4207_ _4207_/A _4207_/B vssd1 vssd1 vccd1 vccd1 _5055_/C sky130_fd_sc_hd__xnor2_1
X_5187_ _6177_/Q _5104_/Y _5106_/Y _6209_/Q vssd1 vssd1 vccd1 vccd1 _5187_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3665__A2 _3664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4862__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4138_ _5937_/Q _5297_/B _4263_/A _5928_/Q vssd1 vssd1 vccd1 vccd1 _4138_/X sky130_fd_sc_hd__o22a_1
XANTENNA__3417__A2 _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4069_ _4069_/A _4069_/B _4069_/C vssd1 vssd1 vccd1 vccd1 _4069_/X sky130_fd_sc_hd__or3_1
XFILLER_0_53_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4225__S0 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4753__A2_N _5424_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold591_A _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout182 fanout183/X vssd1 vssd1 vccd1 vccd1 fanout182/X sky130_fd_sc_hd__clkbuf_8
Xfanout160 hold607/X vssd1 vssd1 vccd1 vccd1 _5164_/A1 sky130_fd_sc_hd__buf_4
Xfanout171 fanout172/X vssd1 vssd1 vccd1 vccd1 fanout171/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3408__A2 _4439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5869__A0 _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold608 _4724_/X vssd1 vssd1 vccd1 vccd1 _6070_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold619 _6038_/Q vssd1 vssd1 vccd1 vccd1 hold619/X sky130_fd_sc_hd__dlygate4sd3_1
X_3440_ _3143_/Y _4044_/B _4054_/C _3439_/Y _3457_/A vssd1 vssd1 vccd1 vccd1 _3440_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_100_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3371_ hold273/X _3353_/X _3372_/B vssd1 vssd1 vccd1 vccd1 _3371_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3383__B _3383_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6090_ _6227_/CLK _6090_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6090_/Q sky130_fd_sc_hd__dfrtp_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5957_/Q _3591_/A _3740_/S _5996_/Q _5179_/S vssd1 vssd1 vccd1 vccd1 _5114_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ _6113_/Q _3657_/A _5040_/X vssd1 vssd1 vccd1 vccd1 _5044_/B sky130_fd_sc_hd__a21o_1
XANTENNA__5097__A1 _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5103__B _5105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_wb_clk_i wb_clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_wb_clk_i/X sky130_fd_sc_hd__clkbuf_16
X_5943_ _6030_/CLK hold65/X vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5874_ hold652/X _4415_/A _5872_/A vssd1 vssd1 vccd1 vccd1 _5875_/C sky130_fd_sc_hd__a21o_1
X_4825_ _6191_/Q _6057_/Q _6038_/Q vssd1 vssd1 vccd1 vccd1 _4825_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3472__A1_N _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4756_ _5502_/A _4755_/Y _3513_/C vssd1 vssd1 vccd1 vccd1 _4926_/S sky130_fd_sc_hd__o21ai_4
X_4687_ _4699_/A _4688_/B vssd1 vssd1 vccd1 vccd1 _4687_/Y sky130_fd_sc_hd__nor2_1
X_3707_ _3706_/X hold484/X _3958_/S vssd1 vssd1 vccd1 vccd1 _3707_/X sky130_fd_sc_hd__mux2_4
X_3638_ _6072_/Q _3638_/B vssd1 vssd1 vccd1 vccd1 _3848_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_3_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4532__A0 _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3569_ _5711_/A _5021_/B _3569_/C vssd1 vssd1 vccd1 vccd1 _3569_/Y sky130_fd_sc_hd__nand3_2
X_5308_ input3/X hold631/X _5313_/S vssd1 vssd1 vccd1 vccd1 _6156_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_101_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4835__A1 _4834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5239_ _3275_/B _5107_/A _5120_/A vssd1 vssd1 vccd1 vccd1 _5239_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_98_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4063__A2 _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3271__B1 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4344__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold604_A _6127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3574__A1 _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4519__S _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output21_A _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5003__A1 _5007_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4610_ _4631_/B _4611_/C vssd1 vssd1 vccd1 vccd1 _4610_/X sky130_fd_sc_hd__and2_1
XFILLER_0_44_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5590_ _5590_/A _5590_/B vssd1 vssd1 vccd1 vccd1 _5590_/Y sky130_fd_sc_hd__xnor2_1
X_4541_ _4540_/X _4539_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4836_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold427 _6184_/Q vssd1 vssd1 vccd1 vccd1 hold427/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold405 _5785_/X vssd1 vssd1 vccd1 vccd1 _6231_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold416 _6139_/Q vssd1 vssd1 vccd1 vccd1 hold416/X sky130_fd_sc_hd__dlygate4sd3_1
X_4472_ _6154_/Q _4779_/B vssd1 vssd1 vccd1 vccd1 _4472_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_13_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold438 _5776_/X vssd1 vssd1 vccd1 vccd1 _6222_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 _5778_/X vssd1 vssd1 vccd1 vccd1 _6224_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6211_ _6211_/CLK _6211_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6211_/Q sky130_fd_sc_hd__dfstp_1
X_3423_ _4485_/B _3419_/X _3421_/Y _4415_/A _3422_/Y vssd1 vssd1 vccd1 vccd1 _3423_/X
+ sky130_fd_sc_hd__a221o_1
X_6142_ _6175_/CLK _6142_/D vssd1 vssd1 vccd1 vccd1 _6142_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _6129_/Q _6127_/Q hold50/X vssd1 vssd1 vccd1 vccd1 _3363_/B sky130_fd_sc_hd__or3_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3285_ _3396_/A _3479_/B vssd1 vssd1 vccd1 vccd1 _3285_/Y sky130_fd_sc_hd__nor2_1
X_6073_ _6170_/CLK _6073_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6073_/Q sky130_fd_sc_hd__dfrtp_4
X_5024_ _5024_/A _5024_/B vssd1 vssd1 vccd1 vccd1 _5448_/B sky130_fd_sc_hd__or2_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5114__A _5116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout175_A fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5926_ _6034_/CLK _5926_/D vssd1 vssd1 vccd1 vccd1 _5926_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5857_ _6117_/Q _5856_/X _5869_/S vssd1 vssd1 vccd1 vccd1 _5857_/X sky130_fd_sc_hd__mux2_1
X_5788_ _6178_/Q hold433/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5788_/X sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4808_ _6056_/Q _4823_/C vssd1 vssd1 vccd1 vccd1 _4809_/B sky130_fd_sc_hd__or2_1
XANTENNA__5545__A2 _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4753__B1 _4451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4739_ _4739_/A _4739_/B vssd1 vssd1 vccd1 vccd1 _4739_/X sky130_fd_sc_hd__or2_1
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5008__B _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4505__A0 _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4600__S0 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout88_A _4116_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4339__S _4345_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3243__S _6179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5481__A1 _6179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3492__B1 _4478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5678__B _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5233__A1 _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_50_wb_clk_i_A _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5233__B2 _6127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5694__A _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4992__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4744__B1 _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3942__A _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4757__B _4779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3070_ _3070_/A _3116_/A vssd1 vssd1 vccd1 vccd1 _4615_/B sky130_fd_sc_hd__nor2_1
XANTENNA__5472__A1 _5050_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5900__RESET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3389__A _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3972_ _3875_/B _3890_/B _4234_/A vssd1 vssd1 vccd1 vccd1 _3972_/X sky130_fd_sc_hd__o21a_1
X_5711_ _5711_/A _5711_/B vssd1 vssd1 vccd1 vccd1 _5711_/X sky130_fd_sc_hd__or2_2
X_5642_ _6064_/Q _5702_/A2 _5702_/B1 _5641_/X vssd1 vssd1 vccd1 vccd1 _5643_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_5_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5573_ _5566_/X _5572_/X _5670_/A vssd1 vssd1 vccd1 vccd1 _5573_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold202 _4357_/X vssd1 vssd1 vccd1 vccd1 _6021_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4524_ _5983_/Q _5991_/Q _5999_/Q _5960_/Q _5076_/A0 _4272_/B vssd1 vssd1 vccd1 vccd1
+ _4524_/X sky130_fd_sc_hd__mux4_1
Xhold224 _5947_/Q vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _6014_/Q vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 _5900_/Q vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 _5767_/Y vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 _6094_/Q vssd1 vssd1 vccd1 vccd1 _5426_/A sky130_fd_sc_hd__buf_1
Xhold246 _6018_/Q vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
X_4455_ _3405_/B _3349_/Y _5314_/A vssd1 vssd1 vccd1 vccd1 _4455_/X sky130_fd_sc_hd__o21a_1
Xhold279 _4291_/X vssd1 vssd1 vccd1 vccd1 _5952_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3406_ _3405_/B hold235/X _5502_/C _3434_/D _3404_/X vssd1 vssd1 vccd1 vccd1 _3406_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4386_ _5502_/B _4383_/Y _4385_/Y _3446_/A _4381_/Y vssd1 vssd1 vccd1 vccd1 _4386_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3337_ _3307_/A _3307_/B _3337_/C _3337_/D vssd1 vssd1 vccd1 vccd1 _3337_/X sky130_fd_sc_hd__and4bb_1
X_6125_ _6130_/CLK _6125_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6125_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _4415_/A _3268_/B _3268_/C vssd1 vssd1 vccd1 vccd1 _4770_/C sky130_fd_sc_hd__nor3_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ _6192_/CLK _6056_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6056_/Q sky130_fd_sc_hd__dfrtp_4
X_5007_ _5007_/A _5007_/B vssd1 vssd1 vccd1 vccd1 _5007_/Y sky130_fd_sc_hd__nand2_1
X_3199_ _4417_/A _3192_/B _3193_/X _3198_/Y _3210_/C vssd1 vssd1 vccd1 vccd1 _3200_/C
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_68_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5215__A1 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3299__A _5838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5909_ _6152_/CLK _5909_/D vssd1 vssd1 vccd1 vccd1 _5909_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold302_A _6048_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5453__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5454__A1 _6177_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4257__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3465__B1 _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5206__A1 _6179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3217__B1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5509__A2 _3370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5142__B1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4240_ hold5/X _4253_/A2 _3960_/Y _4239_/Y vssd1 vssd1 vccd1 vccd1 _4240_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4171_ _4171_/A _4171_/B vssd1 vssd1 vccd1 vccd1 _4173_/B sky130_fd_sc_hd__or2_2
X_3122_ _6130_/Q _4725_/B vssd1 vssd1 vccd1 vccd1 _3309_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3053_ _4398_/A _4417_/B vssd1 vssd1 vccd1 vccd1 _4117_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3471__A3 _5838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3955_ _3650_/X _5384_/A _3952_/X _3954_/X vssd1 vssd1 vccd1 vccd1 _3955_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5625_ _5317_/A _5670_/A _5672_/S vssd1 vssd1 vccd1 vccd1 _5625_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout138_A _6165_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3886_ _3582_/Y _3885_/X _3579_/Y vssd1 vssd1 vccd1 vccd1 _3886_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5381__B1 _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5556_ _4119_/B _5555_/X _4821_/Y vssd1 vssd1 vccd1 vccd1 _5556_/X sky130_fd_sc_hd__a21bo_1
X_5487_ _4030_/Y _5486_/X _5487_/S vssd1 vssd1 vccd1 vccd1 _5487_/X sky130_fd_sc_hd__mux2_1
X_4507_ _4589_/S _4507_/B vssd1 vssd1 vccd1 vccd1 _4512_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5133__B1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4438_ _3193_/A _4436_/X _4437_/X vssd1 vssd1 vccd1 vccd1 _4438_/X sky130_fd_sc_hd__a21o_1
XANTENNA__5684__B2 _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4369_ hold206/X _4211_/X _4372_/S vssd1 vssd1 vccd1 vccd1 _4369_/X sky130_fd_sc_hd__mux2_1
X_6108_ _6206_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ _6256_/CLK hold53/X fanout172/X vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dfrtp_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4947__A0 _4943_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4352__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4411__A2 _4409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3757__A _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5675__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3438__B1 _4043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3989__A1 _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4650__A2 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4938__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4402__A2 _4410_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_19 _5330_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3740_ hold88/A _5982_/Q _3740_/S vssd1 vssd1 vccd1 vccd1 _3740_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5882__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3671_ _6132_/Q _3671_/B vssd1 vssd1 vccd1 vccd1 _5209_/A sky130_fd_sc_hd__nand2_4
X_5410_ _2958_/Y _5026_/Y _5044_/X _5365_/S _5409_/X vssd1 vssd1 vccd1 vccd1 _5410_/Y
+ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5341_ _5341_/A _5457_/A vssd1 vssd1 vccd1 vccd1 _5773_/B sky130_fd_sc_hd__nand2_4
XFILLER_0_23_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4498__A _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5115__B1 _5185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5272_ _5248_/Y _5269_/X _5271_/X vssd1 vssd1 vccd1 vccd1 _5272_/X sky130_fd_sc_hd__a21o_1
X_4223_ _4223_/A _4223_/B vssd1 vssd1 vccd1 vccd1 _4223_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4154_ _5921_/Q _3588_/X _3603_/X _6013_/Q vssd1 vssd1 vccd1 vccd1 _4154_/X sky130_fd_sc_hd__a22o_1
X_3105_ _3105_/A _6258_/Q vssd1 vssd1 vccd1 vccd1 _4056_/A sky130_fd_sc_hd__nand2_4
X_4085_ _4124_/B _4085_/B vssd1 vssd1 vccd1 vccd1 _4094_/C sky130_fd_sc_hd__or2_1
X_3036_ _3193_/A _5502_/B _3276_/A _5502_/C vssd1 vssd1 vccd1 vccd1 _3483_/A sky130_fd_sc_hd__a211o_1
XFILLER_0_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4987_ _5694_/A _4986_/X _4976_/Y vssd1 vssd1 vccd1 vccd1 _4987_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_58_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3938_ _3935_/Y _3936_/X _3937_/Y vssd1 vssd1 vccd1 vccd1 _3938_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_46_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3869_ hold60/A _5910_/Q _3885_/S vssd1 vssd1 vccd1 vccd1 _3869_/X sky130_fd_sc_hd__mux2_1
X_5608_ _5694_/A _5607_/X _4879_/Y vssd1 vssd1 vccd1 vccd1 _5608_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5539_ _5540_/A _5540_/B _5538_/Y vssd1 vssd1 vccd1 vccd1 _5552_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6014_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4347__S _4354_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5686__B _5698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5178__S _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4396__A1 _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3487__A _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3199__A2 _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4148__A1 _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4810__S _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3950__A _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4765__B _6050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4910_ hold311/X _4909_/X _4927_/S vssd1 vssd1 vccd1 vccd1 _4910_/X sky130_fd_sc_hd__mux2_1
X_5890_ input8/X _5890_/B vssd1 vssd1 vccd1 vccd1 _5890_/X sky130_fd_sc_hd__and2_1
X_4841_ _4854_/B _4841_/B vssd1 vssd1 vccd1 vccd1 _4841_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_47_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4772_ _5502_/A _4772_/B _4772_/C _4772_/D vssd1 vssd1 vccd1 vccd1 _4772_/X sky130_fd_sc_hd__or4_1
XFILLER_0_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3723_ _3721_/X _3722_/X _3988_/A vssd1 vssd1 vccd1 vccd1 _3730_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_43_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3654_ _6136_/Q _3653_/X _3654_/S vssd1 vssd1 vccd1 vccd1 _5395_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_3_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3585_ _3513_/A _3571_/X _3559_/B _4963_/A vssd1 vssd1 vccd1 vccd1 _3585_/X sky130_fd_sc_hd__a211o_4
XFILLER_0_100_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4021__A _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5324_ hold38/X _5320_/S _5317_/Y _3539_/B vssd1 vssd1 vccd1 vccd1 _5324_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5255_ _6154_/Q _5253_/Y _5254_/Y _6236_/Q vssd1 vssd1 vccd1 vccd1 _5255_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4206_ _4206_/A _4206_/B vssd1 vssd1 vccd1 vccd1 _4207_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5186_ _5184_/X _5185_/X _5209_/A vssd1 vssd1 vccd1 vccd1 _5186_/X sky130_fd_sc_hd__mux2_1
X_4137_ _3972_/X _4135_/D _4135_/X _4136_/X vssd1 vssd1 vccd1 vccd1 _4145_/B sky130_fd_sc_hd__a211o_1
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4068_ _5502_/B _3127_/B _4043_/C _4048_/A _4067_/X vssd1 vssd1 vccd1 vccd1 _4069_/C
+ sky130_fd_sc_hd__a311o_1
XANTENNA__5811__A1 _3832_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6202__RESET_B fanout184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3822__A0 _6116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3019_ _6259_/Q _6258_/Q vssd1 vssd1 vccd1 vccd1 _4417_/A sky130_fd_sc_hd__or2_4
XFILLER_0_93_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4225__S1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3338__C1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4550__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout183 fanout184/X vssd1 vssd1 vccd1 vccd1 fanout183/X sky130_fd_sc_hd__buf_6
Xfanout161 _5936_/Q vssd1 vssd1 vccd1 vccd1 _4712_/S1 sky130_fd_sc_hd__clkbuf_8
Xfanout150 _4725_/B vssd1 vssd1 vccd1 vccd1 _3715_/B sky130_fd_sc_hd__buf_4
Xfanout172 input13/X vssd1 vssd1 vccd1 vccd1 fanout172/X sky130_fd_sc_hd__buf_4
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3010__A _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3041__A1 _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold609 _6071_/Q vssd1 vssd1 vccd1 vccd1 hold609/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3370_ _4077_/A _3370_/B _3370_/C vssd1 vssd1 vccd1 vccd1 _3372_/B sky130_fd_sc_hd__and3_1
XFILLER_0_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4776__A _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _6116_/Q _3827_/B _3695_/B _6114_/Q vssd1 vssd1 vccd1 vccd1 _5040_/X sky130_fd_sc_hd__a22o_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4057__B1 _4737_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5942_ _6031_/CLK hold73/X vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__dfxtp_1
X_5873_ input1/X _5890_/B vssd1 vssd1 vccd1 vccd1 _5873_/X sky130_fd_sc_hd__and2_1
XFILLER_0_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4824_ _4823_/X _4824_/B _4824_/C vssd1 vssd1 vccd1 vccd1 _4829_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4755_ _3167_/B _3283_/Y _4754_/X vssd1 vssd1 vccd1 vccd1 _4755_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5309__A0 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3706_ _6155_/Q _3705_/Y _6074_/Q vssd1 vssd1 vccd1 vccd1 _3706_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4780__A1 _4104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4686_ _6217_/Q _4976_/B _4714_/S vssd1 vssd1 vccd1 vccd1 _4688_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_31_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3637_ _6072_/Q _3638_/B vssd1 vssd1 vccd1 vccd1 _3647_/C sky130_fd_sc_hd__and2_2
XFILLER_0_3_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3568_ _4124_/B _5313_/S _3567_/Y vssd1 vssd1 vccd1 vccd1 _3569_/C sky130_fd_sc_hd__o21ai_1
X_5307_ input2/X hold632/X _5313_/S vssd1 vssd1 vccd1 vccd1 _6155_/D sky130_fd_sc_hd__mux2_1
X_3499_ _6127_/Q _5900_/Q _5901_/Q _4398_/B _3498_/Y vssd1 vssd1 vccd1 vccd1 _3499_/X
+ sky130_fd_sc_hd__a221o_1
X_5238_ _4077_/A _3353_/B _5217_/A hold586/X vssd1 vssd1 vccd1 vccd1 _5238_/X sky130_fd_sc_hd__a22o_1
X_5169_ _5169_/A _5169_/B vssd1 vssd1 vccd1 vccd1 _5169_/X sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_40_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4360__S _4363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6242_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__6195__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5787__A0 _6177_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4535__S _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5220__A _5220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4270__S _4271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4540_ _5984_/Q hold96/A _6000_/Q _5961_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4540_/X sky130_fd_sc_hd__mux4_1
Xhold406 _6140_/Q vssd1 vssd1 vccd1 vccd1 hold406/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 _5278_/X vssd1 vssd1 vccd1 vccd1 _6139_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4471_ _4589_/S _6154_/Q _4779_/B _4470_/X vssd1 vssd1 vccd1 vccd1 _4501_/A sky130_fd_sc_hd__a31o_1
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold428 _5494_/X vssd1 vssd1 vccd1 vccd1 _6184_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6210_ _6211_/CLK _6210_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6210_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5890__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold439 _6163_/Q vssd1 vssd1 vccd1 vccd1 _3461_/A sky130_fd_sc_hd__buf_2
XANTENNA__3317__A2 _5093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3422_ _3457_/A _3422_/B vssd1 vssd1 vccd1 vccd1 _3422_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6141_ _6175_/CLK _6141_/D vssd1 vssd1 vccd1 vccd1 _6141_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3722__C1 _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _5216_/A _3353_/B vssd1 vssd1 vccd1 vccd1 _3353_/X sky130_fd_sc_hd__or2_4
XFILLER_0_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _3715_/B _3283_/Y _3196_/B vssd1 vssd1 vccd1 vccd1 _3294_/A sky130_fd_sc_hd__o21a_1
X_6072_ _6086_/CLK _6072_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6072_/Q sky130_fd_sc_hd__dfrtp_4
X_5023_ _5023_/A _5023_/B vssd1 vssd1 vccd1 vccd1 _5051_/A sky130_fd_sc_hd__or2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5778__A0 _6240_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5925_ _6033_/CLK _5925_/D vssd1 vssd1 vccd1 vccd1 _5925_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5856_ _6135_/Q _6113_/Q _5868_/S vssd1 vssd1 vccd1 vccd1 _5856_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4807_ _6056_/Q _4823_/C vssd1 vssd1 vccd1 vccd1 _4839_/C sky130_fd_sc_hd__and2_1
XFILLER_0_90_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5787_ _6177_/Q hold443/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5787_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2999_ _2999_/A vssd1 vssd1 vccd1 vccd1 _2999_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_90_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4738_ _4738_/A _4738_/B _4738_/C _4738_/D vssd1 vssd1 vccd1 vccd1 _4738_/X sky130_fd_sc_hd__or4_1
X_4669_ _6024_/Q _5969_/Q _6016_/Q _5949_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4669_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_16_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_7_wb_clk_i_A _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4600__S1 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4992__B2 _4990_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5186__S _5209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4744__A1 _5164_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3468__D1 _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4265__S _4271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3971_ _4234_/A _3890_/B _3892_/B vssd1 vssd1 vccd1 vccd1 _3974_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__4983__A1 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3786__A2 _3785_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5710_ _4124_/B _6166_/Q _5875_/B vssd1 vssd1 vccd1 vccd1 _5711_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__4983__B2 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5641_ _6182_/Q _6198_/Q _5701_/S vssd1 vssd1 vccd1 vccd1 _5641_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5572_ _5584_/B _5572_/B vssd1 vssd1 vccd1 vccd1 _5572_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_53_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4523_ hold112/X _5909_/Q _5895_/Q _6007_/Q _5076_/A0 _4272_/B vssd1 vssd1 vccd1
+ vccd1 _4523_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold214 _6027_/Q vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 _6034_/Q vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold203 _5902_/Q vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold258 _5768_/Y vssd1 vssd1 vccd1 vccd1 _6218_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold269 _5057_/X vssd1 vssd1 vccd1 vccd1 _6094_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _4353_/X vssd1 vssd1 vccd1 vccd1 _6018_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 _3406_/X vssd1 vssd1 vccd1 vccd1 _5900_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4454_ _6048_/Q _3517_/C _3509_/Y _3517_/A vssd1 vssd1 vccd1 vccd1 _4454_/X sky130_fd_sc_hd__a22o_1
X_3405_ _5502_/A _3405_/B vssd1 vssd1 vccd1 vccd1 _3434_/D sky130_fd_sc_hd__nor2_2
X_4385_ _4385_/A _4385_/B vssd1 vssd1 vccd1 vccd1 _4385_/Y sky130_fd_sc_hd__nor2_1
X_6124_ _6129_/CLK _6124_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6124_/Q sky130_fd_sc_hd__dfstp_1
X_3336_ _3302_/A _3563_/A _4618_/C _3306_/A _3303_/A vssd1 vssd1 vccd1 vccd1 _3337_/C
+ sky130_fd_sc_hd__o311a_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ _6190_/CLK _6055_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6055_/Q sky130_fd_sc_hd__dfrtp_4
X_5006_ hold345/X _5005_/Y _5020_/S vssd1 vssd1 vccd1 vccd1 _5006_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3267_ _3220_/X _3258_/X _3266_/X _3211_/Y vssd1 vssd1 vccd1 vccd1 _3268_/C sky130_fd_sc_hd__a22oi_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3474__A1 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3198_ _3545_/A _3198_/B vssd1 vssd1 vccd1 vccd1 _3198_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__3299__B _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4903__S _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4974__A1 _6158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5908_ _6006_/CLK hold95/X vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfxtp_1
X_5839_ _3654_/S _6117_/Q _4022_/X vssd1 vssd1 vccd1 vccd1 _5839_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5151__A1 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5454__A2 _5352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3465__A1 _4750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4178__C1 _3671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5693__A2 _4761_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4170_ _5947_/Q _3605_/X _3615_/X _6030_/Q _4169_/X vssd1 vssd1 vccd1 vccd1 _4171_/B
+ sky130_fd_sc_hd__a221o_1
X_3121_ _4038_/A _4056_/A _4070_/B vssd1 vssd1 vccd1 vccd1 _3121_/X sky130_fd_sc_hd__and3_1
XFILLER_0_93_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3052_ _3052_/A _3081_/B _3178_/B vssd1 vssd1 vccd1 vccd1 _3396_/A sky130_fd_sc_hd__and3_2
XFILLER_0_77_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4956__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3954_ _4036_/B _3645_/X _3953_/X _6119_/Q vssd1 vssd1 vccd1 vccd1 _3954_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3847__B _6117_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3885_ _6001_/Q _5962_/Q _3885_/S vssd1 vssd1 vccd1 vccd1 _3885_/X sky130_fd_sc_hd__mux2_1
X_5624_ _5317_/A _5511_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _5624_/X sky130_fd_sc_hd__o21a_1
XANTENNA__4708__A1 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4959__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4184__A2 _3588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5555_ _6057_/Q _5595_/S _5607_/B1 _5554_/X vssd1 vssd1 vccd1 vccd1 _5555_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5554__S _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5486_ _6161_/Q _5475_/S _5482_/X _5485_/X vssd1 vssd1 vccd1 vccd1 _5486_/X sky130_fd_sc_hd__a22o_1
X_4506_ hold548/X _4505_/X _5296_/S vssd1 vssd1 vccd1 vccd1 _4506_/X sky130_fd_sc_hd__mux2_1
X_4437_ _5838_/A _3264_/X _4040_/B _4485_/B vssd1 vssd1 vccd1 vccd1 _4437_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_1_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4368_ hold173/X _4193_/X _4372_/S vssd1 vssd1 vccd1 vccd1 _4368_/X sky130_fd_sc_hd__mux2_1
X_6107_ _6218_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _3316_/X _3317_/X _3318_/X _4485_/B vssd1 vssd1 vccd1 vccd1 _3319_/Y sky130_fd_sc_hd__o31ai_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _3979_/X hold220/X _4300_/S vssd1 vssd1 vccd1 vccd1 _4299_/X sky130_fd_sc_hd__mux2_1
X_6038_ _6038_/CLK _6038_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _6038_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3103__A _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3013__A _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3610__A1 _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3386__C _5875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3670_ _6132_/Q _3671_/B vssd1 vssd1 vccd1 vccd1 _5116_/A sky130_fd_sc_hd__and2_4
XANTENNA__3683__A _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4779__A _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5340_ _5507_/A wire93/X vssd1 vssd1 vccd1 vccd1 _5340_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_50_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5271_ _6207_/Q _5251_/Y _5252_/Y _6215_/Q _5270_/X vssd1 vssd1 vccd1 vccd1 _5271_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5666__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4222_ _4222_/A _4222_/B vssd1 vssd1 vccd1 vccd1 _4223_/B sky130_fd_sc_hd__xnor2_1
X_4153_ hold62/A _3611_/X _3613_/X hold78/A _4152_/X vssd1 vssd1 vccd1 vccd1 _4156_/A
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4084_ _4084_/A _4084_/B _4084_/C vssd1 vssd1 vccd1 vccd1 _4084_/X sky130_fd_sc_hd__or3_1
X_3104_ _3105_/A _6258_/Q vssd1 vssd1 vccd1 vccd1 _4418_/A sky130_fd_sc_hd__and2_1
X_3035_ _3249_/A _3203_/C vssd1 vssd1 vccd1 vccd1 _3227_/B sky130_fd_sc_hd__or2_1
X_4986_ _6067_/Q _5702_/A2 _5607_/B1 _4985_/X vssd1 vssd1 vccd1 vccd1 _4986_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout150_A _4725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3937_ _3935_/Y _3936_/X _3647_/C vssd1 vssd1 vccd1 vccd1 _3937_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3868_ _6000_/Q _3603_/X _3605_/X _5961_/Q vssd1 vssd1 vccd1 vccd1 _3873_/B sky130_fd_sc_hd__a22o_1
XANTENNA__5284__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5607_ _6061_/Q _5595_/S _5607_/B1 _5606_/X vssd1 vssd1 vccd1 vccd1 _5607_/X sky130_fd_sc_hd__a22o_1
XANTENNA__6061__RESET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3799_ _3798_/B _3798_/C _3798_/D _4234_/A vssd1 vssd1 vccd1 vccd1 _3799_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_14_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5538_ _5538_/A _5538_/B vssd1 vssd1 vccd1 vccd1 _5538_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5469_ _6181_/Q _6180_/Q _6183_/Q _6182_/Q vssd1 vssd1 vccd1 vccd1 _5469_/X sky130_fd_sc_hd__or4_1
XANTENNA__3117__B1 _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3668__A1 _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout63_A _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4712__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4363__S _4363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3487__B _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5648__A2 _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5369__S _5484_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4840_ _6058_/Q _4823_/X _4824_/B vssd1 vssd1 vccd1 vccd1 _4841_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4771_ _4771_/A _4771_/B _4771_/C vssd1 vssd1 vccd1 vccd1 _4824_/B sky130_fd_sc_hd__and3_4
XFILLER_0_82_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3722_ _5893_/Q _3724_/S _3720_/X _3616_/B vssd1 vssd1 vccd1 vccd1 _3722_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5336__A1 _6172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3653_ _5356_/A _6172_/Q _5046_/A _3052_/A _4391_/B vssd1 vssd1 vccd1 vccd1 _3653_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3617__S _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5323_ _3539_/B _5320_/S _5317_/Y _4497_/S vssd1 vssd1 vccd1 vccd1 _6166_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3584_ hold48/A _3573_/B _3671_/B vssd1 vssd1 vccd1 vccd1 _3584_/X sky130_fd_sc_hd__o21a_4
X_5254_ _5289_/S _5254_/B vssd1 vssd1 vccd1 vccd1 _5254_/Y sky130_fd_sc_hd__nor2_2
X_4205_ _4250_/A _4205_/B vssd1 vssd1 vccd1 vccd1 _4206_/B sky130_fd_sc_hd__nand2_1
X_5185_ _3929_/X _4225_/X _5185_/S vssd1 vssd1 vccd1 vccd1 _5185_/X sky130_fd_sc_hd__mux2_1
X_4136_ _3970_/B _3990_/B _4234_/A vssd1 vssd1 vccd1 vccd1 _4136_/X sky130_fd_sc_hd__o21a_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_4067_ _4061_/A _4038_/A _4061_/C _4439_/B _4750_/A vssd1 vssd1 vccd1 vccd1 _4067_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__3822__A1 _6120_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3018_ _4398_/A _3022_/B vssd1 vssd1 vccd1 vccd1 _4728_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5279__S _5289_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3588__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4969_ _4824_/B _4967_/X _4968_/Y _4964_/X vssd1 vssd1 vccd1 vccd1 _4969_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_19_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4838__A0 _4836_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4358__S _4363_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout140 hold656/X vssd1 vssd1 vccd1 vccd1 _3591_/A sky130_fd_sc_hd__buf_4
Xfanout151 hold592/X vssd1 vssd1 vccd1 vccd1 _4725_/B sky130_fd_sc_hd__clkbuf_4
Xfanout173 fanout176/X vssd1 vssd1 vccd1 vccd1 fanout173/X sky130_fd_sc_hd__clkbuf_8
Xfanout162 hold647/X vssd1 vssd1 vccd1 vccd1 _4272_/B sky130_fd_sc_hd__clkbuf_8
Xfanout184 input13/X vssd1 vssd1 vccd1 vccd1 fanout184/X sky130_fd_sc_hd__buf_4
XFILLER_0_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3010__B _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5218__A _5220_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4268__S _4271_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3680__B _6114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4057__A1 _5424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5888__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5941_ _6014_/CLK hold71/X vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_wb_clk_i _5978_/CLK vssd1 vssd1 vccd1 vccd1 _6151_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5872_ _5872_/A _5872_/B vssd1 vssd1 vccd1 vccd1 _5890_/B sky130_fd_sc_hd__nand2_2
X_4823_ _6056_/Q _6057_/Q _4823_/C vssd1 vssd1 vccd1 vccd1 _4823_/X sky130_fd_sc_hd__and3_1
XFILLER_0_7_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4754_ _4759_/B _3396_/D _3711_/B _4753_/X vssd1 vssd1 vccd1 vccd1 _4754_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3705_ _3705_/A vssd1 vssd1 vccd1 vccd1 _3705_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4685_ _4684_/X _4683_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4976_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout113_A _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3636_ _3636_/A _3636_/B vssd1 vssd1 vccd1 vccd1 _3636_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4967__A _6158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5562__S _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3567_ _4124_/B _4497_/S vssd1 vssd1 vccd1 vccd1 _3567_/Y sky130_fd_sc_hd__nand2_1
X_5306_ input1/X hold637/X _5313_/S vssd1 vssd1 vccd1 vccd1 _6154_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3498_ _3498_/A _3498_/B vssd1 vssd1 vccd1 vccd1 _3498_/Y sky130_fd_sc_hd__nor2_1
X_5237_ _4077_/A _5222_/C _5228_/X _5218_/X _4474_/A vssd1 vssd1 vccd1 vccd1 _5237_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5493__A0 _6239_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5168_ _5896_/Q _3591_/A _3739_/S _6008_/Q _5179_/S vssd1 vssd1 vccd1 vccd1 _5169_/B
+ sky130_fd_sc_hd__o221a_1
XANTENNA__4906__S _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5099_ _3302_/A _5098_/X _5097_/X _5094_/X vssd1 vssd1 vccd1 vccd1 _5099_/X sky130_fd_sc_hd__a211o_1
X_4119_ _4119_/A _4119_/B vssd1 vssd1 vccd1 vccd1 _4121_/B sky130_fd_sc_hd__nand2_1
XANTENNA__5796__A1 _3664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3484__C _3488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5720__A1 _3707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3731__B1 _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3021__A _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4551__S _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold418 _6043_/Q vssd1 vssd1 vccd1 vccd1 _5327_/B sky130_fd_sc_hd__clkbuf_2
Xhold407 _5283_/X vssd1 vssd1 vccd1 vccd1 _6140_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4470_ _4589_/S _6204_/Q vssd1 vssd1 vccd1 vccd1 _4470_/X sky130_fd_sc_hd__and2b_1
XANTENNA__3504__C_N _5216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold429 _6230_/Q vssd1 vssd1 vccd1 vccd1 hold429/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3421_ _3428_/B vssd1 vssd1 vccd1 vccd1 _3421_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_40_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6140_ _6175_/CLK _6140_/D vssd1 vssd1 vccd1 vccd1 _6140_/Q sky130_fd_sc_hd__dfxtp_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3352_ _5216_/A _3353_/B vssd1 vssd1 vccd1 vccd1 _3370_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3283_/A _5093_/B vssd1 vssd1 vccd1 vccd1 _3283_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_29_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6071_ _6170_/CLK _6071_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6071_/Q sky130_fd_sc_hd__dfrtp_4
X_5022_ _3533_/S _3496_/X _5052_/D vssd1 vssd1 vccd1 vccd1 _5023_/B sky130_fd_sc_hd__o21ba_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5924_ _6032_/CLK _5924_/D vssd1 vssd1 vccd1 vccd1 _5924_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5855_ hold355/X _5836_/A _5854_/X _5773_/A vssd1 vssd1 vccd1 vccd1 _5855_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5557__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4806_ _6056_/Q _4764_/X _4763_/B vssd1 vssd1 vccd1 vccd1 _4806_/X sky130_fd_sc_hd__a21o_1
X_5786_ _6176_/Q hold514/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5786_/X sky130_fd_sc_hd__mux2_1
X_2998_ _6212_/Q vssd1 vssd1 vccd1 vccd1 _2998_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4737_ _4737_/A _4737_/B vssd1 vssd1 vccd1 vccd1 _4738_/D sky130_fd_sc_hd__nor2_1
X_4668_ hold70/A hold68/A _5924_/Q _6032_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4668_/X sky130_fd_sc_hd__mux4_1
X_3619_ _3617_/X _3618_/X _3983_/S vssd1 vssd1 vccd1 vccd1 _3619_/X sky130_fd_sc_hd__mux2_1
X_4599_ hold534/X _4598_/X _5073_/S vssd1 vssd1 vccd1 vccd1 _4599_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3492__A2 _3503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5769__B2 _4119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4371__S _4372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3016__A _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4680__A1 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3970_ _4234_/A _3970_/B vssd1 vssd1 vccd1 vccd1 _3974_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__4432__A1 _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5640_ _5660_/A _5640_/B vssd1 vssd1 vccd1 vccd1 _5640_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_72_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5571_ _5571_/A _5571_/B _5569_/Y vssd1 vssd1 vccd1 vccd1 _5572_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_5_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4522_ _4589_/S _4522_/B vssd1 vssd1 vccd1 vccd1 _4527_/B sky130_fd_sc_hd__nand2_1
Xhold215 _4363_/X vssd1 vssd1 vccd1 vccd1 _6027_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold226 _4371_/X vssd1 vssd1 vccd1 vccd1 _6034_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold204 _3400_/X vssd1 vssd1 vccd1 vccd1 _5902_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4453_ _3405_/B hold494/X _3434_/D _4750_/A vssd1 vssd1 vccd1 vccd1 _4453_/X sky130_fd_sc_hd__a22o_1
Xhold248 _5968_/Q vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold237 _5983_/Q vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4499__A1 _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold259 _5959_/Q vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
X_3404_ _4433_/A _5838_/B _5489_/D vssd1 vssd1 vccd1 vccd1 _3404_/X sky130_fd_sc_hd__o21a_2
X_4384_ _4737_/A _5502_/D _5838_/C _4044_/B _3545_/A vssd1 vssd1 vccd1 vccd1 _4384_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__5840__S _5869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3335_ _3317_/X _3325_/X _3334_/X _4485_/B vssd1 vssd1 vccd1 vccd1 _3335_/X sky130_fd_sc_hd__o31a_1
X_6123_ _6123_/CLK _6123_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6123_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ _6192_/CLK _6054_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6054_/Q sky130_fd_sc_hd__dfrtp_4
X_3266_ _3540_/A _3422_/B _3265_/X vssd1 vssd1 vccd1 vccd1 _3266_/X sky130_fd_sc_hd__o21a_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5704_/S _5003_/X _5004_/Y vssd1 vssd1 vccd1 vccd1 _5005_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__4120__B1 _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4671__A1 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout180_A fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3197_ _3395_/B _3197_/B _4484_/A vssd1 vssd1 vccd1 vccd1 _3200_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5907_ _6146_/CLK _5907_/D vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5838_ _5838_/A _5838_/B _5838_/C vssd1 vssd1 vccd1 vccd1 _5869_/S sky130_fd_sc_hd__and3_4
X_5769_ _4718_/A _4718_/B _5711_/X _5007_/B _4119_/A vssd1 vssd1 vccd1 vccd1 _5769_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_0_8_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5439__B1 _5363_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4366__S _4372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3465__A2 _5507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4414__B2 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3925__A0 _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5142__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3153__A1 _6130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3120_ _4486_/A _3120_/B vssd1 vssd1 vccd1 vccd1 _4729_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_93_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5250__C_N _4409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3051_ _6252_/Q _6259_/Q _6258_/Q vssd1 vssd1 vccd1 vccd1 _3178_/B sky130_fd_sc_hd__and3_1
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5697__A1_N _5707_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3953_ _4036_/B _3646_/X _3950_/Y _3645_/X vssd1 vssd1 vccd1 vccd1 _3953_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3884_ _5985_/Q _5993_/Q _3885_/S vssd1 vssd1 vccd1 vccd1 _3884_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5623_ _5613_/A _5622_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _5623_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4959__B _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5381__A2 _6046_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5554_ _6057_/Q _6191_/Q _5606_/S vssd1 vssd1 vccd1 vccd1 _5554_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5485_ _5365_/S _5484_/X _5363_/B vssd1 vssd1 vccd1 vccd1 _5485_/X sky130_fd_sc_hd__o21a_1
X_4505_ _6155_/Q _4504_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4505_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5133__A2 _5200_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4436_ _4118_/A _4430_/X _4431_/X _4415_/A _4435_/Y vssd1 vssd1 vccd1 vccd1 _4436_/X
+ sky130_fd_sc_hd__a221o_1
X_4367_ hold255/X _4180_/X _4372_/S vssd1 vssd1 vccd1 vccd1 _6030_/D sky130_fd_sc_hd__mux2_1
X_6106_ _6206_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__4892__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3318_ _4116_/B _3709_/B _3298_/Y vssd1 vssd1 vccd1 vccd1 _3318_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _3930_/X hold187/X _4300_/S vssd1 vssd1 vccd1 vccd1 _4298_/X sky130_fd_sc_hd__mux2_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ _3249_/A _3249_/B vssd1 vssd1 vccd1 vccd1 _3250_/D sky130_fd_sc_hd__nor2_1
X_6037_ _6086_/CLK hold47/X fanout174/X vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__4914__S _5216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3907__B1 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5124__A2 _5115_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5046__A _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold590 _5914_/Q vssd1 vssd1 vccd1 vccd1 hold590/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5832__A0 hold591/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4635__A1 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5919__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3013__B _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4938__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4399__B1 _5838_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4494__S0 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5655__S _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4779__B _4779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5270_ _6157_/Q _5253_/Y _5254_/Y _6239_/Q vssd1 vssd1 vccd1 vccd1 _5270_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5115__A2 _5209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4221_ _4207_/A _4207_/B _4206_/A vssd1 vssd1 vccd1 vccd1 _4222_/B sky130_fd_sc_hd__o21a_1
XANTENNA__4874__A1 _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4152_ _6021_/Q _3599_/X _3601_/X _5966_/Q vssd1 vssd1 vccd1 vccd1 _4152_/X sky130_fd_sc_hd__a22o_1
X_4083_ _3210_/A _4750_/B _4082_/X vssd1 vssd1 vccd1 vccd1 _4084_/C sky130_fd_sc_hd__a21o_1
X_3103_ _4398_/A _4739_/A _3116_/A _3125_/C vssd1 vssd1 vccd1 vccd1 _3157_/C sky130_fd_sc_hd__or4_1
XFILLER_0_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3034_ _3249_/A _3203_/C vssd1 vssd1 vccd1 vccd1 _5502_/C sky130_fd_sc_hd__nor2_2
XANTENNA__3834__C1 _3671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4985_ _6185_/Q _4984_/X _5701_/S vssd1 vssd1 vccd1 vccd1 _4985_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3936_ _3900_/A _3900_/B _3898_/A vssd1 vssd1 vccd1 vccd1 _3936_/X sky130_fd_sc_hd__a21o_1
XANTENNA_fanout143_A _4451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3867_ _5984_/Q _3599_/X _3601_/X hold96/X vssd1 vssd1 vccd1 vccd1 _3873_/A sky130_fd_sc_hd__a22o_1
XANTENNA__3874__A _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5565__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5606_ _6061_/Q _6195_/Q _5606_/S vssd1 vssd1 vccd1 vccd1 _5606_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3798_ _4234_/A _3798_/B _3798_/C _3798_/D vssd1 vssd1 vccd1 vccd1 _3798_/X sky130_fd_sc_hd__or4_1
XANTENNA__3904__A3 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5537_ _5537_/A vssd1 vssd1 vccd1 vccd1 _5552_/A sky130_fd_sc_hd__inv_2
XFILLER_0_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5468_ _6185_/Q _6184_/Q _6187_/Q _6186_/Q vssd1 vssd1 vccd1 vccd1 _5468_/X sky130_fd_sc_hd__or4_1
XFILLER_0_78_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4909__S _4926_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5399_ _5399_/A _5399_/B vssd1 vssd1 vccd1 vccd1 _5400_/B sky130_fd_sc_hd__xnor2_1
X_4419_ _4069_/B _4750_/C _4418_/X _4037_/X vssd1 vssd1 vccd1 vccd1 _4419_/X sky130_fd_sc_hd__o31a_1
XFILLER_0_96_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4712__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5290__A1 hold636/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5290__B2 hold591/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4093__A2 _4750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold522_A _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5042__A1 _6119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6194_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5042__B2 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5345__A2 _5343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6189__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4819__S _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3959__A _3959_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4467__S0 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4770_ _4770_/A _4770_/B _4770_/C vssd1 vssd1 vccd1 vccd1 _5008_/B sky130_fd_sc_hd__and3_4
XANTENNA__4792__A0 _6189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3721_ _6146_/Q _3724_/S _3719_/X _3983_/S vssd1 vssd1 vccd1 vccd1 _3721_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_99_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3652_ _6072_/Q _3652_/B _6073_/Q vssd1 vssd1 vccd1 vccd1 _3920_/A sky130_fd_sc_hd__and3b_4
XANTENNA__5336__A2 _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3583_ _3573_/C _3577_/S _3580_/X _3581_/X vssd1 vssd1 vccd1 vccd1 _3795_/C sky130_fd_sc_hd__o31a_2
X_5322_ _4497_/S _5320_/S _5317_/Y _3383_/A vssd1 vssd1 vccd1 vccd1 _6165_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5253_ _5259_/B _5254_/B vssd1 vssd1 vccd1 vccd1 _5253_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__4847__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4204_ _4250_/A _4205_/B vssd1 vssd1 vccd1 vccd1 _4206_/A sky130_fd_sc_hd__or2_1
X_5184_ _5180_/X _5183_/X _5185_/S vssd1 vssd1 vccd1 vccd1 _5184_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3315__A1_N _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4135_ _4135_/A _4135_/B _4135_/C _4135_/D vssd1 vssd1 vccd1 vccd1 _4135_/X sky130_fd_sc_hd__and4_1
XFILLER_0_64_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4066_ _4737_/A _5502_/D _4054_/C _4065_/X vssd1 vssd1 vccd1 vccd1 _4069_/B sky130_fd_sc_hd__a31o_1
X_3017_ _3507_/C _3137_/A vssd1 vssd1 vccd1 vccd1 _3022_/B sky130_fd_sc_hd__or2_1
XANTENNA__3588__B _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4968_ _4995_/C _4966_/Y _5013_/S vssd1 vssd1 vccd1 vccd1 _4968_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5575__A2 _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4899_ _4895_/B _4898_/X _4963_/A vssd1 vssd1 vccd1 vccd1 _4899_/X sky130_fd_sc_hd__mux2_1
X_3919_ _6139_/Q _6141_/Q _5868_/S vssd1 vssd1 vccd1 vccd1 _5397_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5295__S _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout130 hold625/X vssd1 vssd1 vccd1 vccd1 _3050_/C sky130_fd_sc_hd__buf_2
Xfanout141 _6131_/Q vssd1 vssd1 vccd1 vccd1 _5200_/A2 sky130_fd_sc_hd__buf_4
Xfanout152 _6112_/Q vssd1 vssd1 vccd1 vccd1 _4712_/S0 sky130_fd_sc_hd__buf_6
Xfanout163 hold588/X vssd1 vssd1 vccd1 vccd1 _4415_/A sky130_fd_sc_hd__buf_6
Xfanout174 fanout175/X vssd1 vssd1 vccd1 vccd1 fanout174/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__5263__A1 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3501__A1 _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4057__A2 _4446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5940_ _6035_/CLK hold83/X vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__4284__S _4291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5871_ hold386/X _5836_/A _5870_/X _5773_/A vssd1 vssd1 vccd1 vccd1 _5871_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_47_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4822_ _6057_/Q _4839_/C vssd1 vssd1 vccd1 vccd1 _4824_/C sky130_fd_sc_hd__or2_1
XFILLER_0_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4753_ _3185_/C _5424_/C _4451_/C _4728_/A vssd1 vssd1 vccd1 vccd1 _4753_/X sky130_fd_sc_hd__a2bb2o_1
X_3704_ _3704_/A _3704_/B vssd1 vssd1 vccd1 vccd1 _3705_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4684_ _6025_/Q _5970_/Q _6017_/Q _5950_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4684_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5843__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3635_ _3636_/A _3636_/B vssd1 vssd1 vccd1 vccd1 _3635_/X sky130_fd_sc_hd__or2_1
XANTENNA__4967__B _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3566_ _3457_/A _3560_/X _3565_/X vssd1 vssd1 vccd1 vccd1 _5021_/B sky130_fd_sc_hd__a21oi_2
X_3497_ _5900_/Q _5902_/Q _5901_/Q _5903_/Q vssd1 vssd1 vccd1 vccd1 _3498_/B sky130_fd_sc_hd__or4_1
X_5305_ hold76/X _4034_/X _5305_/S vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__mux2_1
XANTENNA__5144__A _5209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5236_ _4474_/A _5216_/B _5217_/Y hold518/X vssd1 vssd1 vccd1 vccd1 _5236_/X sky130_fd_sc_hd__o22a_1
X_5167_ _6000_/Q _5200_/A2 _5200_/B1 _5961_/Q _3594_/Y vssd1 vssd1 vccd1 vccd1 _5169_/A
+ sky130_fd_sc_hd__o221a_1
X_5098_ _3488_/A _5498_/B _3448_/Y _3082_/Y vssd1 vssd1 vccd1 vccd1 _5098_/X sky130_fd_sc_hd__a211o_1
X_4118_ _4118_/A _4118_/B vssd1 vssd1 vccd1 vccd1 _4118_/Y sky130_fd_sc_hd__nand2_1
X_4049_ _4056_/A _4048_/A _3556_/A vssd1 vssd1 vccd1 vccd1 _4049_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4223__A _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5720__A2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4369__S _4372_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4692__C1 _4619_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5236__A1 _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3302__A _3302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold408 _6120_/Q vssd1 vssd1 vccd1 vccd1 hold408/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold419 _6137_/Q vssd1 vssd1 vccd1 vccd1 hold419/X sky130_fd_sc_hd__dlygate4sd3_1
X_3420_ _4094_/B _4070_/B vssd1 vssd1 vccd1 vccd1 _3428_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_40_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3351_ _3353_/B vssd1 vssd1 vccd1 vccd1 _5216_/B sky130_fd_sc_hd__inv_2
XFILLER_0_21_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3543_/A _4427_/A vssd1 vssd1 vccd1 vccd1 _3334_/A sky130_fd_sc_hd__or2_1
X_6070_ _6170_/CLK _6070_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6070_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _3559_/A _5021_/B _5021_/C vssd1 vssd1 vccd1 vccd1 _5052_/D sky130_fd_sc_hd__and3b_2
XANTENNA__3789__A1 _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4986__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5923_ _6014_/CLK _5923_/D vssd1 vssd1 vccd1 vccd1 _5923_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5854_ _3832_/Y _5834_/X _5837_/X _5853_/X vssd1 vssd1 vccd1 vccd1 _5854_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_75_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4805_ _4990_/A _4805_/B vssd1 vssd1 vccd1 vccd1 _4805_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_90_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5785_ hold404/X _6231_/Q _5789_/S vssd1 vssd1 vccd1 vccd1 _5785_/X sky130_fd_sc_hd__mux2_1
X_2997_ _6062_/Q vssd1 vssd1 vccd1 vccd1 _4901_/A sky130_fd_sc_hd__inv_2
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4736_ _3097_/Y _4725_/X _4735_/Y _4445_/Y _4749_/A vssd1 vssd1 vccd1 vccd1 _4738_/C
+ sky130_fd_sc_hd__a221o_1
X_4667_ hold480/X _4666_/Y _5073_/S vssd1 vssd1 vccd1 vccd1 _4667_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5573__S _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5702__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3618_ hold130/X hold116/X _3724_/S vssd1 vssd1 vccd1 vccd1 _3618_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_101_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4598_ _6161_/Q _4597_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4598_/X sky130_fd_sc_hd__mux2_1
X_3549_ _3545_/Y _3547_/X _3548_/Y _3541_/X vssd1 vssd1 vccd1 vccd1 _3549_/X sky130_fd_sc_hd__a31o_1
X_6199_ _6238_/CLK _6199_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6199_/Q sky130_fd_sc_hd__dfrtp_4
X_5219_ _6075_/Q _6076_/Q vssd1 vssd1 vccd1 vccd1 _5219_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_98_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold268_A _6094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3122__A _6130_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold435_A _6115_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2961__A _6127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3952__A1 _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3265__A_N _3264_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3468__B1 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4968__B1 _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5570_ _5571_/A _5571_/B _5569_/Y vssd1 vssd1 vccd1 vccd1 _5584_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4521_ hold542/X _4520_/X _5296_/S vssd1 vssd1 vccd1 vccd1 _4521_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5145__B1 _5185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold205 _5984_/Q vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 _6150_/Q vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4452_ _5164_/A1 hold192/X _4450_/X _4451_/X vssd1 vssd1 vccd1 vccd1 _4452_/X sky130_fd_sc_hd__a22o_1
Xhold249 _4305_/X vssd1 vssd1 vccd1 vccd1 _5968_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 _5966_/Q vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 _6011_/Q vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
X_3403_ _3405_/B _5424_/B vssd1 vssd1 vccd1 vccd1 _5489_/D sky130_fd_sc_hd__nor2_2
XANTENNA__3207__A _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4383_ _3556_/A _4061_/A _4038_/A _4385_/B vssd1 vssd1 vccd1 vccd1 _4383_/Y sky130_fd_sc_hd__a31oi_2
X_3334_ _3334_/A _3334_/B _3334_/C _3334_/D vssd1 vssd1 vccd1 vccd1 _3334_/X sky130_fd_sc_hd__or4_1
XFILLER_0_0_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6122_ _6171_/CLK _6122_/D fanout173/X vssd1 vssd1 vccd1 vccd1 _6122_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3264_/X _3265_/B _3439_/B _5502_/A vssd1 vssd1 vccd1 vccd1 _3265_/X sky130_fd_sc_hd__and4b_1
X_6053_ _6144_/CLK _6053_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _6053_/Q sky130_fd_sc_hd__dfrtp_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5004_ _6160_/Q _5704_/S vssd1 vssd1 vccd1 vccd1 _5004_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4120__A1 _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _3396_/A _3196_/B vssd1 vssd1 vccd1 vccd1 _4484_/A sky130_fd_sc_hd__or2_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout173_A fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4038__A _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6055__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5620__A1 _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3877__A _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5906_ _6151_/CLK hold87/X vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5837_ _5837_/A _5837_/B vssd1 vssd1 vccd1 vccd1 _5837_/X sky130_fd_sc_hd__or2_2
XANTENNA__6175__SET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5768_ _5767_/A _5766_/X hold257/X vssd1 vssd1 vccd1 vccd1 _5768_/Y sky130_fd_sc_hd__o21ai_1
X_4719_ hold458/X _4612_/B _4718_/X _4474_/X vssd1 vssd1 vccd1 vccd1 _4719_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_16_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5699_ _5687_/A _5691_/A _5698_/Y vssd1 vssd1 vccd1 vccd1 _5699_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5803__A1_N _6238_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_wb_clk_i _5978_/CLK vssd1 vssd1 vccd1 vccd1 _6038_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__3698__B1 _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2956__A _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5478__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5507__A _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4886__C1 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3153__A2 _4725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4557__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_10_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3050_ _3210_/A _4485_/A _3050_/C vssd1 vssd1 vccd1 vccd1 _3081_/B sky130_fd_sc_hd__and3b_1
XANTENNA__5850__A1 _3785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4102__B2 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3952_ _6141_/Q _3648_/A _3920_/A _5394_/A _3624_/Y vssd1 vssd1 vccd1 vccd1 _3952_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3883_ _5897_/Q _3588_/X _3615_/X _6009_/Q vssd1 vssd1 vccd1 vccd1 _3888_/B sky130_fd_sc_hd__a22o_1
XFILLER_0_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5622_ _5621_/X _5616_/Y _5670_/A vssd1 vssd1 vccd1 vccd1 _5622_/X sky130_fd_sc_hd__mux2_1
X_5553_ _5552_/A _5552_/B _5552_/C vssd1 vssd1 vccd1 vccd1 _5571_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4504_ _4502_/X _4503_/X _5872_/A vssd1 vssd1 vccd1 vccd1 _4504_/X sky130_fd_sc_hd__mux2_1
X_5484_ _5483_/X hold361/X _5484_/S vssd1 vssd1 vccd1 vccd1 _5484_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4435_ _5424_/B _4435_/B vssd1 vssd1 vccd1 vccd1 _4435_/Y sky130_fd_sc_hd__nor2_1
X_4366_ hold252/X _4165_/X _4372_/S vssd1 vssd1 vccd1 vccd1 _6029_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6105_ _6208_/CLK hold37/X vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dfxtp_1
X_3317_ _3283_/A _5093_/B _3498_/A _3196_/B vssd1 vssd1 vccd1 vccd1 _3317_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ _3880_/X hold262/X _4300_/S vssd1 vssd1 vccd1 vccd1 _5961_/D sky130_fd_sc_hd__mux2_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3498_/A _3511_/C _4117_/C vssd1 vssd1 vccd1 vccd1 _3298_/A sky130_fd_sc_hd__and3_2
X_6036_ _6086_/CLK _6036_/D fanout174/X vssd1 vssd1 vccd1 vccd1 _6036_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__4991__A _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5841__A1 _3664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3179_ _3210_/A _4398_/A _4038_/B _3203_/B _4485_/A vssd1 vssd1 vccd1 vccd1 _3543_/A
+ sky130_fd_sc_hd__o2111a_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5298__S _5305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5109__B1 _5085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4580__B2 _4474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold580 _6257_/Q vssd1 vssd1 vccd1 vccd1 hold580/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold591 _6243_/Q vssd1 vssd1 vccd1 vccd1 hold591/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__4096__B1 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4399__A1 _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4494__S1 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4220_ _4220_/A _4220_/B vssd1 vssd1 vccd1 vccd1 _4222_/A sky130_fd_sc_hd__nand2_1
XANTENNA__3126__A2 _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4287__S _4291_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4151_ hold177/X _4150_/X _4262_/S vssd1 vssd1 vccd1 vccd1 _4151_/X sky130_fd_sc_hd__mux2_1
X_4082_ _3556_/A _3477_/B _3543_/B _4416_/A _4094_/B vssd1 vssd1 vccd1 vccd1 _4082_/X
+ sky130_fd_sc_hd__a311o_1
X_3102_ _4735_/A _3113_/B _3125_/C _3203_/D vssd1 vssd1 vccd1 vccd1 _3157_/B sky130_fd_sc_hd__or4_1
XANTENNA__3204__B _3370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3033_ _4735_/A _3249_/B vssd1 vssd1 vccd1 vccd1 _3203_/C sky130_fd_sc_hd__or2_1
XFILLER_0_77_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4984_ _6201_/Q _4815_/B _4978_/X _4983_/X vssd1 vssd1 vccd1 vccd1 _4984_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_58_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3935_ _3939_/B _3935_/B vssd1 vssd1 vccd1 vccd1 _3935_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5605_ _5603_/X _5605_/B vssd1 vssd1 vccd1 vccd1 _5605_/X sky130_fd_sc_hd__and2b_1
X_3866_ _3759_/A _5052_/B _3798_/X _3799_/X _3756_/Y vssd1 vssd1 vccd1 vccd1 _4135_/A
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_46_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3797_ _3798_/B _3798_/C _3798_/D vssd1 vssd1 vccd1 vccd1 _3800_/B sky130_fd_sc_hd__or3_2
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5536_ _5538_/A _5538_/B vssd1 vssd1 vccd1 vccd1 _5537_/A sky130_fd_sc_hd__nor2_1
XANTENNA__4051__A _4725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5467_ _6234_/Q _6178_/Q _5773_/B vssd1 vssd1 vccd1 vccd1 _5467_/X sky130_fd_sc_hd__mux2_1
X_4418_ _4418_/A _4750_/B _4418_/C _4417_/X vssd1 vssd1 vccd1 vccd1 _4418_/X sky130_fd_sc_hd__or4b_1
X_5398_ _5398_/A _5398_/B vssd1 vssd1 vccd1 vccd1 _5399_/B sky130_fd_sc_hd__xnor2_1
X_4349_ _4180_/X hold213/X _4354_/S vssd1 vssd1 vccd1 vccd1 _6014_/D sky130_fd_sc_hd__mux2_1
XANTENNA__5814__B2 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6019_ _6035_/CLK _6019_/D vssd1 vssd1 vccd1 vccd1 _6019_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5042__A2 _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4896__A _6236_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5491__S _5497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4164__S0 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4835__S _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3816__B1 _6138_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3292__A1 _3488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4467__S1 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3720_ _3573_/C _3986_/A2 _3584_/X _3585_/X _6005_/Q vssd1 vssd1 vccd1 vccd1 _3720_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3694__B _4735_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3651_ _6073_/Q _6072_/Q _3652_/B vssd1 vssd1 vccd1 vccd1 _5033_/A sky130_fd_sc_hd__nand3_2
XANTENNA__5741__B1 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4544__A1 _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3582_ _3573_/C _3577_/S _3580_/X _3581_/X vssd1 vssd1 vccd1 vccd1 _3582_/Y sky130_fd_sc_hd__o31ai_4
XANTENNA__3978__S0 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5321_ _6164_/Q _5320_/S _5317_/Y _3461_/A vssd1 vssd1 vccd1 vccd1 _5321_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_23_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5252_ _5289_/S _5252_/B vssd1 vssd1 vccd1 vccd1 _5252_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5183_ _4255_/S _5181_/X _5182_/X _5200_/A2 vssd1 vssd1 vccd1 vccd1 _5183_/X sky130_fd_sc_hd__o22a_1
X_4203_ _4205_/B vssd1 vssd1 vccd1 vccd1 _4203_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4134_ _3974_/B _4134_/B vssd1 vssd1 vccd1 vccd1 _4135_/D sky130_fd_sc_hd__and2b_1
XANTENNA__3215__A _5838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4065_ _4398_/B _3301_/B _3298_/A vssd1 vssd1 vccd1 vccd1 _4065_/X sky130_fd_sc_hd__o21a_1
X_3016_ _3507_/C _3137_/A vssd1 vssd1 vccd1 vccd1 _3484_/A sky130_fd_sc_hd__nor2_1
XANTENNA__3588__C _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4967_ _6158_/Q _5013_/S vssd1 vssd1 vccd1 vccd1 _4967_/X sky130_fd_sc_hd__or2_1
XANTENNA__4480__S _4596_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4898_ _6196_/Q _6062_/Q _6038_/Q vssd1 vssd1 vccd1 vccd1 _4898_/X sky130_fd_sc_hd__mux2_1
X_3918_ _6140_/Q _3648_/A _3650_/X _5386_/B vssd1 vssd1 vccd1 vccd1 _3918_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4783__A1 _6188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3849_ _5333_/B _3849_/B vssd1 vssd1 vccd1 vccd1 _3851_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_34_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3109__B _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5519_ _5518_/X _5514_/A _5566_/S vssd1 vssd1 vccd1 vccd1 _5519_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_42_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3743__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6251__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout120 _3193_/A vssd1 vssd1 vccd1 vccd1 _3643_/A sky130_fd_sc_hd__buf_4
Xfanout131 _6254_/Q vssd1 vssd1 vccd1 vccd1 _4485_/A sky130_fd_sc_hd__clkbuf_8
Xfanout142 hold652/X vssd1 vssd1 vccd1 vccd1 _4077_/A sky130_fd_sc_hd__buf_4
XANTENNA__3125__A _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout164 _3539_/A vssd1 vssd1 vccd1 vccd1 _4460_/A sky130_fd_sc_hd__buf_6
Xfanout153 hold648/X vssd1 vssd1 vccd1 vccd1 _5076_/A0 sky130_fd_sc_hd__buf_6
Xfanout175 fanout176/X vssd1 vssd1 vccd1 vccd1 fanout175/X sky130_fd_sc_hd__buf_4
XANTENNA__5340__A _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold632_A _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5015__A2 _4766_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5250__A _5250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5903__RESET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5870_ _4030_/Y _5834_/X _5837_/X _5869_/X vssd1 vssd1 vccd1 vccd1 _5870_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_87_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4821_ _4990_/A _4821_/B vssd1 vssd1 vccd1 vccd1 _4821_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4752_ _5245_/A hold628/X _4927_/S _4751_/X vssd1 vssd1 vccd1 vccd1 _6074_/D sky130_fd_sc_hd__a22o_1
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3568__A2 _5313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4683_ hold72/A _5933_/Q _5925_/Q _6033_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4683_/X sky130_fd_sc_hd__mux4_1
X_3703_ _5033_/A _5383_/B _5374_/B _3624_/Y vssd1 vssd1 vccd1 vccd1 _3704_/B sky130_fd_sc_hd__a2bb2o_1
XANTENNA__5714__B1 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4517__B2 _4474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3634_ _5333_/B _3633_/X _3634_/S vssd1 vssd1 vccd1 vccd1 _3636_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5190__A1 _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3565_ _3711_/B _3564_/Y _3554_/X _4618_/B vssd1 vssd1 vccd1 vccd1 _3565_/X sky130_fd_sc_hd__o211a_1
X_3496_ _5502_/A _3713_/B _3496_/C vssd1 vssd1 vccd1 vccd1 _3496_/X sky130_fd_sc_hd__or3_4
X_5304_ hold179/X _3979_/X _5305_/S vssd1 vssd1 vccd1 vccd1 _5304_/X sky130_fd_sc_hd__mux2_1
X_5235_ _4077_/A _5222_/C hold517/X _5218_/X hold50/X vssd1 vssd1 vccd1 vccd1 _5235_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5166_ _6158_/Q _5121_/Y _5122_/Y _6192_/Q vssd1 vssd1 vccd1 vccd1 _5176_/B sky130_fd_sc_hd__a22o_1
X_5097_ _4038_/A _4726_/A _3277_/A _3203_/B _5096_/X vssd1 vssd1 vccd1 vccd1 _5097_/X
+ sky130_fd_sc_hd__a221o_1
X_4117_ _4118_/A _4117_/B _4117_/C vssd1 vssd1 vccd1 vccd1 _5007_/A sky130_fd_sc_hd__and3_2
XANTENNA__3599__B _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3256__A1 _3302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4048_ _4048_/A _4048_/B _4418_/C _4045_/X vssd1 vssd1 vccd1 vccd1 _4048_/X sky130_fd_sc_hd__or4b_1
XANTENNA__4453__B1 _3434_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5999_ _6149_/CLK _5999_/D vssd1 vssd1 vccd1 vccd1 _5999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4756__A1 _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2959__A _6172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3495__A1 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold409 _5215_/X vssd1 vssd1 vccd1 vccd1 _6120_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5245__A _5245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3350_ _5314_/A _5566_/S _3503_/C vssd1 vssd1 vccd1 vccd1 _3353_/B sky130_fd_sc_hd__or3_4
XANTENNA__3722__A2 _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ hold319/X _5019_/X _5020_/S vssd1 vssd1 vccd1 vccd1 _5020_/X sky130_fd_sc_hd__mux2_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _3281_/A _3281_/B _3281_/C vssd1 vssd1 vccd1 vccd1 _3290_/B sky130_fd_sc_hd__or3_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4295__S _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5922_ _6030_/CLK _5922_/D vssd1 vssd1 vccd1 vccd1 _5922_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__3789__A2 _3745_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5853_ _6116_/Q _5852_/X _5869_/S vssd1 vssd1 vccd1 vccd1 _5853_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_61_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5784_ _6174_/Q hold429/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5784_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_63_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4804_ hold341/X _4803_/X _4927_/S vssd1 vssd1 vccd1 vccd1 _4804_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2996_ _2996_/A vssd1 vssd1 vccd1 vccd1 _5590_/A sky130_fd_sc_hd__inv_2
XFILLER_0_56_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4735_ _4735_/A _4759_/A vssd1 vssd1 vccd1 vccd1 _4735_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3410__A1 _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4043__B _5502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4666_ _4522_/B _4619_/X _4665_/Y vssd1 vssd1 vccd1 vccd1 _4666_/Y sky130_fd_sc_hd__a21oi_1
X_4597_ _4595_/X _4596_/X _5762_/A vssd1 vssd1 vccd1 vccd1 _4597_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_12_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3617_ hold86/X hold84/X _3724_/S vssd1 vssd1 vccd1 vccd1 _3617_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4910__A1 _4909_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3548_ _4061_/A _3709_/B vssd1 vssd1 vccd1 vccd1 _3548_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_101_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3479_ _3479_/A _3479_/B _4427_/A vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__or3_1
X_6198_ _6203_/CLK _6198_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6198_/Q sky130_fd_sc_hd__dfrtp_4
X_5218_ _5220_/A _5218_/B vssd1 vssd1 vccd1 vccd1 _5218_/X sky130_fd_sc_hd__and2_2
X_5149_ _6238_/Q _5108_/Y _5129_/Y _6214_/Q _5148_/X vssd1 vssd1 vccd1 vccd1 _5150_/C
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5602__B _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3229__A1 _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3403__A _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5769__A3 _5711_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3122__B _4725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4234__A _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3401__A1 _6127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4074__D_N _5250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5154__B2 _6199_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4520_ _6156_/Q _4519_/X _4598_/S vssd1 vssd1 vccd1 vccd1 _4520_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5145__A1 _5116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold206 _6032_/Q vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_25_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold217 _5980_/Q vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
X_4451_ _3405_/B _4438_/X _4451_/C _5917_/Q vssd1 vssd1 vccd1 vccd1 _4451_/X sky130_fd_sc_hd__and4bb_1
Xhold228 _6025_/Q vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold239 _5928_/Q vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__dlygate4sd3_1
X_3402_ hold57/X _3402_/B _5979_/D hold41/X vssd1 vssd1 vccd1 vccd1 _6077_/D sky130_fd_sc_hd__or4_1
X_6121_ _6243_/CLK _6121_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6121_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__3207__B _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4382_ _4451_/C _4391_/B _4038_/A vssd1 vssd1 vccd1 vccd1 _4385_/B sky130_fd_sc_hd__a21oi_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _3333_/A _3333_/B vssd1 vssd1 vccd1 vccd1 _3334_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ _6190_/CLK _6052_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6052_/Q sky130_fd_sc_hd__dfrtp_1
X_3264_ _5838_/B _3264_/B vssd1 vssd1 vccd1 vccd1 _3264_/X sky130_fd_sc_hd__or2_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3459__A1 hold567/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5003_ _5007_/A _5002_/Y _4990_/Y vssd1 vssd1 vccd1 vccd1 _5003_/X sky130_fd_sc_hd__o21a_1
XANTENNA__6208__SET_B fanout177/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _4486_/A _4056_/B vssd1 vssd1 vccd1 vccd1 _5093_/A sky130_fd_sc_hd__or2_2
XANTENNA__5849__S _5869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5081__B1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5905_ _6144_/CLK _5905_/D vssd1 vssd1 vccd1 vccd1 _5905_/Q sky130_fd_sc_hd__dfxtp_1
X_5836_ _5836_/A vssd1 vssd1 vccd1 vccd1 _5836_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_48_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6095__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5767_ _5767_/A _5767_/B vssd1 vssd1 vccd1 vccd1 _5767_/Y sky130_fd_sc_hd__nand2_1
X_2979_ _2979_/A vssd1 vssd1 vccd1 vccd1 _3849_/B sky130_fd_sc_hd__inv_2
XANTENNA__3893__A _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5698_ _5698_/A _5698_/B vssd1 vssd1 vccd1 vccd1 _5698_/Y sky130_fd_sc_hd__xnor2_1
X_4718_ _4718_/A _4718_/B vssd1 vssd1 vccd1 vccd1 _4718_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4649_ hold520/X _4612_/B _4648_/Y _4474_/X vssd1 vssd1 vccd1 vccd1 _4649_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_97_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3698__A1 _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6035_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout79_A _3594_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5494__S _5497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4178__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5127__A1 _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5127__B2 _6188_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5507__B _5507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4886__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4838__S _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3310__B1 _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5669__S _5705_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_A _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4573__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3951_ _6140_/Q _5046_/A _5868_/S vssd1 vssd1 vccd1 vccd1 _5394_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3882_ _6150_/Q _3611_/X _3613_/X hold98/A vssd1 vssd1 vccd1 vccd1 _3888_/A sky130_fd_sc_hd__a22o_1
XFILLER_0_42_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5366__A1 _3707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5621_ _5620_/X _5613_/A _5705_/S vssd1 vssd1 vccd1 vccd1 _5621_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4169__A2 _3588_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5552_ _5552_/A _5552_/B _5552_/C vssd1 vssd1 vccd1 vccd1 _5559_/A sky130_fd_sc_hd__and3_1
XFILLER_0_5_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3377__B1 _4725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4503_ hold548/X input2/X _4596_/S vssd1 vssd1 vccd1 vccd1 _4503_/X sky130_fd_sc_hd__mux2_1
X_5483_ _6235_/Q _6179_/Q _5773_/B vssd1 vssd1 vccd1 vccd1 _5483_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4434_ _3715_/B _3713_/A _4445_/B _4043_/C _4739_/B vssd1 vssd1 vccd1 vccd1 _4435_/B
+ sky130_fd_sc_hd__o221a_1
X_4365_ hold122/X _4150_/X _4372_/S vssd1 vssd1 vccd1 vccd1 _4365_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_6104_ _6208_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ _3290_/B _3334_/A _3314_/X _3315_/X _3498_/A vssd1 vssd1 vccd1 vccd1 _3316_/X
+ sky130_fd_sc_hd__o41a_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ _6035_/CLK _6035_/D vssd1 vssd1 vccd1 vccd1 _6035_/Q sky130_fd_sc_hd__dfxtp_1
X_4296_ _3836_/X hold139/X _4300_/S vssd1 vssd1 vccd1 vccd1 _4296_/X sky130_fd_sc_hd__mux2_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _3715_/B _5093_/B vssd1 vssd1 vccd1 vccd1 _3247_/Y sky130_fd_sc_hd__nand2_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4991__B _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3178_ _3203_/A _3178_/B _3178_/C vssd1 vssd1 vccd1 vccd1 _3477_/B sky130_fd_sc_hd__and3_2
XFILLER_0_95_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5579__S _5705_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5819_ _6241_/Q _5791_/X _5818_/X _5764_/B vssd1 vssd1 vccd1 vccd1 _5819_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3907__A2 _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4512__A _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5109__A1 _5120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4580__A2 _4612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4868__A0 _4865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold570 _5733_/X vssd1 vssd1 vccd1 vccd1 _6209_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 _3390_/X vssd1 vssd1 vccd1 vccd1 hold581/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 _6124_/Q vssd1 vssd1 vccd1 vccd1 hold592/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4096__A1 _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3798__A _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5596__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4406__B _4446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4568__S _4598_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4150_ _4242_/S _4133_/X _4148_/Y _4149_/X vssd1 vssd1 vccd1 vccd1 _4150_/X sky130_fd_sc_hd__a22o_2
X_3101_ _3113_/B _3203_/D vssd1 vssd1 vccd1 vccd1 _3101_/Y sky130_fd_sc_hd__nor2_1
X_4081_ _4398_/B _4726_/A _4618_/C _3228_/B vssd1 vssd1 vccd1 vccd1 _4084_/B sky130_fd_sc_hd__a22o_1
X_3032_ _6259_/Q _6258_/Q _3193_/A vssd1 vssd1 vccd1 vccd1 _3249_/B sky130_fd_sc_hd__or3b_4
X_4983_ _4999_/A1 _4980_/X _4982_/X _4824_/B vssd1 vssd1 vccd1 vccd1 _4983_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_58_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3934_ _6141_/Q _3934_/B vssd1 vssd1 vccd1 vccd1 _3935_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3865_ _3597_/X _3864_/A _3539_/Y vssd1 vssd1 vccd1 vccd1 _3865_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_73_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5604_ _5604_/A _5604_/B _5602_/Y vssd1 vssd1 vccd1 vccd1 _5605_/B sky130_fd_sc_hd__or3b_1
X_3796_ _5895_/Q _3588_/X _3793_/X _3794_/X _3795_/X vssd1 vssd1 vccd1 vccd1 _3798_/D
+ sky130_fd_sc_hd__a2111o_1
X_5535_ _6156_/Q _5507_/Y _5508_/X vssd1 vssd1 vccd1 vccd1 _5538_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5466_ hold576/X _5465_/X _5488_/S vssd1 vssd1 vccd1 vccd1 _5466_/X sky130_fd_sc_hd__mux2_1
X_4417_ _4417_/A _4417_/B _4759_/A vssd1 vssd1 vccd1 vccd1 _4417_/X sky130_fd_sc_hd__or3_1
X_5397_ _5397_/A _5397_/B vssd1 vssd1 vccd1 vccd1 _5398_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4348_ _4165_/X hold277/X _4354_/S vssd1 vssd1 vccd1 vccd1 _6013_/D sky130_fd_sc_hd__mux2_1
X_4279_ hold70/X _4211_/X _4282_/S vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__mux2_1
XANTENNA__4078__A1 _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6018_ _6032_/CLK _6018_/D vssd1 vssd1 vccd1 vccd1 _6018_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold410_A _6116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold508_A _6135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5772__S _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5750__A1 _3785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_33_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6251_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4896__B _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6198__RESET_B fanout184/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3816__A1 _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4164__S1 _5200_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6127__RESET_B fanout171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3321__A _5424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3292__A2 _3543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3650_ _6073_/Q _6072_/Q _3652_/B vssd1 vssd1 vccd1 vccd1 _3650_/X sky130_fd_sc_hd__and3_2
XFILLER_0_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3694__C _3694_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3581_ _3513_/A _3571_/X _3559_/A _4963_/A vssd1 vssd1 vccd1 vccd1 _3581_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3978__S1 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5320_ _5319_/X _3461_/A _5320_/S vssd1 vssd1 vccd1 vccd1 _5320_/X sky130_fd_sc_hd__mux2_1
X_5251_ _5259_/B _5252_/B vssd1 vssd1 vccd1 vccd1 _5251_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__4298__S _4300_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4202_ _4202_/A _4202_/B vssd1 vssd1 vccd1 vccd1 _4205_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_11_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5182_ _6017_/Q _5925_/Q _5182_/S vssd1 vssd1 vccd1 vccd1 _5182_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4133_ hold145/X hold151/X hold239/X hold169/X _5200_/B1 _5182_/S vssd1 vssd1 vccd1
+ vccd1 _4133_/X sky130_fd_sc_hd__mux4_1
XANTENNA__3215__B _4759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3930__S _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4064_ _4045_/X _4063_/Y _3694_/C vssd1 vssd1 vccd1 vccd1 _4069_/A sky130_fd_sc_hd__a21oi_1
X_3015_ _4038_/B _4043_/A vssd1 vssd1 vccd1 vccd1 _3137_/A sky130_fd_sc_hd__nand2_2
XANTENNA__5009__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4480__A1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5857__S _5869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4966_ _6066_/Q _4966_/B vssd1 vssd1 vccd1 vccd1 _4966_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4897_ _6212_/Q _5009_/A2 _4769_/Y _4895_/B _4896_/X vssd1 vssd1 vccd1 vccd1 _4897_/X
+ sky130_fd_sc_hd__a221o_1
X_3917_ _5386_/B vssd1 vssd1 vccd1 vccd1 _5032_/B sky130_fd_sc_hd__inv_2
XFILLER_0_61_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3440__C1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3848_ _6139_/Q _3848_/B _3851_/B vssd1 vssd1 vccd1 vccd1 _3859_/A sky130_fd_sc_hd__or3b_1
XANTENNA__5732__A1 _3926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3779_ _3646_/X _3778_/B _3778_/Y _3645_/X vssd1 vssd1 vccd1 vccd1 _3779_/X sky130_fd_sc_hd__a211o_1
XANTENNA__3743__B1 _3739_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5518_ _5517_/X hold527/X _5609_/S vssd1 vssd1 vccd1 vccd1 _5518_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5496__A0 _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5449_ _6072_/Q _3652_/B _5448_/A _5333_/Y _5448_/Y vssd1 vssd1 vccd1 vccd1 _5449_/X
+ sky130_fd_sc_hd__a221o_1
Xfanout121 _4061_/A vssd1 vssd1 vccd1 vccd1 _3193_/A sky130_fd_sc_hd__buf_2
Xfanout110 _5772_/S vssd1 vssd1 vccd1 vccd1 _5875_/A sky130_fd_sc_hd__clkbuf_8
Xfanout132 hold638/X vssd1 vssd1 vccd1 vccd1 _4094_/D sky130_fd_sc_hd__clkbuf_4
Xfanout143 _4451_/C vssd1 vssd1 vccd1 vccd1 _4765_/A sky130_fd_sc_hd__clkbuf_8
Xfanout165 _3539_/A vssd1 vssd1 vccd1 vccd1 _4485_/B sky130_fd_sc_hd__clkbuf_8
Xfanout154 hold609/X vssd1 vssd1 vccd1 vccd1 _5333_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__5248__B1 _4409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout176 input13/X vssd1 vssd1 vccd1 vccd1 fanout176/X sky130_fd_sc_hd__buf_4
XANTENNA__5799__B2 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5799__A1 _6237_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5340__B wire93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout61_A _4763_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3795__B _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5723__A1 _3785_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3734__B1 _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5487__A0 _4030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3501__A3 _6094_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5239__B1 _5120_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5250__B _5250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4462__A1 _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4581__S _4596_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4820_ hold309/X _4819_/X _4927_/S vssd1 vssd1 vccd1 vccd1 _4820_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4751_ _4618_/B _4749_/X _4750_/X _4118_/A _4415_/X vssd1 vssd1 vccd1 vccd1 _4751_/X
+ sky130_fd_sc_hd__a221o_1
X_4682_ hold501/X _4681_/Y _5073_/S vssd1 vssd1 vccd1 vccd1 _4682_/X sky130_fd_sc_hd__mux2_1
X_3702_ _3912_/B _3820_/A _6136_/Q vssd1 vssd1 vccd1 vccd1 _5383_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_7_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5714__A1 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4517__A2 _4612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3633_ _6070_/Q _5333_/B vssd1 vssd1 vccd1 vccd1 _3633_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_3_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3564_ _3562_/Y _3563_/Y _3090_/Y vssd1 vssd1 vccd1 vccd1 _3564_/Y sky130_fd_sc_hd__a21oi_1
X_5303_ hold216/X _3930_/X _5305_/S vssd1 vssd1 vccd1 vccd1 _6150_/D sky130_fd_sc_hd__mux2_1
X_3495_ _3715_/B _3494_/X _3462_/Y vssd1 vssd1 vccd1 vccd1 _5954_/D sky130_fd_sc_hd__o21ai_1
X_5234_ hold50/X _3353_/B _5217_/A hold497/X vssd1 vssd1 vccd1 vccd1 _5234_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3226__A _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5165_ _6208_/Q _5106_/Y _5108_/Y _6240_/Q vssd1 vssd1 vccd1 vccd1 _5176_/A sky130_fd_sc_hd__a22o_1
XANTENNA__6049__RESET_B fanout176/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4116_ _4460_/A _4116_/B vssd1 vssd1 vccd1 vccd1 _4116_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5096_ _3545_/A _4044_/B _4383_/Y _3488_/B _5095_/X vssd1 vssd1 vccd1 vccd1 _5096_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3599__C _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4453__A1 _3405_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4047_ _4439_/B _4053_/A _4046_/Y vssd1 vssd1 vccd1 vccd1 _4418_/C sky130_fd_sc_hd__a21o_1
XANTENNA__4453__B2 _4750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5587__S _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5998_ _6006_/CLK _5998_/D vssd1 vssd1 vccd1 vccd1 _5998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4949_ _6064_/Q _4948_/C _6065_/Q vssd1 vssd1 vccd1 vccd1 _4950_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3136__A _4726_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2975__A _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5351__A _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4444__A1 _4433_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5497__S _5497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3280_ _5502_/B _3477_/C _4424_/D _4483_/B vssd1 vssd1 vccd1 vccd1 _3281_/C sky130_fd_sc_hd__or4_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5921_ _6029_/CLK _5921_/D vssd1 vssd1 vccd1 vccd1 _5921_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4986__A2 _5702_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5852_ _6120_/Q _6138_/Q _5868_/S vssd1 vssd1 vccd1 vccd1 _5852_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_48_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5783_ _6173_/Q hold478/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5783_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4199__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4803_ _4802_/X _6055_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _4803_/X sky130_fd_sc_hd__mux2_1
X_2995_ _6193_/Q vssd1 vssd1 vccd1 vccd1 _5582_/A sky130_fd_sc_hd__inv_2
XFILLER_0_8_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4734_ _3556_/A _4749_/C _4733_/X vssd1 vssd1 vccd1 vccd1 _4738_/B sky130_fd_sc_hd__o21a_1
XANTENNA__4043__C _4043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4665_ _5764_/B _4663_/X _4664_/X vssd1 vssd1 vccd1 vccd1 _4665_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4596_ hold534/X input8/X _4596_/S vssd1 vssd1 vccd1 vccd1 _4596_/X sky130_fd_sc_hd__mux2_1
X_3616_ _3988_/A _3616_/B _3793_/D vssd1 vssd1 vccd1 vccd1 _4364_/A sky130_fd_sc_hd__or3_4
XANTENNA_fanout111_A _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3547_ _5093_/A _3246_/A _3246_/B _3543_/Y _3546_/X vssd1 vssd1 vccd1 vccd1 _3547_/X
+ sky130_fd_sc_hd__o311a_1
X_3478_ _3478_/A _4772_/D vssd1 vssd1 vccd1 vccd1 _4759_/C sky130_fd_sc_hd__nor2_1
XANTENNA__4123__A0 _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6197_ _6238_/CLK _6197_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6197_/Q sky130_fd_sc_hd__dfrtp_4
X_5217_ _5217_/A vssd1 vssd1 vccd1 vccd1 _5217_/Y sky130_fd_sc_hd__inv_2
XANTENNA__3106__D _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5148_ _6198_/Q _5119_/Y _5146_/X _5109_/Y vssd1 vssd1 vccd1 vccd1 _5148_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3403__B _5424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5079_ _3477_/B _4406_/Y _5078_/X vssd1 vssd1 vccd1 vccd1 _5080_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__3229__A2 _4451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4665__A1 _5764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3468__A2 _3713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5090__A1 _4451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5020__S _5020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold207 _4369_/X vssd1 vssd1 vccd1 vccd1 _6032_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4450_ _4118_/A _4449_/X _4448_/X _4443_/Y vssd1 vssd1 vccd1 vccd1 _4450_/X sky130_fd_sc_hd__a211o_1
Xhold229 _4361_/X vssd1 vssd1 vccd1 vccd1 _6025_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_200 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3401_ _6127_/Q _2964_/Y _3366_/X _3353_/X hold40/X vssd1 vssd1 vccd1 vccd1 hold41/A
+ sky130_fd_sc_hd__a32o_1
X_4381_ _4417_/A _4381_/B vssd1 vssd1 vccd1 vccd1 _4381_/Y sky130_fd_sc_hd__nor2_1
Xhold218 _4311_/X vssd1 vssd1 vccd1 vccd1 _5980_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6120_ _6178_/CLK _6120_/D vssd1 vssd1 vccd1 vccd1 _6120_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_0_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3332_ _3324_/A _3324_/B _3283_/A vssd1 vssd1 vccd1 vccd1 _3333_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_21_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5853__A0 _6116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6051_ _6144_/CLK _6051_/D fanout172/X vssd1 vssd1 vccd1 vccd1 _6051_/Q sky130_fd_sc_hd__dfrtp_1
X_3263_ _4446_/A _4044_/B _5424_/A vssd1 vssd1 vccd1 vccd1 _3264_/B sky130_fd_sc_hd__a21oi_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _6068_/Q _5702_/A2 _5607_/B1 _5001_/X vssd1 vssd1 vccd1 vccd1 _5002_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_0_56_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3194_ _4486_/A _4056_/B vssd1 vssd1 vccd1 vccd1 _3196_/B sky130_fd_sc_hd__nor2_2
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4038__C _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4408__A1 _4391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5081__A1 _3302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5904_ _6144_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
X_5835_ _5837_/A _5834_/X _5773_/A vssd1 vssd1 vccd1 vccd1 _5836_/A sky130_fd_sc_hd__a21oi_4
XANTENNA_fanout159_A _5164_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5865__S _5869_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5766_ _5765_/X _5763_/X _5771_/S _3959_/A vssd1 vssd1 vccd1 vccd1 _5766_/X sky130_fd_sc_hd__o2bb2a_1
X_2978_ _2978_/A vssd1 vssd1 vccd1 vccd1 _3805_/B sky130_fd_sc_hd__inv_2
XFILLER_0_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5697_ _5707_/S _5696_/X _5624_/X _5685_/A vssd1 vssd1 vccd1 vccd1 _5697_/X sky130_fd_sc_hd__o2bb2a_1
X_4717_ _4716_/A _4716_/B _4716_/C vssd1 vssd1 vccd1 vccd1 _4718_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4648_ _4648_/A _4648_/B vssd1 vssd1 vccd1 vccd1 _4648_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__5136__A2 _5105_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4070__A _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3147__A1 _4391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3698__A2 _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4579_ _4579_/A _4579_/B vssd1 vssd1 vccd1 vccd1 _4579_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5613__B _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6249_ _6251_/CLK _6249_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6249_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5844__A0 _6114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4583__A0 _6160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4886__B2 _4879_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5835__B1 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3310__A1 _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3950_ _4036_/B _3950_/B vssd1 vssd1 vccd1 vccd1 _3950_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_58_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3881_ hold155/X _3880_/X _4035_/S vssd1 vssd1 vccd1 vccd1 _3881_/X sky130_fd_sc_hd__mux2_1
X_5620_ _5619_/X _6154_/Q _5704_/S vssd1 vssd1 vccd1 vccd1 _5620_/X sky130_fd_sc_hd__mux2_1
X_5551_ _5551_/A _5551_/B vssd1 vssd1 vccd1 vccd1 _5552_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__3377__A1 _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4502_ hold548/X _4612_/B _4501_/X _4474_/X vssd1 vssd1 vccd1 vccd1 _4502_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5482_ _5025_/A _5479_/X _5481_/X _4019_/X vssd1 vssd1 vccd1 vccd1 _5482_/X sky130_fd_sc_hd__a211o_1
XFILLER_0_13_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4433_ _4433_/A _4433_/B _5838_/B _4749_/A vssd1 vssd1 vccd1 vccd1 _4739_/B sky130_fd_sc_hd__or4_1
XFILLER_0_67_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4364_ _4364_/A _4364_/B vssd1 vssd1 vccd1 vccd1 _4372_/S sky130_fd_sc_hd__nor2_4
X_6103_ _6148_/CLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
X_4295_ _3789_/X hold259/X _4300_/S vssd1 vssd1 vccd1 vccd1 _5959_/D sky130_fd_sc_hd__mux2_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _4618_/C _3285_/Y _3288_/B _3395_/B vssd1 vssd1 vccd1 vccd1 _3315_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ _6034_/CLK _6034_/D vssd1 vssd1 vccd1 vccd1 _6034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _3246_/A _3246_/B vssd1 vssd1 vccd1 vccd1 _3542_/B sky130_fd_sc_hd__or2_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3177_ _3177_/A _3281_/A _3177_/C vssd1 vssd1 vccd1 vccd1 _3177_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5818_ hold476/X _5457_/A _5352_/Y _2990_/Y vssd1 vssd1 vccd1 vccd1 _5818_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5749_ _4119_/A _4928_/B _4648_/Y _5762_/C vssd1 vssd1 vccd1 vccd1 _5749_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6245__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5109__A2 _5107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5046__D _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold571 _6215_/Q vssd1 vssd1 vccd1 vccd1 hold571/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold560 _4569_/X vssd1 vssd1 vccd1 vccd1 _6059_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold593 _6238_/Q vssd1 vssd1 vccd1 vccd1 hold593/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold582 _3391_/X vssd1 vssd1 vccd1 vccd1 _5916_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3144__A _3694_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5293__A1 _5245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2983__A _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3753__S _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4849__S _4927_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3100_ _3203_/D vssd1 vssd1 vccd1 vccd1 _3178_/C sky130_fd_sc_hd__inv_2
X_4080_ _4043_/A _4750_/A _4416_/C _4079_/X vssd1 vssd1 vccd1 vccd1 _4084_/A sky130_fd_sc_hd__a211o_1
XFILLER_0_37_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4584__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3031_ _3249_/A _3070_/A vssd1 vssd1 vccd1 vccd1 _4398_/C sky130_fd_sc_hd__or2_1
XANTENNA__3834__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4492__C1 _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4982_ _6159_/Q _4981_/X _5013_/S vssd1 vssd1 vccd1 vccd1 _4982_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3933_ _6141_/Q _3934_/B vssd1 vssd1 vccd1 vccd1 _3939_/B sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_3_wb_clk_i _5978_/CLK vssd1 vssd1 vccd1 vccd1 _6152_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3864_ _3864_/A vssd1 vssd1 vccd1 vccd1 _3864_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_46_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5603_ _5604_/A _5604_/B _5602_/Y vssd1 vssd1 vccd1 vccd1 _5603_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3795_ _6007_/Q _3968_/A _3795_/C _3885_/S vssd1 vssd1 vccd1 vccd1 _3795_/X sky130_fd_sc_hd__and4_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5534_ hold512/X _5533_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _5534_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5465_ _3926_/X _5464_/X _5487_/S vssd1 vssd1 vccd1 vccd1 _5465_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4416_ _4416_/A _4416_/B _4416_/C vssd1 vssd1 vccd1 vccd1 _4750_/C sky130_fd_sc_hd__or3_1
X_5396_ _5396_/A _5396_/B vssd1 vssd1 vccd1 vccd1 _5398_/A sky130_fd_sc_hd__xor2_1
XANTENNA__3522__A1 _5317_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4347_ _4150_/X hold267/X _4354_/S vssd1 vssd1 vccd1 vccd1 _6012_/D sky130_fd_sc_hd__mux2_1
X_4278_ hold82/X _4193_/X _4282_/S vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__mux2_1
XANTENNA__5275__A1 _6158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6017_ _6033_/CLK _6017_/D vssd1 vssd1 vccd1 vccd1 _6017_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__5275__B2 _6240_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3229_ _4398_/A _4451_/C _3227_/B _3224_/X _3228_/Y vssd1 vssd1 vccd1 vccd1 _3229_/X
+ sky130_fd_sc_hd__o311a_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4507__B _4507_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5027__A1 _2960_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5750__A2 _5771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5354__A _5705_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold390 _6062_/Q vssd1 vssd1 vccd1 vccd1 hold390/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3602__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3816__A2 _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5018__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4624__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5741__A2 _5771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3580_ hold23/A _4253_/A2 _4034_/S vssd1 vssd1 vccd1 vccd1 _3580_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_51_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5250_ _5250_/A _5250_/B _4409_/X vssd1 vssd1 vccd1 vccd1 _5252_/B sky130_fd_sc_hd__or3b_1
X_4201_ hold265/X _3605_/X _3615_/X hold206/X _4200_/X vssd1 vssd1 vccd1 vccd1 _4202_/B
+ sky130_fd_sc_hd__a221o_1
X_5181_ _5950_/Q _6033_/Q _5182_/S vssd1 vssd1 vccd1 vccd1 _5181_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3395__A_N _6048_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4132_ _4132_/A _4364_/B vssd1 vssd1 vccd1 vccd1 _4262_/S sky130_fd_sc_hd__nor2_4
X_4063_ _4735_/A _4124_/A _4046_/Y vssd1 vssd1 vccd1 vccd1 _4063_/Y sky130_fd_sc_hd__o21ai_1
X_3014_ _5356_/A _3694_/C vssd1 vssd1 vccd1 vccd1 _3777_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_93_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4965_ _6066_/Q _4966_/B vssd1 vssd1 vccd1 vccd1 _4995_/C sky130_fd_sc_hd__and2_1
XFILLER_0_80_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout141_A _6131_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3916_ _4005_/A _3916_/B vssd1 vssd1 vccd1 vccd1 _5386_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4896_ _6236_/Q _5008_/B vssd1 vssd1 vccd1 vccd1 _4896_/X sky130_fd_sc_hd__and2_1
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3847_ _5024_/A _6117_/Q vssd1 vssd1 vccd1 vccd1 _3851_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3991__A1 _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5732__A2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3778_ _3950_/B _3778_/B vssd1 vssd1 vccd1 vccd1 _3778_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5517_ _4119_/B _5516_/X _4757_/Y vssd1 vssd1 vccd1 vccd1 _5517_/X sky130_fd_sc_hd__a21bo_1
X_5448_ _5448_/A _5448_/B vssd1 vssd1 vccd1 vccd1 _5448_/Y sky130_fd_sc_hd__nor2_1
Xfanout100 _5341_/A vssd1 vssd1 vccd1 vccd1 _5764_/B sky130_fd_sc_hd__clkbuf_8
Xfanout111 _5772_/S vssd1 vssd1 vccd1 vccd1 _5073_/S sky130_fd_sc_hd__buf_6
X_5379_ _5378_/A _5378_/B _3848_/B vssd1 vssd1 vccd1 vccd1 _5379_/X sky130_fd_sc_hd__a21o_1
Xfanout122 hold580/X vssd1 vssd1 vccd1 vccd1 _4061_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout144 hold643/X vssd1 vssd1 vccd1 vccd1 _4451_/C sky130_fd_sc_hd__buf_4
Xfanout155 _5164_/A1 vssd1 vssd1 vccd1 vccd1 _3405_/B sky130_fd_sc_hd__buf_6
Xfanout133 _6253_/Q vssd1 vssd1 vccd1 vccd1 _3210_/A sky130_fd_sc_hd__buf_4
Xfanout177 fanout184/X vssd1 vssd1 vccd1 vccd1 fanout177/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__5248__A1 _5250_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout166 _3539_/A vssd1 vssd1 vccd1 vccd1 _4118_/A sky130_fd_sc_hd__buf_2
XANTENNA__3422__A _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4471__A2 _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout54_A _5705_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3795__C _3795_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5723__A2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3734__A1 _5249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5084__A _5085_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4998__A0 _6160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4750_ _4750_/A _4750_/B _4750_/C vssd1 vssd1 vccd1 vccd1 _4750_/X sky130_fd_sc_hd__or3_1
X_4681_ _4538_/B _4619_/X _4680_/Y vssd1 vssd1 vccd1 vccd1 _4681_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3701_ _6138_/Q _6176_/Q vssd1 vssd1 vccd1 vccd1 _3820_/A sky130_fd_sc_hd__or2_1
X_3632_ _6070_/Q _5333_/B vssd1 vssd1 vccd1 vccd1 _3647_/B sky130_fd_sc_hd__or2_1
XFILLER_0_70_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5302_ hold60/X _3880_/X _5305_/S vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__mux2_1
XFILLER_0_51_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3507__A _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3563_ _3563_/A _3713_/B vssd1 vssd1 vccd1 vccd1 _3563_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3494_ _3491_/B _3523_/B vssd1 vssd1 vccd1 vccd1 _3494_/X sky130_fd_sc_hd__and2b_1
X_5233_ _4077_/A _5222_/C _5219_/Y _5218_/X _6127_/Q vssd1 vssd1 vccd1 vccd1 _5233_/X
+ sky130_fd_sc_hd__a32o_1
XANTENNA__3226__B _4451_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5164_ _5164_/A1 _2978_/A _5086_/Y _5163_/X vssd1 vssd1 vccd1 vccd1 _5164_/X sky130_fd_sc_hd__a22o_1
X_4115_ hold58/X _4034_/X _4115_/S vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__mux2_1
X_5095_ _3446_/A _4391_/B _3477_/B _3543_/B vssd1 vssd1 vccd1 vccd1 _5095_/X sky130_fd_sc_hd__o211a_1
X_4046_ _4385_/A _4046_/B vssd1 vssd1 vccd1 vccd1 _4046_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_91_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5650__A1 _6199_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5868__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3256__A3 _5093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5997_ _6151_/CLK _5997_/D vssd1 vssd1 vccd1 vccd1 _5997_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4948_ _6064_/Q _6065_/Q _4948_/C vssd1 vssd1 vccd1 vccd1 _4966_/B sky130_fd_sc_hd__and3_1
XANTENNA__3413__B1 _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4879_ _4990_/A _4879_/B vssd1 vssd1 vccd1 vccd1 _4879_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4913__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4947__S _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5351__B _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4682__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4444__A2 _5838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2991__A _6189_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3327__A _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4380__A1 _4038_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3062__A _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5632__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5920_ _6149_/CLK _5920_/D vssd1 vssd1 vccd1 vccd1 _5920_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5851_ hold317/X _5836_/A _5850_/X _5773_/A vssd1 vssd1 vccd1 vccd1 _5851_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5782_ _6172_/Q hold456/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5782_/X sky130_fd_sc_hd__mux2_1
X_2994_ _6192_/Q vssd1 vssd1 vccd1 vccd1 _5569_/A sky130_fd_sc_hd__inv_2
XFILLER_0_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4802_ _4119_/B _4801_/X _4789_/Y vssd1 vssd1 vccd1 vccd1 _4802_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_61_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4733_ _4737_/A _4433_/B _4759_/A _3264_/B vssd1 vssd1 vccd1 vccd1 _4733_/X sky130_fd_sc_hd__a31o_1
XFILLER_0_16_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4664_ hold480/X _5762_/A _4619_/X vssd1 vssd1 vccd1 vccd1 _4664_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4595_ hold534/X _4612_/B _4594_/Y _4474_/X vssd1 vssd1 vccd1 vccd1 _4595_/X sky130_fd_sc_hd__a22o_1
X_3615_ _3968_/A _3983_/S _3982_/S vssd1 vssd1 vccd1 vccd1 _3615_/X sky130_fd_sc_hd__and3_4
XFILLER_0_43_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3546_ _4385_/A _3185_/C _4046_/B vssd1 vssd1 vccd1 vccd1 _3546_/X sky130_fd_sc_hd__a21o_1
XANTENNA_fanout104_A _5011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5216_ _5216_/A _5216_/B vssd1 vssd1 vccd1 vccd1 _5217_/A sky130_fd_sc_hd__and2_2
X_3477_ _3477_/A _3477_/B _3477_/C vssd1 vssd1 vccd1 vccd1 _4772_/D sky130_fd_sc_hd__or3_1
X_6196_ _6219_/CLK _6196_/D fanout178/X vssd1 vssd1 vccd1 vccd1 _6196_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA__5871__B2 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5147_ _6174_/Q _5104_/Y _5121_/Y _6156_/Q vssd1 vssd1 vccd1 vccd1 _5150_/B sky130_fd_sc_hd__a22o_1
XANTENNA__3882__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5078_ _5078_/A _5078_/B _5078_/C vssd1 vssd1 vccd1 vccd1 _5078_/X sky130_fd_sc_hd__or3_1
X_4029_ hold408/X _3958_/S _4028_/X vssd1 vssd1 vccd1 vccd1 _4030_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__5598__S _5705_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3700__A _6176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2986__A _6156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5311__A0 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5862__A1 _3926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5301__S _5305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4050__B1 _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold208 hold660/X vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold219 _6006_/Q vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_3400_ _5875_/A hold203/X _3397_/X _3399_/X vssd1 vssd1 vccd1 vccd1 _3400_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_0_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4380_ _4038_/A _4379_/X _3081_/B vssd1 vssd1 vccd1 vccd1 _4381_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3331_ _3396_/A _3545_/A _3286_/Y vssd1 vssd1 vccd1 vccd1 _3333_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3540_/A _3303_/A _3563_/A _3261_/X vssd1 vssd1 vccd1 vccd1 _3265_/B sky130_fd_sc_hd__a22o_1
X_6050_ _6123_/CLK _6050_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _6050_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ hold332/X _5000_/X _5701_/S vssd1 vssd1 vccd1 vccd1 _5001_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3504__B _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3193_ _3193_/A _4038_/A _3193_/C vssd1 vssd1 vccd1 vccd1 _3193_/X sky130_fd_sc_hd__and3_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3459__A3 _3713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5903_ _6130_/CLK _5903_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _5903_/Q sky130_fd_sc_hd__dfrtp_1
X_5834_ _6043_/Q _5834_/B _5834_/C _5834_/D vssd1 vssd1 vccd1 vccd1 _5834_/X sky130_fd_sc_hd__or4_4
XFILLER_0_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3919__A1 _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5765_ _5762_/A _4119_/A _4990_/B _5771_/S _5764_/X vssd1 vssd1 vccd1 vccd1 _5765_/X
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_56_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2977_ _2977_/A vssd1 vssd1 vccd1 vccd1 _3761_/B sky130_fd_sc_hd__inv_2
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5696_ _5004_/Y _5629_/Y _5695_/X _5691_/X _5511_/X vssd1 vssd1 vccd1 vccd1 _5696_/X
+ sky130_fd_sc_hd__a32o_1
X_4716_ _4716_/A _4716_/B _4716_/C vssd1 vssd1 vccd1 vccd1 _4718_/A sky130_fd_sc_hd__and3_1
X_4647_ _4647_/A _4647_/B _4647_/C vssd1 vssd1 vccd1 vccd1 _4648_/B sky130_fd_sc_hd__and3_1
XFILLER_0_71_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__4070__B _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4578_ _4561_/B _4563_/B _4561_/A vssd1 vssd1 vccd1 vccd1 _4579_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__4497__S _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3529_ _6070_/Q _5333_/B vssd1 vssd1 vccd1 vccd1 _3638_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6248_ _6251_/CLK _6248_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6248_/Q sky130_fd_sc_hd__dfrtp_1
X_6179_ _6235_/CLK _6179_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6179_/Q sky130_fd_sc_hd__dfstp_2
XFILLER_0_79_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6203_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5357__A _5484_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5780__A0 _6242_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5835__A1 _5837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3880_ _3878_/X _3879_/X _4034_/S vssd1 vssd1 vccd1 vccd1 _3880_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_45_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5771__A0 _4030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4574__A1 _4865_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5550_ _5551_/A _5551_/B vssd1 vssd1 vccd1 vccd1 _5571_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5481_ _6179_/Q _5026_/A _5480_/X _3920_/A _5330_/B vssd1 vssd1 vccd1 vccd1 _5481_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4501_ _4501_/A _4501_/B vssd1 vssd1 vccd1 vccd1 _4501_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_26_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4432_ _3210_/C _4056_/B _3306_/C _4445_/B vssd1 vssd1 vccd1 vccd1 _4738_/A sky130_fd_sc_hd__o211a_1
XANTENNA__3129__A2 _4398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4363_ _4261_/X hold214/X _4363_/S vssd1 vssd1 vccd1 vccd1 _4363_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4110__S _4115_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6102_ _6102_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfxtp_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ _4045_/A _3193_/X _4124_/A _3488_/B vssd1 vssd1 vccd1 vccd1 _3314_/X sky130_fd_sc_hd__a2bb2o_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4294_ _3737_/X hold321/X _4300_/S vssd1 vssd1 vccd1 vccd1 _4294_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5826__A1 _3959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6033_ _6033_/CLK _6033_/D vssd1 vssd1 vccd1 vccd1 _6033_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3643_/A _3237_/Y _3242_/X _3243_/X _4451_/C vssd1 vssd1 vccd1 vccd1 _3246_/B
+ sky130_fd_sc_hd__o2111a_2
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _4615_/B _4439_/A _3709_/B _3176_/D vssd1 vssd1 vccd1 vccd1 _3177_/C sky130_fd_sc_hd__or4_1
XANTENNA__3250__A _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout171_A fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5817_ hold594/X _5816_/X _5832_/S vssd1 vssd1 vccd1 vccd1 _6240_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_91_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5748_ hold538/X _5741_/Y _5747_/X _5767_/A vssd1 vssd1 vccd1 vccd1 _5748_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5679_ _5679_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5682_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_32_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold561 _6196_/Q vssd1 vssd1 vccd1 vccd1 _5613_/A sky130_fd_sc_hd__buf_1
Xhold572 _5754_/X vssd1 vssd1 vccd1 vccd1 _6215_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold550 _6210_/Q vssd1 vssd1 vccd1 vccd1 hold550/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold594 _6240_/Q vssd1 vssd1 vccd1 vccd1 hold594/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 _6211_/Q vssd1 vssd1 vccd1 vccd1 hold583/X sky130_fd_sc_hd__buf_1
XANTENNA_fanout84_A _3739_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5293__A2 _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold648_A _6112_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4253__B1 _3671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5087__A _5107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3819__B1 _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3030_ _3249_/A _3070_/A vssd1 vssd1 vccd1 vccd1 _3276_/A sky130_fd_sc_hd__nor2_2
X_4981_ _6067_/Q _4995_/C vssd1 vssd1 vccd1 vccd1 _4981_/X sky130_fd_sc_hd__xor2_1
XFILLER_0_58_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3932_ _6071_/Q _6119_/Q vssd1 vssd1 vccd1 vccd1 _3934_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_46_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3863_ _3862_/X _3849_/B _3958_/S vssd1 vssd1 vccd1 vccd1 _3864_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_73_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5602_ _5602_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5602_/Y sky130_fd_sc_hd__xnor2_1
X_3794_ _5960_/Q _3988_/A _3795_/C _3885_/S vssd1 vssd1 vccd1 vccd1 _3794_/X sky130_fd_sc_hd__and4_1
X_5533_ _5532_/X _5527_/Y _5670_/A vssd1 vssd1 vccd1 vccd1 _5533_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5464_ _3705_/A _5363_/C _5459_/X _5463_/X vssd1 vssd1 vccd1 vccd1 _5464_/X sky130_fd_sc_hd__a2bb2o_1
X_5395_ _5395_/A _5395_/B vssd1 vssd1 vccd1 vccd1 _5399_/A sky130_fd_sc_hd__xor2_1
X_4415_ _4415_/A _4415_/B vssd1 vssd1 vccd1 vccd1 _4415_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4346_ _4346_/A _4364_/B vssd1 vssd1 vccd1 vccd1 _4354_/S sky130_fd_sc_hd__or2_4
X_4277_ hold66/X _4180_/X _4282_/S vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__mux2_1
X_6016_ _6033_/CLK _6016_/D vssd1 vssd1 vccd1 vccd1 _6016_/Q sky130_fd_sc_hd__dfxtp_1
X_3228_ _3283_/A _3228_/B vssd1 vssd1 vccd1 vccd1 _3228_/Y sky130_fd_sc_hd__nand2_1
X_3159_ _3277_/A _3117_/X _3111_/X vssd1 vssd1 vccd1 vccd1 _3159_/X sky130_fd_sc_hd__a21o_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4786__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold598_A _6236_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold380 _6185_/Q vssd1 vssd1 vccd1 vccd1 hold380/X sky130_fd_sc_hd__buf_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold391 _4623_/X vssd1 vssd1 vccd1 vccd1 _6062_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4685__S _4697_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3602__B _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4417__C _4759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_42_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6170_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4433__B _4433_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3985__C1 _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4624__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3201__A1 _3715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4200_ _5924_/Q _3588_/X _3603_/X _6016_/Q vssd1 vssd1 vccd1 vccd1 _4200_/X sky130_fd_sc_hd__a22o_1
X_5180_ _3739_/S _5178_/X _5179_/X _3591_/A vssd1 vssd1 vccd1 vccd1 _5180_/X sky130_fd_sc_hd__o22a_1
X_4131_ _3671_/B _3539_/Y _3569_/Y _4130_/X _5023_/A vssd1 vssd1 vccd1 vccd1 _4364_/B
+ sky130_fd_sc_hd__a41o_4
XFILLER_0_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4062_ _3127_/B _4054_/X _4061_/X _3457_/A _3469_/Y vssd1 vssd1 vccd1 vccd1 _4062_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3512__B _5424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3013_ _4735_/A _4061_/A vssd1 vssd1 vccd1 vccd1 _4043_/A sky130_fd_sc_hd__nor2_1
X_4964_ _4104_/B _4962_/X _4963_/X _4999_/A1 vssd1 vssd1 vccd1 vccd1 _4964_/X sky130_fd_sc_hd__o211a_1
X_3915_ _3944_/A _4012_/A _6173_/Q vssd1 vssd1 vccd1 vccd1 _3916_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_46_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4895_ _4990_/A _4895_/B vssd1 vssd1 vccd1 vccd1 _4895_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3846_ _5033_/A _5386_/A _3845_/X vssd1 vssd1 vccd1 vccd1 _3846_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_46_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5193__A1 _6178_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3674__S _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3777_ _3777_/A _3777_/B vssd1 vssd1 vccd1 vccd1 _3778_/B sky130_fd_sc_hd__nor2_1
XANTENNA__3743__A2 _3591_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5516_ _6054_/Q _5595_/S _5607_/B1 _5515_/X vssd1 vssd1 vccd1 vccd1 _5516_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_42_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5447_ _5794_/B _5445_/Y _5446_/X _5365_/S vssd1 vssd1 vccd1 vccd1 _5447_/X sky130_fd_sc_hd__a31o_1
X_5378_ _5378_/A _5378_/B vssd1 vssd1 vccd1 vccd1 _5378_/Y sky130_fd_sc_hd__nor2_1
Xfanout112 _5772_/S vssd1 vssd1 vccd1 vccd1 _5488_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout101 _3378_/Y vssd1 vssd1 vccd1 vccd1 _5341_/A sky130_fd_sc_hd__clkbuf_8
Xfanout156 _5023_/A vssd1 vssd1 vccd1 vccd1 _5767_/A sky130_fd_sc_hd__clkbuf_8
Xfanout123 _4739_/A vssd1 vssd1 vccd1 vccd1 _5356_/A sky130_fd_sc_hd__buf_4
Xfanout145 _4038_/A vssd1 vssd1 vccd1 vccd1 _4398_/B sky130_fd_sc_hd__clkbuf_8
X_4329_ _3668_/X _2966_/A _4336_/S vssd1 vssd1 vccd1 vccd1 _4329_/X sky130_fd_sc_hd__mux2_1
Xfanout134 hold640/X vssd1 vssd1 vccd1 vccd1 _3112_/A sky130_fd_sc_hd__clkbuf_4
Xfanout178 fanout184/X vssd1 vssd1 vccd1 vccd1 fanout178/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__5248__A2 _5250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout167 _5507_/A vssd1 vssd1 vccd1 vccd1 _3539_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4471__A3 _4779_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3967__C1 _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3431__A1 _3193_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3613__A _3968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5239__A2 _5107_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5304__S _5305_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5355__A1_N _5341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3700_ _6176_/Q _3910_/C vssd1 vssd1 vccd1 vccd1 _3912_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4680_ _5764_/B _4678_/X _4679_/X vssd1 vssd1 vccd1 vccd1 _4680_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5175__A1 _6176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3631_ _6070_/Q _5333_/B vssd1 vssd1 vccd1 vccd1 _3652_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4922__A1 _6197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3562_ _3540_/A _3561_/X _4446_/A vssd1 vssd1 vccd1 vccd1 _3562_/Y sky130_fd_sc_hd__o21ai_1
X_5301_ hold112/X _3836_/X _5305_/S vssd1 vssd1 vccd1 vccd1 _5301_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3507__B _5502_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3493_ _3491_/X _3492_/Y _3715_/B vssd1 vssd1 vccd1 vccd1 _5955_/D sky130_fd_sc_hd__mux2_1
X_5232_ hold604/X _3353_/B _5217_/A _5231_/X vssd1 vssd1 vccd1 vccd1 _5232_/X sky130_fd_sc_hd__a22o_1
XANTENNA__3489__B2 _5424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5163_ _5163_/A _5163_/B _5163_/C _5163_/D vssd1 vssd1 vccd1 vccd1 _5163_/X sky130_fd_sc_hd__or4_1
X_4114_ hold284/X _3979_/X _4115_/S vssd1 vssd1 vccd1 vccd1 _5912_/D sky130_fd_sc_hd__mux2_1
X_5094_ _3228_/B _3442_/X _5093_/Y _4618_/C vssd1 vssd1 vccd1 vccd1 _5094_/X sky130_fd_sc_hd__o31a_1
X_4045_ _4045_/A _4125_/C vssd1 vssd1 vccd1 vccd1 _4045_/X sky130_fd_sc_hd__or2_1
XFILLER_0_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3661__B2 _6113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3669__S _4035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5402__A2 _6174_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__6058__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5996_ _6151_/CLK _5996_/D vssd1 vssd1 vccd1 vccd1 _5996_/Q sky130_fd_sc_hd__dfxtp_1
X_4947_ _4943_/B _4946_/X _4963_/A vssd1 vssd1 vccd1 vccd1 _4947_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4878_ hold330/X _4877_/X _4927_/S vssd1 vssd1 vccd1 vccd1 _4878_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5166__A1 _6158_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3829_ _3624_/Y _5375_/B _3825_/X _3828_/X vssd1 vssd1 vccd1 vccd1 _3829_/Y sky130_fd_sc_hd__a211oi_2
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3716__A2 _4043_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4913__B2 _4915_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3433__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4524__S0 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold630_A _6160_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4904__A1 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4904__B2 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4840__B1 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5850_ _3785_/Y _5834_/X _5837_/X _5849_/X vssd1 vssd1 vccd1 vccd1 _5850_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_75_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5781_ _6243_/Q hold468/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5781_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4199__A2 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2993_ _2993_/A vssd1 vssd1 vccd1 vccd1 _5551_/A sky130_fd_sc_hd__inv_2
XFILLER_0_8_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4801_ _4800_/X _6055_/Q _5595_/S vssd1 vssd1 vccd1 vccd1 _4801_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4732_ _4725_/X _4730_/X _4731_/X _4412_/B vssd1 vssd1 vccd1 vccd1 _4732_/X sky130_fd_sc_hd__a22o_1
X_4663_ hold480/X _4612_/B _4662_/X _4474_/X vssd1 vssd1 vccd1 vccd1 _4663_/X sky130_fd_sc_hd__a22o_1
X_3614_ _3988_/A _3983_/S _3793_/D vssd1 vssd1 vccd1 vccd1 _4263_/A sky130_fd_sc_hd__or3_4
XANTENNA__4113__S _4115_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4594_ _4594_/A _4594_/B vssd1 vssd1 vccd1 vccd1 _4594_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3545_ _3545_/A _5078_/B vssd1 vssd1 vccd1 vccd1 _3545_/Y sky130_fd_sc_hd__nor2_2
X_3476_ _3303_/A _5424_/C _3475_/X vssd1 vssd1 vccd1 vccd1 _3476_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_86_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5215_ _5023_/A hold408/X _5086_/Y _5214_/X vssd1 vssd1 vccd1 vccd1 _5215_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_6195_ _6211_/CLK _6195_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6195_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5871__A2 _5836_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5146_ _3745_/X _5105_/B _5145_/X vssd1 vssd1 vccd1 vccd1 _5146_/X sky130_fd_sc_hd__a21o_1
X_5077_ _3082_/Y _3543_/B _4750_/A _4391_/B _4416_/C vssd1 vssd1 vccd1 vccd1 _5078_/C
+ sky130_fd_sc_hd__a221o_1
X_4028_ _3958_/S _4028_/B vssd1 vssd1 vccd1 vccd1 _4028_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_79_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5979_ _6129_/CLK _5979_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _5979_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4898__A0 _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4958__S _5020_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5643__A _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3570__B1 _5023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4259__A _5209_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3322__B1 _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5614__A2 _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3928__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold209 _5921_/Q vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4868__S _5011_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3330_ _3289_/A _3328_/Y _3395_/B vssd1 vssd1 vccd1 vccd1 _3334_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _6202_/Q _4766_/Y _4992_/X _4999_/X vssd1 vssd1 vccd1 vccd1 _5000_/X sky130_fd_sc_hd__a211o_1
X_3261_ _3303_/A _3554_/A _4044_/B vssd1 vssd1 vccd1 vccd1 _3261_/X sky130_fd_sc_hd__a21o_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ _4417_/A _3192_/B vssd1 vssd1 vccd1 vccd1 _4439_/B sky130_fd_sc_hd__nor2_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5161__S0 _5185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5902_ _6130_/CLK _5902_/D fanout171/X vssd1 vssd1 vccd1 vccd1 _5902_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__5081__A3 _4036_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4108__S _4115_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5369__A1 _6170_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5833_ _6043_/Q _5834_/B _5834_/C _5834_/D vssd1 vssd1 vccd1 vccd1 _5837_/B sky130_fd_sc_hd__nor4_1
XFILLER_0_17_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5764_ _5767_/B _5764_/B vssd1 vssd1 vccd1 vccd1 _5764_/X sky130_fd_sc_hd__or2_1
X_2976_ _6137_/Q vssd1 vssd1 vccd1 vccd1 _2976_/Y sky130_fd_sc_hd__inv_2
XANTENNA__4041__A1 _4070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5695_ _4990_/Y _5694_/Y _5704_/S vssd1 vssd1 vccd1 vccd1 _5695_/X sky130_fd_sc_hd__a21o_1
X_4715_ _4715_/A _4715_/B vssd1 vssd1 vccd1 vccd1 _4716_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4646_ _4647_/A _4647_/C _4647_/B vssd1 vssd1 vccd1 vccd1 _4648_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4577_ _4575_/X _4577_/B vssd1 vssd1 vccd1 vccd1 _4579_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3147__A3 _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4778__S _5216_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__6243__SET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3528_ _6041_/Q _5790_/D vssd1 vssd1 vccd1 vccd1 _5834_/B sky130_fd_sc_hd__nand2_1
X_6247_ _6247_/CLK _6247_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6247_/Q sky130_fd_sc_hd__dfrtp_1
X_3459_ hold567/X _4446_/A _3713_/A _3458_/X vssd1 vssd1 vccd1 vccd1 _3459_/X sky130_fd_sc_hd__a31o_1
X_6178_ _6178_/CLK _6178_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6178_/Q sky130_fd_sc_hd__dfstp_2
X_5129_ _5129_/A _5129_/B vssd1 vssd1 vccd1 vccd1 _5129_/Y sky130_fd_sc_hd__nor2_2
XANTENNA__6294__A _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3711__A _4759_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3605__B _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5312__S _5313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3068__A _3434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5480_ _6179_/Q _5394_/B _5480_/S vssd1 vssd1 vccd1 vccd1 _5480_/X sky130_fd_sc_hd__mux2_1
X_4500_ _4498_/X _4500_/B vssd1 vssd1 vccd1 vccd1 _4501_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4598__S _4598_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_1 _3306_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4431_ _4070_/B _4731_/S _3320_/B vssd1 vssd1 vccd1 vccd1 _4431_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_1_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4362_ _4242_/X hold133/X _4363_/S vssd1 vssd1 vccd1 vccd1 _4362_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_1_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6101_ _6208_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _4485_/B _3294_/X _3298_/Y _3312_/X vssd1 vssd1 vccd1 vccd1 _3343_/A sky130_fd_sc_hd__a31o_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4293_ _3668_/X hold296/X _4300_/S vssd1 vssd1 vccd1 vccd1 _4293_/X sky130_fd_sc_hd__mux2_1
X_6032_ _6032_/CLK _6032_/D vssd1 vssd1 vccd1 vccd1 _6032_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _3643_/A _3237_/Y _3242_/X _3243_/X vssd1 vssd1 vccd1 vccd1 _5093_/B sky130_fd_sc_hd__o211a_2
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3531__A _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3175_ _5502_/B _3479_/B _3488_/B vssd1 vssd1 vccd1 vccd1 _3176_/D sky130_fd_sc_hd__or3_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3250__B _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5816_ _5815_/X _3864_/Y _5831_/S vssd1 vssd1 vccd1 vccd1 _5816_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_91_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5747_ _3707_/X _5771_/S _5742_/Y _5746_/X vssd1 vssd1 vccd1 vccd1 _5747_/X sky130_fd_sc_hd__o22a_1
X_2959_ _6172_/Q vssd1 vssd1 vccd1 vccd1 _2959_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5678_ _6201_/Q _5685_/B vssd1 vssd1 vccd1 vccd1 _5678_/Y sky130_fd_sc_hd__nand2_1
X_4629_ _4699_/A _4629_/B vssd1 vssd1 vccd1 vccd1 _4630_/B sky130_fd_sc_hd__nand2_1
Xhold562 _5623_/X vssd1 vssd1 vccd1 vccd1 _6196_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold551 _5736_/X vssd1 vssd1 vccd1 vccd1 _6210_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold540 _6057_/Q vssd1 vssd1 vccd1 vccd1 hold540/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 _6242_/Q vssd1 vssd1 vccd1 vccd1 hold595/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 _6116_/Q vssd1 vssd1 vccd1 vccd1 hold573/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 _5739_/X vssd1 vssd1 vccd1 vccd1 _6211_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_49_wb_clk_i_A _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout77_A _3717_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5753__A1 _3832_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5307__S _5313_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5505__A1 _6127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5646__A1_N _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4492__A1 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4881__S _4963_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4980_ _4976_/B _4979_/X _5011_/S vssd1 vssd1 vccd1 vccd1 _4980_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4244__A1 _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5441__B1 _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3931_ hold232/X _3930_/X _4035_/S vssd1 vssd1 vccd1 vccd1 _5897_/D sky130_fd_sc_hd__mux2_1
XANTENNA__4795__A2 _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3862_ _4538_/B _3861_/X _6074_/Q vssd1 vssd1 vccd1 vccd1 _3862_/X sky130_fd_sc_hd__mux2_1
XANTENNA__5744__A1 _3664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5601_ _6161_/Q _5507_/Y _5508_/X vssd1 vssd1 vccd1 vccd1 _5698_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_39_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3793_ _5999_/Q _3988_/A _3795_/C _3793_/D vssd1 vssd1 vccd1 vccd1 _3793_/X sky130_fd_sc_hd__and4_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5532_ _5531_/X hold512/X _5566_/S vssd1 vssd1 vccd1 vccd1 _5532_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5463_ _5330_/B _5462_/X _5363_/C vssd1 vssd1 vccd1 vccd1 _5463_/X sky130_fd_sc_hd__o21a_1
X_5394_ _5394_/A _5394_/B vssd1 vssd1 vccd1 vccd1 _5400_/A sky130_fd_sc_hd__xor2_1
X_4414_ _3121_/X _3309_/B _4413_/X _3715_/B vssd1 vssd1 vccd1 vccd1 _4415_/B sky130_fd_sc_hd__a22o_1
X_4345_ hold227/X _4034_/X _4345_/S vssd1 vssd1 vccd1 vccd1 _6011_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_94_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4276_ hold62/X _4165_/X _4282_/S vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__mux2_1
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6015_ _6035_/CLK _6015_/D vssd1 vssd1 vccd1 vccd1 _6015_/Q sky130_fd_sc_hd__dfxtp_1
X_3227_ _3426_/A _3227_/B vssd1 vssd1 vccd1 vccd1 _3228_/B sky130_fd_sc_hd__nor2_1
X_3158_ _3158_/A _3158_/B _3158_/C _3157_/X vssd1 vssd1 vccd1 vccd1 _3158_/X sky130_fd_sc_hd__or4b_1
XFILLER_0_96_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3089_ _6258_/Q _6259_/Q _3643_/A vssd1 vssd1 vccd1 vccd1 _3125_/C sky130_fd_sc_hd__nand3b_4
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5735__A1 _3959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5196__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3436__A _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5499__B1 _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_wb_clk_i_A _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold381 _5495_/X vssd1 vssd1 vccd1 vccd1 _6185_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold370 _3393_/X vssd1 vssd1 vccd1 vccd1 _5917_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold392 _6190_/Q vssd1 vssd1 vccd1 vccd1 _2992_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__3171__A _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3602__C _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5726__A1 _3832_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_11_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6029_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__4433__C _5838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4130_ _6041_/Q _6042_/Q _6043_/Q _5834_/C _5834_/D vssd1 vssd1 vccd1 vccd1 _4130_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4177__A _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5111__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4061_ _4061_/A _6125_/Q _4061_/C _4061_/D vssd1 vssd1 vccd1 vccd1 _4061_/X sky130_fd_sc_hd__and4_1
XANTENNA__5662__B1 _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4465__B2 _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3512__C _5424_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3012_ _3182_/A _3012_/B vssd1 vssd1 vccd1 vccd1 _4728_/A sky130_fd_sc_hd__nor2_1
X_4963_ _4963_/A _4963_/B vssd1 vssd1 vccd1 vccd1 _4963_/X sky130_fd_sc_hd__or2_1
XFILLER_0_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3914_ _6140_/Q _3914_/B vssd1 vssd1 vccd1 vccd1 _4012_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_46_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5717__A1 _3664_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4894_ hold313/X _4893_/X _4927_/S vssd1 vssd1 vccd1 vccd1 _4894_/X sky130_fd_sc_hd__mux2_1
X_3845_ _6139_/Q _3648_/A _3920_/A _5397_/A _3843_/X vssd1 vssd1 vccd1 vccd1 _3845_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3776_ _3648_/A _5403_/A _5396_/A _3920_/A _3624_/Y vssd1 vssd1 vccd1 vccd1 _3776_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout127_A _3426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5515_ _6054_/Q _6188_/Q _5606_/S vssd1 vssd1 vccd1 vccd1 _5515_/X sky130_fd_sc_hd__mux2_1
X_5446_ hold514/X _5773_/B _5444_/Y _5457_/A vssd1 vssd1 vccd1 vccd1 _5446_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4153__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout113 _5772_/S vssd1 vssd1 vccd1 vccd1 _5832_/S sky130_fd_sc_hd__clkbuf_4
Xfanout102 _5872_/A vssd1 vssd1 vccd1 vccd1 _5762_/A sky130_fd_sc_hd__buf_4
X_5377_ _5377_/A _5377_/B vssd1 vssd1 vccd1 vccd1 _5378_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4328_ _5297_/A _4346_/A vssd1 vssd1 vccd1 vccd1 _4336_/S sky130_fd_sc_hd__or2_4
Xfanout124 _3556_/A vssd1 vssd1 vccd1 vccd1 _4739_/A sky130_fd_sc_hd__buf_4
Xfanout146 _6125_/Q vssd1 vssd1 vccd1 vccd1 _4038_/A sky130_fd_sc_hd__clkbuf_8
Xfanout135 _6252_/Q vssd1 vssd1 vccd1 vccd1 _3203_/B sky130_fd_sc_hd__clkbuf_8
Xfanout179 fanout180/X vssd1 vssd1 vccd1 vccd1 fanout179/X sky130_fd_sc_hd__clkbuf_8
X_4259_ _5209_/A _4259_/B _4259_/C vssd1 vssd1 vccd1 vccd1 _4259_/X sky130_fd_sc_hd__or3_1
Xfanout157 _5164_/A1 vssd1 vssd1 vccd1 vccd1 _5023_/A sky130_fd_sc_hd__clkbuf_8
Xfanout168 _5916_/Q vssd1 vssd1 vccd1 vccd1 _5507_/A sky130_fd_sc_hd__buf_4
XANTENNA__4456__A1 _4478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold506_A _6205_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4916__C1 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5978__CLK _5978_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3613__B _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4447__A1 _3446_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3775__S _5868_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4460__A _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3630_ _6072_/Q _6172_/Q vssd1 vssd1 vccd1 vccd1 _3634_/S sky130_fd_sc_hd__and2b_1
XANTENNA__4922__A2 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3561_ _3507_/C _3125_/C _4398_/B vssd1 vssd1 vccd1 vccd1 _3561_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5300_ hold74/X _3789_/X _5305_/S vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__mux2_1
XANTENNA__3507__C _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3492_ _3461_/A _3503_/C _4478_/A vssd1 vssd1 vccd1 vccd1 _3492_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__4686__A1 _4976_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5231_ _5225_/B _5228_/B _5220_/Y _5218_/X _4765_/A vssd1 vssd1 vccd1 vccd1 _5231_/X
+ sky130_fd_sc_hd__a32o_1
X_5162_ _6239_/Q _5108_/Y _5109_/Y _5161_/X vssd1 vssd1 vccd1 vccd1 _5163_/D sky130_fd_sc_hd__a22o_1
X_4113_ hold98/X _3930_/X _4115_/S vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__mux2_1
X_5093_ _5093_/A _5093_/B vssd1 vssd1 vccd1 vccd1 _5093_/Y sky130_fd_sc_hd__nor2_1
X_4044_ _4085_/B _4044_/B vssd1 vssd1 vccd1 vccd1 _4125_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5995_ _6146_/CLK _5995_/D vssd1 vssd1 vccd1 vccd1 _5995_/Q sky130_fd_sc_hd__dfxtp_1
X_4946_ _6199_/Q _6065_/Q _6038_/Q vssd1 vssd1 vccd1 vccd1 _4946_/X sky130_fd_sc_hd__mux2_1
X_4877_ _4876_/X _6060_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _4877_/X sky130_fd_sc_hd__mux2_1
X_3828_ hold573/X _3826_/X _3827_/X _3645_/X _3824_/X vssd1 vssd1 vccd1 vccd1 _3828_/X
+ sky130_fd_sc_hd__a221o_1
X_3759_ _3759_/A _5052_/B vssd1 vssd1 vccd1 vccd1 _3759_/X sky130_fd_sc_hd__or2_1
X_5429_ hold567/X _5488_/S _5427_/Y _5428_/Y vssd1 vssd1 vccd1 vccd1 _5429_/X sky130_fd_sc_hd__o22a_1
XANTENNA__6297__A _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5874__B1 _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3433__B _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4524__S1 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold623_A _6157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3404__A2 _5838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4062__C1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5865__A0 _6119_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3624__A _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4439__B _4439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4800_ _5606_/S _4799_/X _4790_/X vssd1 vssd1 vccd1 vccd1 _4800_/X sky130_fd_sc_hd__a21o_1
X_5780_ _6242_/Q hold472/X _5789_/S vssd1 vssd1 vccd1 vccd1 _5780_/X sky130_fd_sc_hd__mux2_1
X_2992_ _2992_/A vssd1 vssd1 vccd1 vccd1 _5538_/A sky130_fd_sc_hd__inv_2
X_4731_ _6259_/Q _4739_/A _4731_/S vssd1 vssd1 vccd1 vccd1 _4731_/X sky130_fd_sc_hd__mux2_1
X_4662_ _4662_/A _4662_/B vssd1 vssd1 vccd1 vccd1 _4662_/X sky130_fd_sc_hd__xor2_1
XANTENNA__4190__A _4223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6191__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3613_ _3968_/A _3616_/B _3982_/S vssd1 vssd1 vccd1 vccd1 _3613_/X sky130_fd_sc_hd__and3_4
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3159__A1 _3277_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4593_ _4577_/B _4579_/B _4575_/X vssd1 vssd1 vccd1 vccd1 _4594_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3544_ _3488_/A _3543_/B _5498_/B _3221_/X _3396_/A vssd1 vssd1 vccd1 vccd1 _5078_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_3_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3475_ _3563_/A _3422_/B _4446_/B vssd1 vssd1 vccd1 vccd1 _3475_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5214_ _6211_/Q _5106_/Y _5108_/Y _6243_/Q _5213_/X vssd1 vssd1 vccd1 vccd1 _5214_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5856__A0 _6135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6194_ _6194_/CLK _6194_/D fanout184/X vssd1 vssd1 vccd1 vccd1 _6194_/Q sky130_fd_sc_hd__dfrtp_2
X_5145_ _5116_/A _4179_/X _5185_/S _5144_/X vssd1 vssd1 vccd1 vccd1 _5145_/X sky130_fd_sc_hd__o211a_1
XANTENNA__3882__A2 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5076_ _5076_/A0 _5075_/Y _5296_/S vssd1 vssd1 vccd1 vccd1 _6112_/D sky130_fd_sc_hd__mux2_1
X_4027_ _6161_/Q _4026_/X _6074_/Q vssd1 vssd1 vccd1 vccd1 _4028_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_47_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5978_ _5978_/CLK _5978_/D fanout170/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4929_ _6238_/Q _5008_/B vssd1 vssd1 vccd1 vccd1 _4929_/X sky130_fd_sc_hd__and2_1
XFILLER_0_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4304__S _4309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5362__C _5424_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold573_A _6116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__3561__A1 _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3354__A _6129_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3313__A1 _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _6125_/Q _3446_/A vssd1 vssd1 vccd1 vccd1 _4446_/B sky130_fd_sc_hd__nand2_4
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3191_ _3302_/A _4070_/B _4412_/A vssd1 vssd1 vccd1 vccd1 _3198_/B sky130_fd_sc_hd__a21oi_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5161__S1 _5116_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4813__A1 _6156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4813__B2 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5901_ _6167_/CLK _5901_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _5901_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5832_ hold591/X _5831_/X _5832_/S vssd1 vssd1 vccd1 vccd1 _6243_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5763_ _5761_/Y _5762_/X _4119_/A vssd1 vssd1 vccd1 vccd1 _5763_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_56_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4714_ _6219_/Q _5007_/B _4714_/S vssd1 vssd1 vccd1 vccd1 _4715_/B sky130_fd_sc_hd__mux2_1
X_2975_ _6136_/Q vssd1 vssd1 vccd1 vccd1 _2975_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4041__A2 _4446_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5694_ _5694_/A _5694_/B vssd1 vssd1 vccd1 vccd1 _5694_/Y sky130_fd_sc_hd__nand2_1
X_4645_ _4609_/A _4609_/B _4628_/Y _4630_/B vssd1 vssd1 vccd1 vccd1 _4647_/C sky130_fd_sc_hd__o31a_1
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3963__S _3983_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4576_ _4575_/A _4575_/B _4575_/C vssd1 vssd1 vccd1 vccd1 _4577_/B sky130_fd_sc_hd__a21o_1
XANTENNA__5541__A2 _5606_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3527_ _3527_/A _4129_/B vssd1 vssd1 vccd1 vccd1 _5740_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3552__A1 _3457_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_wb_clk_i_A clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__3264__A _5838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6246_ _6246_/CLK _6246_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6246_/Q sky130_fd_sc_hd__dfrtp_1
XANTENNA__3304__A1 _5424_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3458_ hold567/X _5424_/A _2960_/Y vssd1 vssd1 vccd1 vccd1 _3458_/X sky130_fd_sc_hd__o21a_1
X_6177_ _6233_/CLK _6177_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6177_/Q sky130_fd_sc_hd__dfstp_2
X_3389_ _4415_/A _3389_/B hold92/X _3517_/B vssd1 vssd1 vccd1 vccd1 _3389_/X sky130_fd_sc_hd__or4b_1
XANTENNA__5798__A2_N _5352_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5128_ _5164_/A1 hold363/X _5086_/Y _5127_/X vssd1 vssd1 vccd1 vccd1 _5128_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4804__A1 _4803_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5059_ _5059_/A vssd1 vssd1 vccd1 vccd1 _6096_/D sky130_fd_sc_hd__inv_2
XFILLER_0_94_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__6042__RESET_B fanout183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4568__A0 _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold419_A _6137_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4032__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4034__S _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_36_wb_clk_i clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6246_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5296__A1 _5250_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4654__S0 _4712_/S0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4023__A2 _6141_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3349__A _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__3068__B _4116_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_2 _3404_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ _3488_/B _4759_/A _4446_/B _3193_/C _4429_/X vssd1 vssd1 vccd1 vccd1 _4430_/X
+ sky130_fd_sc_hd__a221o_1
X_4361_ _4226_/X hold228/X _4363_/S vssd1 vssd1 vccd1 vccd1 _4361_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_67_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6100_ _6208_/CLK hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4292_ _5297_/A _4292_/B vssd1 vssd1 vccd1 vccd1 _4300_/S sky130_fd_sc_hd__or2_4
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ _5838_/A _3321_/B _3311_/Y _5918_/Q _6130_/Q vssd1 vssd1 vccd1 vccd1 _3312_/X
+ sky130_fd_sc_hd__a221o_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_6031_ _6031_/CLK _6031_/D vssd1 vssd1 vccd1 vccd1 _6031_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _4085_/B _3116_/B _6179_/Q vssd1 vssd1 vccd1 vccd1 _3243_/X sky130_fd_sc_hd__mux2_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _4417_/A _3182_/B vssd1 vssd1 vccd1 vccd1 _3463_/A sky130_fd_sc_hd__or2_1
XFILLER_0_76_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3250__C _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5815_ hold427/X _5794_/Y _5814_/X _5794_/B vssd1 vssd1 vccd1 vccd1 _5815_/X sky130_fd_sc_hd__a22o_1
XANTENNA_fanout157_A _5164_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__3259__A _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5746_ _4119_/A _4915_/B _4632_/X _5762_/C vssd1 vssd1 vccd1 vccd1 _5746_/X sky130_fd_sc_hd__o22a_1
X_2958_ _6174_/Q vssd1 vssd1 vccd1 vccd1 _2958_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3222__B1 _4124_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5677_ _5679_/A _5685_/B vssd1 vssd1 vccd1 vccd1 _5682_/A sky130_fd_sc_hd__and2_1
XFILLER_0_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5474__A _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4628_ _4699_/A _4629_/B vssd1 vssd1 vccd1 vccd1 _4628_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold530 _4456_/X vssd1 vssd1 vccd1 vccd1 _6050_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4722__B1 _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold563 _6208_/Q vssd1 vssd1 vccd1 vccd1 hold563/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 _6060_/Q vssd1 vssd1 vccd1 vccd1 hold552/X sky130_fd_sc_hd__buf_1
X_4559_ _4575_/A _4559_/B _4559_/C vssd1 vssd1 vccd1 vccd1 _4561_/A sky130_fd_sc_hd__nand3_1
Xhold541 _4537_/X vssd1 vssd1 vccd1 vccd1 _6057_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 _6241_/Q vssd1 vssd1 vccd1 vccd1 _2990_/A sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5278__A1 _5245_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold574 _6256_/Q vssd1 vssd1 vccd1 vccd1 hold574/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold585 _6076_/Q vssd1 vssd1 vccd1 vccd1 _5228_/B sky130_fd_sc_hd__buf_1
X_6229_ _6251_/CLK _6229_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6229_/Q sky130_fd_sc_hd__dfstp_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold369_A _5917_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4253__A2 _4253_/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5450__B2 _6176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4272__B _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5753__A2 _5771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4961__B1 _4769_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3616__B _3616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput50 _5953_/Q vssd1 vssd1 vccd1 vccd1 io_out[6] sky130_fd_sc_hd__buf_12
XFILLER_0_101_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4477__C1 _3252_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5441__A1 _3832_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3930_ _3928_/X _3929_/X _4034_/S vssd1 vssd1 vccd1 vccd1 _3930_/X sky130_fd_sc_hd__mux2_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__3452__B1 _3210_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3861_ _3623_/X _3860_/A _3846_/X vssd1 vssd1 vccd1 vccd1 _3861_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_46_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5744__A2 _5771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5600_ _2996_/A _5599_/X _5672_/S vssd1 vssd1 vccd1 vccd1 _5600_/X sky130_fd_sc_hd__mux2_1
X_3792_ hold112/X _3611_/X _3613_/X hold163/X vssd1 vssd1 vccd1 vccd1 _3798_/C sky130_fd_sc_hd__a22o_1
XFILLER_0_26_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5531_ _5530_/X _6055_/Q _5609_/S vssd1 vssd1 vccd1 vccd1 _5531_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_81_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5462_ _6177_/Q _5026_/A _5460_/X _5025_/A _5461_/X vssd1 vssd1 vccd1 vccd1 _5462_/X
+ sky130_fd_sc_hd__a221o_1
X_5393_ _5392_/A _5392_/B _5033_/A vssd1 vssd1 vccd1 vccd1 _5393_/X sky130_fd_sc_hd__a21o_1
XANTENNA__3526__B _5566_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4413_ _4413_/A _4729_/B _4413_/C _4413_/D vssd1 vssd1 vccd1 vccd1 _4413_/X sky130_fd_sc_hd__or4_1
X_4344_ hold285/X _3979_/X _4345_/S vssd1 vssd1 vccd1 vccd1 _6010_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_1_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_6014_ _6014_/CLK _6014_/D vssd1 vssd1 vccd1 vccd1 _6014_/Q sky130_fd_sc_hd__dfxtp_1
X_4275_ hold169/X _4150_/X _4282_/S vssd1 vssd1 vccd1 vccd1 _4275_/X sky130_fd_sc_hd__mux2_1
X_3226_ _4124_/A _4451_/C vssd1 vssd1 vccd1 vccd1 _3283_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3691__A0 _6114_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3157_ _4433_/A _3157_/B _3157_/C _3157_/D vssd1 vssd1 vccd1 vccd1 _3157_/X sky130_fd_sc_hd__and4b_1
XFILLER_0_68_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3088_ _3105_/A _6258_/Q vssd1 vssd1 vccd1 vccd1 _4412_/A sky130_fd_sc_hd__or2_4
XFILLER_0_49_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5735__A2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5196__B1 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5729_ _3864_/Y _5715_/B _5715_/Y _5728_/X vssd1 vssd1 vccd1 vccd1 _5729_/X sky130_fd_sc_hd__o22a_1
XANTENNA__4312__S _4318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5499__A1 _5609_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3436__B _4618_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold371 _6180_/Q vssd1 vssd1 vccd1 vccd1 hold371/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold360 _4459_/X vssd1 vssd1 vccd1 vccd1 _6052_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold382 _6078_/Q vssd1 vssd1 vccd1 vccd1 hold382/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold393 _5548_/X vssd1 vssd1 vccd1 vccd1 _6190_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5671__A1 _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4982__S _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4934__A0 _6156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5726__A2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3737__A1 _4034_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3627__A _6135_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3362__A _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5111__B1 _3740_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4060_ _4618_/B _4050_/X _4059_/X vssd1 vssd1 vccd1 vccd1 _5250_/A sky130_fd_sc_hd__o21a_4
XANTENNA__5662__A1 _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4465__A2 _4618_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3011_ _3511_/C vssd1 vssd1 vccd1 vccd1 _3012_/B sky130_fd_sc_hd__inv_2
XFILLER_0_59_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4962_ _6200_/Q _6066_/Q _5216_/A vssd1 vssd1 vccd1 vccd1 _4962_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_86_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3913_ _6140_/Q _3914_/B vssd1 vssd1 vccd1 vccd1 _4009_/C sky130_fd_sc_hd__or2_1
X_4893_ _4892_/X _6061_/Q _4926_/S vssd1 vssd1 vccd1 vccd1 _4893_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3844_ _6138_/Q _6140_/Q _5868_/S vssd1 vssd1 vccd1 vccd1 _5397_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_73_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5717__A2 _5715_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3775_ _6136_/Q _6138_/Q _5868_/S vssd1 vssd1 vccd1 vccd1 _5396_/A sky130_fd_sc_hd__mux2_1
XANTENNA__3537__A _4460_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5514_ _5514_/A _5514_/B vssd1 vssd1 vccd1 vccd1 _5514_/X sky130_fd_sc_hd__xor2_1
X_5445_ _5445_/A _5872_/A vssd1 vssd1 vccd1 vccd1 _5445_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5376_ _5376_/A _5376_/B vssd1 vssd1 vccd1 vccd1 _5377_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout103 _3377_/X vssd1 vssd1 vccd1 vccd1 _5872_/A sky130_fd_sc_hd__buf_8
Xfanout125 hold574/X vssd1 vssd1 vccd1 vccd1 _3556_/A sky130_fd_sc_hd__buf_4
Xfanout136 hold556/X vssd1 vssd1 vccd1 vccd1 _4497_/S sky130_fd_sc_hd__buf_8
Xfanout147 _3302_/A vssd1 vssd1 vccd1 vccd1 _3540_/A sky130_fd_sc_hd__buf_4
Xfanout114 _2968_/Y vssd1 vssd1 vccd1 vccd1 _5772_/S sky130_fd_sc_hd__clkbuf_8
X_4327_ _4034_/X hold168/X _4327_/S vssd1 vssd1 vccd1 vccd1 _5995_/D sky130_fd_sc_hd__mux2_1
X_4258_ hold294/X _5200_/A2 _4255_/S hold278/X _4256_/S vssd1 vssd1 vccd1 vccd1 _4259_/C
+ sky130_fd_sc_hd__o221a_1
Xfanout158 _5245_/A vssd1 vssd1 vccd1 vccd1 _5773_/A sky130_fd_sc_hd__clkbuf_8
Xfanout169 hold590/X vssd1 vssd1 vccd1 vccd1 _4697_/S sky130_fd_sc_hd__buf_6
XANTENNA__5653__A1 _6157_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4456__A2 _3517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3209_ _4433_/A _5838_/B vssd1 vssd1 vccd1 vccd1 _3306_/C sky130_fd_sc_hd__nor2_1
X_4189_ _4195_/B _4189_/B vssd1 vssd1 vccd1 vccd1 _5055_/B sky130_fd_sc_hd__xnor2_1
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4815__B _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4307__S _4309_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3881__S _4035_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold190 _4320_/X vssd1 vssd1 vccd1 vccd1 _5988_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4725__B _4725_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5837__A _5837_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4907__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4460__B _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3560_ _3171_/X _3545_/Y _3547_/X _3541_/X vssd1 vssd1 vccd1 vccd1 _3560_/X sky130_fd_sc_hd__a31o_1
XANTENNA__4383__A1 _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5230_ _4765_/A _3353_/B _5217_/A _5229_/X vssd1 vssd1 vccd1 vccd1 _5230_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3491_ _3523_/B _3491_/B vssd1 vssd1 vccd1 vccd1 _3491_/X sky130_fd_sc_hd__or2_1
X_5161_ _3835_/X _4192_/X _5157_/X _5160_/X _5185_/S _5116_/A vssd1 vssd1 vccd1 vccd1
+ _5161_/X sky130_fd_sc_hd__mux4_2
XANTENNA__3804__B _6116_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4112_ hold120/X _3880_/X _4115_/S vssd1 vssd1 vccd1 vccd1 _4112_/X sky130_fd_sc_hd__mux2_1
X_5092_ _4749_/A _5090_/X _5091_/X _4618_/B vssd1 vssd1 vccd1 vccd1 _5092_/X sky130_fd_sc_hd__o31a_1
XANTENNA__5635__B2 _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4043_ _4043_/A _5502_/B _4043_/C vssd1 vssd1 vccd1 vccd1 _4048_/B sky130_fd_sc_hd__and3_1
XFILLER_0_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5994_ _6010_/CLK _5994_/D vssd1 vssd1 vccd1 vccd1 _5994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4945_ _6215_/Q _5009_/A2 _4769_/Y _4943_/B _4944_/X vssd1 vssd1 vccd1 vccd1 _4945_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4876_ _4119_/B _4875_/X _4865_/Y vssd1 vssd1 vccd1 vccd1 _4876_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_19_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3827_ _6116_/Q _3827_/B vssd1 vssd1 vccd1 vccd1 _3827_/X sky130_fd_sc_hd__or2_1
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3758_ _3759_/A _5052_/B vssd1 vssd1 vccd1 vccd1 _3758_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3689_ _3848_/B _3686_/X _3687_/Y _3688_/X vssd1 vssd1 vccd1 vccd1 _3689_/X sky130_fd_sc_hd__a31o_1
X_5428_ _3785_/A _5487_/S _5488_/S vssd1 vssd1 vccd1 vccd1 _5428_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_2_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5359_ _6173_/Q _5341_/A _5794_/B _5358_/X vssd1 vssd1 vccd1 vccd1 _5359_/X sky130_fd_sc_hd__o211a_1
XANTENNA__5874__A1 hold652/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3433__C _5341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3730__A _4234_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold616_A _6176_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3363__D_N _3370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5617__A1 _6196_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output33_A _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2991_ _6189_/Q vssd1 vssd1 vccd1 vccd1 _5524_/A sky130_fd_sc_hd__inv_2
XFILLER_0_56_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4730_ _3446_/A _3192_/B _4413_/D _4729_/X vssd1 vssd1 vccd1 vccd1 _4730_/X sky130_fd_sc_hd__a211o_1
X_4661_ _4699_/A _4643_/B _4648_/A vssd1 vssd1 vccd1 vccd1 _4662_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_16_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3612_ _3988_/A _3983_/S _3982_/S vssd1 vssd1 vccd1 vccd1 _5297_/B sky130_fd_sc_hd__or3_4
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4592_ _4590_/X _4592_/B vssd1 vssd1 vccd1 vccd1 _4594_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_29_wb_clk_i_A clkbuf_2_3__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_3543_ _3543_/A _3543_/B vssd1 vssd1 vccd1 vccd1 _3543_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3474_ _3715_/B _3473_/X _3462_/Y vssd1 vssd1 vccd1 vccd1 _3474_/Y sky130_fd_sc_hd__o21ai_1
X_5213_ _6203_/Q _5119_/Y _5211_/X _5109_/Y _5212_/X vssd1 vssd1 vccd1 vccd1 _5213_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__5856__A1 _6113_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6193_ _6194_/CLK _6193_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6193_/Q sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_2_2__f_wb_clk_i_A clkbuf_0_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5144_ _5209_/A _5144_/B _5144_/C vssd1 vssd1 vccd1 vccd1 _5144_/X sky130_fd_sc_hd__or3_1
XANTENNA__5608__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5075_ _4771_/B _4121_/B _4120_/Y vssd1 vssd1 vccd1 vccd1 _5075_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__5241__S _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4026_ _3624_/Y _5372_/B _4019_/X _4025_/X vssd1 vssd1 vccd1 vccd1 _4026_/X sky130_fd_sc_hd__a211o_1
XANTENNA__4746__A1_N _4485_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5977_ _6038_/CLK _5977_/D fanout170/X vssd1 vssd1 vccd1 vccd1 _5977_/Q sky130_fd_sc_hd__dfrtp_1
X_4928_ _4990_/A _4928_/B vssd1 vssd1 vccd1 vccd1 _4928_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__4595__B2 _4474_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4859_ _6193_/Q _4767_/X _4857_/X _4858_/X vssd1 vssd1 vccd1 vccd1 _4859_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3570__A2 _3671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4320__S _4327_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5362__D _5424_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5783__A0 _6173_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3354__B _6127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _4036_/B _3543_/B _4045_/A vssd1 vssd1 vccd1 vccd1 _3197_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__3370__A _4077_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4466__A _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3077__A1 _3507_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4813__A2 _5008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5900_ _6167_/CLK _5900_/D fanout176/X vssd1 vssd1 vccd1 vccd1 _5900_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3482__D1 _4439_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5831_ _5830_/X _4030_/Y _5831_/S vssd1 vssd1 vccd1 vccd1 _5831_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5774__A0 _6236_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5762_ _5762_/A _5762_/B _5762_/C vssd1 vssd1 vccd1 vccd1 _5762_/X sky130_fd_sc_hd__or3_1
XANTENNA__4405__S _5488_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2974_ _5333_/B vssd1 vssd1 vccd1 vccd1 _3894_/A sky130_fd_sc_hd__inv_2
X_4713_ _4712_/X _4711_/X _5914_/Q vssd1 vssd1 vccd1 vccd1 _5007_/B sky130_fd_sc_hd__mux2_2
Xclkbuf_leaf_6_wb_clk_i _5978_/CLK vssd1 vssd1 vccd1 vccd1 _6148_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5693_ _6068_/Q _4761_/X _5702_/B1 _5692_/X vssd1 vssd1 vccd1 vccd1 _5694_/B sky130_fd_sc_hd__a22o_1
X_4644_ _4676_/A _4644_/B vssd1 vssd1 vccd1 vccd1 _4647_/B sky130_fd_sc_hd__nand2_1
X_4575_ _4575_/A _4575_/B _4575_/C vssd1 vssd1 vccd1 vccd1 _4575_/X sky130_fd_sc_hd__and3_1
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout102_A _5872_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3526_ _3532_/B _5566_/S vssd1 vssd1 vccd1 vccd1 _6123_/D sky130_fd_sc_hd__and2_1
XANTENNA__5829__B2 _5341_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5829__A1 hold591/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_6245_ _6246_/CLK _6245_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6245_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3457_ _3457_/A _5424_/C _4433_/A vssd1 vssd1 vccd1 vccd1 _4377_/B sky130_fd_sc_hd__or3b_1
X_6176_ _6247_/CLK _6176_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6176_/Q sky130_fd_sc_hd__dfstp_4
X_3388_ _3392_/A _3388_/B vssd1 vssd1 vccd1 vccd1 _3517_/B sky130_fd_sc_hd__or2_2
XANTENNA__4376__A _5773_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5127_ _6196_/Q _5119_/Y _5122_/Y _6188_/Q _5126_/X vssd1 vssd1 vccd1 vccd1 _5127_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__3280__A _5502_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5058_ _2999_/Y _5249_/A _5296_/S vssd1 vssd1 vccd1 vccd1 _5059_/A sky130_fd_sc_hd__mux2_1
X_4009_ _5046_/A _6141_/Q _4009_/C vssd1 vssd1 vccd1 vccd1 _4011_/A sky130_fd_sc_hd__or3_1
XFILLER_0_79_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5765__B1 _5771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4315__S _4318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4740__A1 _3488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5670__A _5670_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4179__S0 _5182_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__clkbuf_2
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4654__S1 _4712_/S1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3349__B _3503_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 _3421_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4360_ _4211_/X hold171/X _4363_/S vssd1 vssd1 vccd1 vccd1 _4360_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3311_ _3320_/B vssd1 vssd1 vccd1 vccd1 _3311_/Y sky130_fd_sc_hd__inv_2
X_4291_ _4261_/X hold278/X _4291_/S vssd1 vssd1 vccd1 vccd1 _4291_/X sky130_fd_sc_hd__mux2_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ _6030_/CLK _6030_/D vssd1 vssd1 vccd1 vccd1 _6030_/Q sky130_fd_sc_hd__dfxtp_1
X_3242_ _6174_/Q _3239_/X _3241_/X vssd1 vssd1 vccd1 vccd1 _3242_/X sky130_fd_sc_hd__o21ba_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _4417_/A _3182_/B vssd1 vssd1 vccd1 vccd1 _3488_/B sky130_fd_sc_hd__nor2_4
XFILLER_0_83_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4798__A1 _6205_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5814_ hold594/X _5791_/X _5813_/X _5764_/B vssd1 vssd1 vccd1 vccd1 _5814_/X sky130_fd_sc_hd__a22o_1
XANTENNA__5211__A2 _5185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5745_ hold486/X _5741_/Y _5744_/X _5767_/A vssd1 vssd1 vccd1 vccd1 _5745_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3222__A1 _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2957_ _4415_/A vssd1 vssd1 vccd1 vccd1 _2957_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5676_ _5675_/X _6159_/Q _5704_/S vssd1 vssd1 vccd1 vccd1 _5676_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__5474__B _6154_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4627_ _6213_/Q _4915_/B _4714_/S vssd1 vssd1 vccd1 vccd1 _4629_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_44_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold520 _6064_/Q vssd1 vssd1 vccd1 vccd1 hold520/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__4722__A1 _6161_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold553 _4584_/X vssd1 vssd1 vccd1 vccd1 _6060_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4558_ _6209_/Q _4850_/B _4589_/S vssd1 vssd1 vccd1 vccd1 _4559_/C sky130_fd_sc_hd__mux2_1
Xhold542 _6056_/Q vssd1 vssd1 vccd1 vccd1 hold542/X sky130_fd_sc_hd__buf_1
Xhold531 _6188_/Q vssd1 vssd1 vccd1 vccd1 _5514_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold597 _5822_/X vssd1 vssd1 vccd1 vccd1 _6241_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 _5730_/X vssd1 vssd1 vccd1 vccd1 _6208_/D sky130_fd_sc_hd__dlygate4sd3_1
X_4489_ _4565_/S _4564_/S vssd1 vssd1 vccd1 vccd1 _4612_/B sky130_fd_sc_hd__and2_4
Xhold586 _5237_/X vssd1 vssd1 vccd1 vccd1 hold586/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3509_ _3517_/B _3517_/C vssd1 vssd1 vccd1 vccd1 _3509_/Y sky130_fd_sc_hd__nor2_1
Xhold575 _3460_/Y vssd1 vssd1 vccd1 vccd1 _6095_/D sky130_fd_sc_hd__dlygate4sd3_1
X_6228_ _6233_/CLK _6228_/D fanout180/X vssd1 vssd1 vccd1 vccd1 _6228_/Q sky130_fd_sc_hd__dfstp_1
X_6159_ _6238_/CLK _6159_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6159_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold529_A _6050_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3169__B _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4961__B2 _4963_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput40 _6246_/Q vssd1 vssd1 vccd1 vccd1 io_out[26] sky130_fd_sc_hd__buf_12
Xoutput51 _6078_/Q vssd1 vssd1 vccd1 vccd1 io_out[8] sky130_fd_sc_hd__buf_12
XFILLER_0_101_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4572__S0 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4229__B1 _3613_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3452__A1 _3192_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3860_ _3860_/A vssd1 vssd1 vccd1 vccd1 _5373_/A sky130_fd_sc_hd__inv_2
X_3791_ _5983_/Q _3599_/X _3601_/X _5991_/Q vssd1 vssd1 vccd1 vccd1 _3798_/B sky130_fd_sc_hd__a22o_1
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4952__A1 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4952__B2 _4824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5530_ _4119_/B _5529_/X _4789_/Y vssd1 vssd1 vccd1 vccd1 _5530_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5461_ _6118_/Q _3192_/B _3646_/X _3918_/X _3920_/X vssd1 vssd1 vccd1 vccd1 _5461_/X
+ sky130_fd_sc_hd__a311o_1
XFILLER_0_54_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4412_ _4412_/A _4412_/B vssd1 vssd1 vccd1 vccd1 _4413_/D sky130_fd_sc_hd__nor2_1
X_5392_ _5392_/A _5392_/B vssd1 vssd1 vccd1 vccd1 _5392_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4919__A _6155_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4343_ hold135/X _3930_/X _4345_/S vssd1 vssd1 vccd1 vccd1 _4343_/X sky130_fd_sc_hd__mux2_1
X_4274_ _5297_/B _4364_/B vssd1 vssd1 vccd1 vccd1 _4282_/S sky130_fd_sc_hd__nor2_4
X_6013_ _6034_/CLK _6013_/D vssd1 vssd1 vccd1 vccd1 _6013_/Q sky130_fd_sc_hd__dfxtp_1
X_3225_ _4124_/A _4765_/A vssd1 vssd1 vccd1 vccd1 _4618_/C sky130_fd_sc_hd__and2_4
XFILLER_0_94_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__3691__A1 _6118_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3156_ _3135_/B _3182_/B _4412_/A _3125_/X _3155_/X vssd1 vssd1 vccd1 vccd1 _3157_/D
+ sky130_fd_sc_hd__o311a_1
X_3087_ _3105_/A _6258_/Q vssd1 vssd1 vccd1 vccd1 _3277_/A sky130_fd_sc_hd__nor2_4
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5728_ _4119_/A _4836_/B _4547_/Y _5762_/C vssd1 vssd1 vccd1 vccd1 _5728_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_9_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3989_ _3968_/A _3983_/X _3988_/X vssd1 vssd1 vccd1 vccd1 _3990_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5659_ _5659_/A _5659_/B vssd1 vssd1 vccd1 vccd1 _5664_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold361 _6187_/Q vssd1 vssd1 vccd1 vccd1 hold361/X sky130_fd_sc_hd__buf_1
Xhold350 _5492_/X vssd1 vssd1 vccd1 vccd1 _6182_/D sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold372 _5490_/X vssd1 vssd1 vccd1 vccd1 _6180_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 _6202_/Q vssd1 vssd1 vccd1 vccd1 _5685_/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold383 _4788_/X vssd1 vssd1 vccd1 vccd1 _6078_/D sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3733__A _5249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout82_A _3739_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3985__A2 _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5187__A1 _6177_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3908__A _6172_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4503__S _4596_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__5813__A1_N _6240_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5828__A1_N _6243_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_20_wb_clk_i clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1 _6219_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__3362__B _6047_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5662__A2 _6197_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3010_ _3426_/A _3507_/C vssd1 vssd1 vccd1 vccd1 _3511_/C sky130_fd_sc_hd__nor2_2
XANTENNA__4474__A _4474_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4961_ _6216_/Q _5009_/A2 _4769_/Y _4963_/B _4960_/X vssd1 vssd1 vccd1 vccd1 _4961_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4622__B1 _5767_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3425__A1 _5875_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3912_ _6139_/Q _3912_/B _3912_/C vssd1 vssd1 vccd1 vccd1 _3914_/B sky130_fd_sc_hd__or3_1
X_4892_ _4119_/B _4891_/X _4879_/Y vssd1 vssd1 vccd1 vccd1 _4892_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3843_ _3645_/X _3842_/X _3841_/X vssd1 vssd1 vccd1 vccd1 _3843_/X sky130_fd_sc_hd__o21a_1
XANTENNA__3818__A _6136_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4925__A1 _5694_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3774_ _6115_/Q _6119_/Q _6070_/Q vssd1 vssd1 vccd1 vccd1 _5403_/A sky130_fd_sc_hd__mux2_1
XFILLER_0_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3537__B _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5513_ _6188_/Q _5514_/B vssd1 vssd1 vccd1 vccd1 _5526_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5444_ _4375_/Y _5344_/X _5443_/X vssd1 vssd1 vccd1 vccd1 _5444_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4153__A2 _3611_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5375_ _5375_/A _5375_/B vssd1 vssd1 vccd1 vccd1 _5376_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout104 _5011_/S vssd1 vssd1 vccd1 vccd1 _4963_/A sky130_fd_sc_hd__buf_6
Xfanout115 _5480_/S vssd1 vssd1 vccd1 vccd1 _5502_/A sky130_fd_sc_hd__buf_6
Xfanout137 _6165_/Q vssd1 vssd1 vccd1 vccd1 _4589_/S sky130_fd_sc_hd__buf_4
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout126 _3050_/C vssd1 vssd1 vccd1 vccd1 _4737_/A sky130_fd_sc_hd__buf_4
X_4326_ _3979_/X hold260/X _4327_/S vssd1 vssd1 vccd1 vccd1 _4326_/X sky130_fd_sc_hd__mux2_1
X_4257_ hold211/X _5200_/A2 _4255_/S hold242/X _5182_/S vssd1 vssd1 vccd1 vccd1 _4259_/B
+ sky130_fd_sc_hd__o221a_1
Xfanout159 _5164_/A1 vssd1 vssd1 vccd1 vccd1 _5245_/A sky130_fd_sc_hd__buf_4
Xfanout148 _3302_/A vssd1 vssd1 vccd1 vccd1 _4124_/B sky130_fd_sc_hd__buf_4
X_4188_ _4195_/A _4176_/B _4172_/Y vssd1 vssd1 vccd1 vccd1 _4189_/B sky130_fd_sc_hd__a21bo_1
X_3208_ _3208_/A _3208_/B vssd1 vssd1 vccd1 vccd1 _5838_/B sky130_fd_sc_hd__nor2_4
X_3139_ _4460_/C _3545_/A vssd1 vssd1 vccd1 vccd1 _4772_/C sky130_fd_sc_hd__or2_1
XFILLER_0_96_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3967__A2 _3724_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__4916__A1 _4104_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4323__S _4327_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold596_A _6241_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4559__A _4575_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 _5304_/X vssd1 vssd1 vccd1 vccd1 _6151_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _5893_/Q vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4993__S _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5580__A1 _6159_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4383__A2 _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_A clkbuf_leaf_9_wb_clk_i/A vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3490_ _6299_/A _3525_/C _3473_/X vssd1 vssd1 vccd1 vccd1 _3491_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5064__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5160_ _5160_/A _5160_/B vssd1 vssd1 vccd1 vccd1 _5160_/X sky130_fd_sc_hd__or2_1
XFILLER_0_75_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4111_ hold163/X _3836_/X _4115_/S vssd1 vssd1 vccd1 vccd1 _4111_/X sky130_fd_sc_hd__mux2_1
X_5091_ _4737_/A _4124_/B _3143_/Y _4383_/Y _4433_/B vssd1 vssd1 vccd1 vccd1 _5091_/X
+ sky130_fd_sc_hd__a32o_1
X_4042_ _4094_/B _4416_/A _4416_/B _4750_/B vssd1 vssd1 vccd1 vccd1 _4048_/A sky130_fd_sc_hd__or4_2
XFILLER_0_91_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5993_ _6006_/CLK _5993_/D vssd1 vssd1 vccd1 vccd1 _5993_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4944_ _6239_/Q _5008_/B vssd1 vssd1 vccd1 vccd1 _4944_/X sky130_fd_sc_hd__and2_1
XFILLER_0_74_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4071__A1 _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4875_ _4874_/X _6060_/Q _5595_/S vssd1 vssd1 vccd1 vccd1 _4875_/X sky130_fd_sc_hd__mux2_1
XANTENNA__3548__A _4061_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3826_ _3656_/Y _3646_/X _3827_/B vssd1 vssd1 vccd1 vccd1 _3826_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3757_ _4234_/A _3757_/B vssd1 vssd1 vccd1 vccd1 _5052_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3688_ _5024_/B _3682_/Y _3687_/A _3639_/X vssd1 vssd1 vccd1 vccd1 _3688_/X sky130_fd_sc_hd__a22o_1
X_5427_ _5425_/X _5426_/Y _5326_/X vssd1 vssd1 vccd1 vccd1 _5427_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__5323__A1 _3539_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5323__B2 _4497_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5358_ hold478/X _5773_/B _5355_/X _5457_/A vssd1 vssd1 vccd1 vccd1 _5358_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_10_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5874__A2 _4415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4309_ _4261_/X hold250/X _4309_/S vssd1 vssd1 vccd1 vccd1 _4309_/X sky130_fd_sc_hd__mux2_1
XANTENNA__4509__S0 _5076_/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5289_ _3990_/B _4250_/B _5289_/S vssd1 vssd1 vccd1 vccd1 _5289_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_97_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4318__S _4318_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5657__B _5685_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__5612__S _5672_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5173__S0 _5185_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2990_ _2990_/A vssd1 vssd1 vccd1 vccd1 _2990_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_61_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__3368__A _4765_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5002__B1 _5607_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4660_ _4658_/Y _4676_/B vssd1 vssd1 vccd1 vccd1 _4662_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__4898__S _6038_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3611_ _3968_/A _3616_/B _3793_/D vssd1 vssd1 vccd1 vccd1 _3611_/X sky130_fd_sc_hd__and3_4
X_4591_ _4699_/A _4591_/B vssd1 vssd1 vccd1 vccd1 _4592_/B sky130_fd_sc_hd__or2_1
XFILLER_0_101_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3542_ _5093_/A _3542_/B vssd1 vssd1 vccd1 vccd1 _5078_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_3473_ hold588/X _3472_/X _3466_/Y _6299_/A vssd1 vssd1 vccd1 vccd1 _3473_/X sky130_fd_sc_hd__o211a_1
X_5212_ _6161_/Q _5121_/Y _5129_/Y _6219_/Q _5206_/X vssd1 vssd1 vccd1 vccd1 _5212_/X
+ sky130_fd_sc_hd__a221o_1
X_6192_ _6192_/CLK _6192_/D fanout177/X vssd1 vssd1 vccd1 vccd1 _6192_/Q sky130_fd_sc_hd__dfrtp_4
X_5143_ _5922_/Q _5200_/A2 _5200_/B1 _6030_/Q _5182_/S vssd1 vssd1 vccd1 vccd1 _5144_/C
+ sky130_fd_sc_hd__o221a_1
X_5074_ hold25/X _4250_/B _5772_/S vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__mux2_1
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4025_ _3655_/B _4020_/Y _4021_/X _5394_/B _3920_/A vssd1 vssd1 vccd1 vccd1 _4025_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5976_ _6038_/CLK hold45/X fanout170/X vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4927_ hold357/X _4926_/X _4927_/S vssd1 vssd1 vccd1 vccd1 _4927_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__4595__A2 _4612_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4858_ _6159_/Q _5008_/B _4853_/X _4999_/A1 _4856_/Y vssd1 vssd1 vccd1 vccd1 _4858_/X
+ sky130_fd_sc_hd__a221o_1
X_3809_ _3809_/A _3809_/B vssd1 vssd1 vccd1 vccd1 _3811_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_7_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4789_ _4990_/A _4789_/B vssd1 vssd1 vccd1 vccd1 _4789_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5480__A0 _6179_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5535__A1 _6156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3651__A _6073_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__3370__B _3370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3482__C1 _4094_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5830_ hold361/X _5794_/Y _5829_/X _5794_/B vssd1 vssd1 vccd1 vccd1 _5830_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_76_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5761_ _5767_/B _5762_/C vssd1 vssd1 vccd1 vccd1 _5761_/Y sky130_fd_sc_hd__nand2b_1
X_2973_ _6073_/Q vssd1 vssd1 vccd1 vccd1 _5025_/A sky130_fd_sc_hd__inv_2
X_4712_ _6027_/Q _5972_/Q _6019_/Q _5952_/Q _4712_/S0 _4712_/S1 vssd1 vssd1 vccd1
+ vccd1 _4712_/X sky130_fd_sc_hd__mux4_1
XFILLER_0_17_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5692_ _6186_/Q _6202_/Q _5701_/S vssd1 vssd1 vccd1 vccd1 _5692_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4643_ _4699_/A _4643_/B vssd1 vssd1 vccd1 vccd1 _4644_/B sky130_fd_sc_hd__or2_1
XFILLER_0_71_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4574_ _6210_/Q _4865_/B _4589_/S vssd1 vssd1 vccd1 vccd1 _4575_/C sky130_fd_sc_hd__mux2_1
XFILLER_0_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3525_ _3715_/B _6299_/A _3525_/C vssd1 vssd1 vccd1 vccd1 _5953_/D sky130_fd_sc_hd__or3_1
XFILLER_0_24_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_6244_ _6246_/CLK _6244_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6244_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3456_ _3453_/X _3455_/X _3441_/X vssd1 vssd1 vccd1 vccd1 _6299_/A sky130_fd_sc_hd__o21ai_4
X_6175_ _6175_/CLK _6175_/D fanout183/X vssd1 vssd1 vccd1 vccd1 _6175_/Q sky130_fd_sc_hd__dfstp_1
X_3387_ _3446_/A _3405_/B _5313_/S vssd1 vssd1 vccd1 vccd1 _4457_/B sky130_fd_sc_hd__or3_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_5126_ _6154_/Q _5121_/Y _5123_/Y _5088_/Y _5125_/X vssd1 vssd1 vccd1 vccd1 _5126_/X
+ sky130_fd_sc_hd__a221o_1
X_5057_ _5426_/A _5051_/A _5056_/X vssd1 vssd1 vccd1 vccd1 _5057_/X sky130_fd_sc_hd__a21bo_1
X_4008_ _4008_/A _4008_/B vssd1 vssd1 vccd1 vccd1 _4008_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3473__C1 _6299_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5765__A1 _5762_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5959_ _6006_/CLK _5959_/D vssd1 vssd1 vccd1 vccd1 _5959_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5517__A1 _4119_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4331__S _4336_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__4740__A2 _4759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__6051__RESET_B fanout172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_45_wb_clk_i clkbuf_2_2__f_wb_clk_i/X vssd1 vssd1 vccd1 vccd1 _6167_/CLK
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__5756__A1 _3864_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4964__C1 _4999_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5508__A1 _5507_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _4124_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3310_ _3192_/B _4731_/S _3446_/A vssd1 vssd1 vccd1 vccd1 _3320_/B sky130_fd_sc_hd__o21a_2
X_4290_ _4242_/X hold282/X _4291_/S vssd1 vssd1 vccd1 vccd1 _5951_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5072__S _5772_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3241_ _5356_/A _3643_/A _6174_/Q _3777_/A vssd1 vssd1 vccd1 vccd1 _3241_/X sky130_fd_sc_hd__and4b_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3172_ _3411_/B _3172_/B vssd1 vssd1 vccd1 vccd1 _3479_/B sky130_fd_sc_hd__or2_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5813_ _6240_/Q _5352_/A _5457_/A hold448/X vssd1 vssd1 vccd1 vccd1 _5813_/X sky130_fd_sc_hd__a2bb2o_1
XANTENNA__5747__A1 _3707_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4940__A _6156_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5744_ _3664_/X _5771_/S _5742_/Y _5743_/X vssd1 vssd1 vccd1 vccd1 _5744_/X sky130_fd_sc_hd__o22a_1
XFILLER_0_57_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2956_ _5507_/A vssd1 vssd1 vccd1 vccd1 _5480_/S sky130_fd_sc_hd__inv_2
XANTENNA__3222__A2 _6127_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5675_ _5694_/A _5674_/X _4976_/Y vssd1 vssd1 vccd1 vccd1 _5675_/X sky130_fd_sc_hd__a21bo_1
XANTENNA__4970__A2 _4815_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4626_ _4625_/X _4624_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4915_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_4_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3556__A _3556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold510 _6067_/Q vssd1 vssd1 vccd1 vccd1 hold510/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold521 _4653_/X vssd1 vssd1 vccd1 vccd1 _6064_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 _6219_/Q vssd1 vssd1 vccd1 vccd1 hold554/X sky130_fd_sc_hd__buf_1
XANTENNA__4722__A2 _4620_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold532 _6047_/Q vssd1 vssd1 vccd1 vccd1 _5314_/A sky130_fd_sc_hd__buf_2
X_4557_ _4556_/X _4555_/X _4697_/S vssd1 vssd1 vccd1 vccd1 _4850_/B sky130_fd_sc_hd__mux2_2
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold543 _4521_/X vssd1 vssd1 vccd1 vccd1 _6056_/D sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 _6216_/Q vssd1 vssd1 vccd1 vccd1 hold565/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold576 _6177_/Q vssd1 vssd1 vccd1 vccd1 hold576/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold587 _5238_/X vssd1 vssd1 vccd1 vccd1 _6130_/D sky130_fd_sc_hd__dlygate4sd3_1
X_3508_ _3508_/A _6121_/Q _3508_/C vssd1 vssd1 vccd1 vccd1 _3508_/X sky130_fd_sc_hd__and3_1
X_4488_ _5875_/B _4761_/A vssd1 vssd1 vccd1 vccd1 _4564_/S sky130_fd_sc_hd__nand2_2
Xhold598 _6236_/Q vssd1 vssd1 vccd1 vccd1 hold598/X sky130_fd_sc_hd__dlygate4sd3_1
X_6227_ _6227_/CLK _6227_/D fanout182/X vssd1 vssd1 vccd1 vccd1 _6227_/Q sky130_fd_sc_hd__dfstp_1
XANTENNA__5132__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3439_ _4737_/A _3439_/B vssd1 vssd1 vccd1 vccd1 _3439_/Y sky130_fd_sc_hd__nor2_1
X_6158_ _6238_/CLK _6158_/D fanout179/X vssd1 vssd1 vccd1 vccd1 _6158_/Q sky130_fd_sc_hd__dfrtp_4
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _5120_/A _5107_/A _5085_/B vssd1 vssd1 vccd1 vccd1 _5109_/Y sky130_fd_sc_hd__a21oi_4
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_6089_ _6251_/CLK _6089_/D fanout181/X vssd1 vssd1 vccd1 vccd1 _6089_/Q sky130_fd_sc_hd__dfrtp_2
XANTENNA__4326__S _4327_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__5199__C1 _4256_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__5738__A1 _4030_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__4850__A _4990_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput41 _6247_/Q vssd1 vssd1 vccd1 vccd1 io_out[27] sky130_fd_sc_hd__buf_12
Xoutput30 _6087_/Q vssd1 vssd1 vccd1 vccd1 io_out[17] sky130_fd_sc_hd__buf_12
Xoutput52 _6079_/Q vssd1 vssd1 vccd1 vccd1 io_out[9] sky130_fd_sc_hd__buf_12
XFILLER_0_101_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4477__A1 _4478_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__4572__S1 _4272_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__5729__A1 _3864_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__3835__S0 _5179_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3790_ hold240/X _3789_/X _4035_/S vssd1 vssd1 vccd1 vccd1 _5894_/D sky130_fd_sc_hd__mux2_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__5067__S _5073_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_5460_ _6118_/Q _5373_/B _5460_/S vssd1 vssd1 vccd1 vccd1 _5460_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_4411_ _5317_/A _4409_/X _4410_/Y _5327_/B _5773_/A vssd1 vssd1 vccd1 vccd1 _6043_/D
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5391_ _6173_/Q _3909_/B _4005_/A _5390_/Y vssd1 vssd1 vccd1 vccd1 _5392_/B sky130_fd_sc_hd__o211a_1
XFILLER_0_10_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__4919__B _5013_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4342_ hold199/X _3880_/X _4345_/S vssd1 vssd1 vccd1 vccd1 _4342_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4273_ _3405_/B _4771_/C _4121_/X _4272_/X vssd1 vssd1 vccd1 vccd1 _5936_/D sky130_fd_sc_hd__o31a_1
X_6012_ _6030_/CLK _6012_/D vssd1 vssd1 vccd1 vccd1 _6012_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__4000__A _5046_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3224_ _3323_/C _3223_/X _3249_/A vssd1 vssd1 vccd1 vccd1 _3224_/X sky130_fd_sc_hd__a21o_1
.ends

