magic
tech sky130B
magscale 1 2
timestamp 1717343180
<< obsli1 >>
rect 1104 2159 38824 217617
<< obsm1 >>
rect 106 2128 39914 217648
<< metal2 >>
rect 2042 219200 2098 220000
rect 2962 219200 3018 220000
rect 3882 219200 3938 220000
rect 4802 219200 4858 220000
rect 5722 219200 5778 220000
rect 6642 219200 6698 220000
rect 7562 219200 7618 220000
rect 8482 219200 8538 220000
rect 9402 219200 9458 220000
rect 10322 219200 10378 220000
rect 11242 219200 11298 220000
rect 12162 219200 12218 220000
rect 13082 219200 13138 220000
rect 14002 219200 14058 220000
rect 14922 219200 14978 220000
rect 15842 219200 15898 220000
rect 16762 219200 16818 220000
rect 17682 219200 17738 220000
rect 18602 219200 18658 220000
rect 19522 219200 19578 220000
rect 20442 219200 20498 220000
rect 21362 219200 21418 220000
rect 22282 219200 22338 220000
rect 23202 219200 23258 220000
rect 24122 219200 24178 220000
rect 25042 219200 25098 220000
rect 25962 219200 26018 220000
rect 26882 219200 26938 220000
rect 27802 219200 27858 220000
rect 28722 219200 28778 220000
rect 29642 219200 29698 220000
rect 30562 219200 30618 220000
rect 31482 219200 31538 220000
rect 32402 219200 32458 220000
rect 33322 219200 33378 220000
rect 34242 219200 34298 220000
rect 35162 219200 35218 220000
rect 36082 219200 36138 220000
rect 37002 219200 37058 220000
rect 37922 219200 37978 220000
rect 846 0 902 800
rect 2042 0 2098 800
rect 3238 0 3294 800
rect 4434 0 4490 800
rect 5630 0 5686 800
rect 6826 0 6882 800
rect 8022 0 8078 800
rect 9218 0 9274 800
rect 10414 0 10470 800
rect 11610 0 11666 800
rect 12806 0 12862 800
rect 14002 0 14058 800
rect 15198 0 15254 800
rect 16394 0 16450 800
rect 17590 0 17646 800
rect 18786 0 18842 800
rect 19982 0 20038 800
rect 21178 0 21234 800
rect 22374 0 22430 800
rect 23570 0 23626 800
rect 24766 0 24822 800
rect 25962 0 26018 800
rect 27158 0 27214 800
rect 28354 0 28410 800
rect 29550 0 29606 800
rect 30746 0 30802 800
rect 31942 0 31998 800
rect 33138 0 33194 800
rect 34334 0 34390 800
rect 35530 0 35586 800
rect 36726 0 36782 800
rect 37922 0 37978 800
rect 39118 0 39174 800
<< obsm2 >>
rect 110 219144 1986 219314
rect 2154 219144 2906 219314
rect 3074 219144 3826 219314
rect 3994 219144 4746 219314
rect 4914 219144 5666 219314
rect 5834 219144 6586 219314
rect 6754 219144 7506 219314
rect 7674 219144 8426 219314
rect 8594 219144 9346 219314
rect 9514 219144 10266 219314
rect 10434 219144 11186 219314
rect 11354 219144 12106 219314
rect 12274 219144 13026 219314
rect 13194 219144 13946 219314
rect 14114 219144 14866 219314
rect 15034 219144 15786 219314
rect 15954 219144 16706 219314
rect 16874 219144 17626 219314
rect 17794 219144 18546 219314
rect 18714 219144 19466 219314
rect 19634 219144 20386 219314
rect 20554 219144 21306 219314
rect 21474 219144 22226 219314
rect 22394 219144 23146 219314
rect 23314 219144 24066 219314
rect 24234 219144 24986 219314
rect 25154 219144 25906 219314
rect 26074 219144 26826 219314
rect 26994 219144 27746 219314
rect 27914 219144 28666 219314
rect 28834 219144 29586 219314
rect 29754 219144 30506 219314
rect 30674 219144 31426 219314
rect 31594 219144 32346 219314
rect 32514 219144 33266 219314
rect 33434 219144 34186 219314
rect 34354 219144 35106 219314
rect 35274 219144 36026 219314
rect 36194 219144 36946 219314
rect 37114 219144 37866 219314
rect 38034 219144 39988 219314
rect 110 856 39988 219144
rect 110 734 790 856
rect 958 734 1986 856
rect 2154 734 3182 856
rect 3350 734 4378 856
rect 4546 734 5574 856
rect 5742 734 6770 856
rect 6938 734 7966 856
rect 8134 734 9162 856
rect 9330 734 10358 856
rect 10526 734 11554 856
rect 11722 734 12750 856
rect 12918 734 13946 856
rect 14114 734 15142 856
rect 15310 734 16338 856
rect 16506 734 17534 856
rect 17702 734 18730 856
rect 18898 734 19926 856
rect 20094 734 21122 856
rect 21290 734 22318 856
rect 22486 734 23514 856
rect 23682 734 24710 856
rect 24878 734 25906 856
rect 26074 734 27102 856
rect 27270 734 28298 856
rect 28466 734 29494 856
rect 29662 734 30690 856
rect 30858 734 31886 856
rect 32054 734 33082 856
rect 33250 734 34278 856
rect 34446 734 35474 856
rect 35642 734 36670 856
rect 36838 734 37866 856
rect 38034 734 39062 856
rect 39230 734 39988 856
<< metal3 >>
rect 0 207272 800 207392
rect 0 206184 800 206304
rect 0 205096 800 205216
rect 0 204008 800 204128
rect 0 202920 800 203040
rect 0 201832 800 201952
rect 0 200744 800 200864
rect 0 199656 800 199776
rect 0 198568 800 198688
rect 0 197480 800 197600
rect 0 196392 800 196512
rect 0 195304 800 195424
rect 0 194216 800 194336
rect 0 193128 800 193248
rect 0 192040 800 192160
rect 0 190952 800 191072
rect 0 189864 800 189984
rect 39200 189320 40000 189440
rect 0 188776 800 188896
rect 39200 188776 40000 188896
rect 39200 188232 40000 188352
rect 0 187688 800 187808
rect 39200 187688 40000 187808
rect 39200 187144 40000 187264
rect 0 186600 800 186720
rect 39200 186600 40000 186720
rect 39200 186056 40000 186176
rect 0 185512 800 185632
rect 39200 185512 40000 185632
rect 39200 184968 40000 185088
rect 0 184424 800 184544
rect 39200 184424 40000 184544
rect 39200 183880 40000 184000
rect 0 183336 800 183456
rect 39200 183336 40000 183456
rect 39200 182792 40000 182912
rect 0 182248 800 182368
rect 39200 182248 40000 182368
rect 39200 181704 40000 181824
rect 0 181160 800 181280
rect 39200 181160 40000 181280
rect 39200 180616 40000 180736
rect 0 180072 800 180192
rect 39200 180072 40000 180192
rect 39200 179528 40000 179648
rect 0 178984 800 179104
rect 39200 178984 40000 179104
rect 39200 178440 40000 178560
rect 0 177896 800 178016
rect 39200 177896 40000 178016
rect 39200 177352 40000 177472
rect 0 176808 800 176928
rect 39200 176808 40000 176928
rect 39200 176264 40000 176384
rect 0 175720 800 175840
rect 39200 175720 40000 175840
rect 39200 175176 40000 175296
rect 0 174632 800 174752
rect 39200 174632 40000 174752
rect 39200 174088 40000 174208
rect 0 173544 800 173664
rect 39200 173544 40000 173664
rect 39200 173000 40000 173120
rect 0 172456 800 172576
rect 39200 172456 40000 172576
rect 39200 171912 40000 172032
rect 0 171368 800 171488
rect 39200 171368 40000 171488
rect 39200 170824 40000 170944
rect 0 170280 800 170400
rect 39200 170280 40000 170400
rect 39200 169736 40000 169856
rect 0 169192 800 169312
rect 39200 169192 40000 169312
rect 39200 168648 40000 168768
rect 0 168104 800 168224
rect 39200 168104 40000 168224
rect 39200 167560 40000 167680
rect 0 167016 800 167136
rect 39200 167016 40000 167136
rect 39200 166472 40000 166592
rect 0 165928 800 166048
rect 39200 165928 40000 166048
rect 39200 165384 40000 165504
rect 0 164840 800 164960
rect 39200 164840 40000 164960
rect 39200 164296 40000 164416
rect 0 163752 800 163872
rect 39200 163752 40000 163872
rect 39200 163208 40000 163328
rect 0 162664 800 162784
rect 39200 162664 40000 162784
rect 39200 162120 40000 162240
rect 0 161576 800 161696
rect 39200 161576 40000 161696
rect 39200 161032 40000 161152
rect 0 160488 800 160608
rect 39200 160488 40000 160608
rect 39200 159944 40000 160064
rect 0 159400 800 159520
rect 39200 159400 40000 159520
rect 39200 158856 40000 158976
rect 0 158312 800 158432
rect 39200 158312 40000 158432
rect 39200 157768 40000 157888
rect 0 157224 800 157344
rect 39200 157224 40000 157344
rect 39200 156680 40000 156800
rect 0 156136 800 156256
rect 39200 156136 40000 156256
rect 39200 155592 40000 155712
rect 0 155048 800 155168
rect 39200 155048 40000 155168
rect 39200 154504 40000 154624
rect 0 153960 800 154080
rect 39200 153960 40000 154080
rect 39200 153416 40000 153536
rect 0 152872 800 152992
rect 39200 152872 40000 152992
rect 39200 152328 40000 152448
rect 0 151784 800 151904
rect 39200 151784 40000 151904
rect 39200 151240 40000 151360
rect 0 150696 800 150816
rect 39200 150696 40000 150816
rect 39200 150152 40000 150272
rect 0 149608 800 149728
rect 39200 149608 40000 149728
rect 39200 149064 40000 149184
rect 0 148520 800 148640
rect 39200 148520 40000 148640
rect 39200 147976 40000 148096
rect 0 147432 800 147552
rect 39200 147432 40000 147552
rect 39200 146888 40000 147008
rect 0 146344 800 146464
rect 39200 146344 40000 146464
rect 39200 145800 40000 145920
rect 0 145256 800 145376
rect 39200 145256 40000 145376
rect 39200 144712 40000 144832
rect 0 144168 800 144288
rect 39200 144168 40000 144288
rect 39200 143624 40000 143744
rect 0 143080 800 143200
rect 39200 143080 40000 143200
rect 39200 142536 40000 142656
rect 0 141992 800 142112
rect 39200 141992 40000 142112
rect 39200 141448 40000 141568
rect 0 140904 800 141024
rect 39200 140904 40000 141024
rect 39200 140360 40000 140480
rect 0 139816 800 139936
rect 39200 139816 40000 139936
rect 39200 139272 40000 139392
rect 0 138728 800 138848
rect 39200 138728 40000 138848
rect 39200 138184 40000 138304
rect 0 137640 800 137760
rect 39200 137640 40000 137760
rect 39200 137096 40000 137216
rect 0 136552 800 136672
rect 39200 136552 40000 136672
rect 39200 136008 40000 136128
rect 0 135464 800 135584
rect 39200 135464 40000 135584
rect 39200 134920 40000 135040
rect 0 134376 800 134496
rect 39200 134376 40000 134496
rect 39200 133832 40000 133952
rect 0 133288 800 133408
rect 39200 133288 40000 133408
rect 39200 132744 40000 132864
rect 0 132200 800 132320
rect 39200 132200 40000 132320
rect 39200 131656 40000 131776
rect 0 131112 800 131232
rect 39200 131112 40000 131232
rect 39200 130568 40000 130688
rect 0 130024 800 130144
rect 39200 130024 40000 130144
rect 39200 129480 40000 129600
rect 0 128936 800 129056
rect 39200 128936 40000 129056
rect 39200 128392 40000 128512
rect 0 127848 800 127968
rect 39200 127848 40000 127968
rect 39200 127304 40000 127424
rect 0 126760 800 126880
rect 39200 126760 40000 126880
rect 39200 126216 40000 126336
rect 0 125672 800 125792
rect 39200 125672 40000 125792
rect 39200 125128 40000 125248
rect 0 124584 800 124704
rect 39200 124584 40000 124704
rect 39200 124040 40000 124160
rect 0 123496 800 123616
rect 39200 123496 40000 123616
rect 39200 122952 40000 123072
rect 0 122408 800 122528
rect 39200 122408 40000 122528
rect 39200 121864 40000 121984
rect 0 121320 800 121440
rect 39200 121320 40000 121440
rect 39200 120776 40000 120896
rect 0 120232 800 120352
rect 39200 120232 40000 120352
rect 39200 119688 40000 119808
rect 0 119144 800 119264
rect 39200 119144 40000 119264
rect 39200 118600 40000 118720
rect 0 118056 800 118176
rect 39200 118056 40000 118176
rect 39200 117512 40000 117632
rect 0 116968 800 117088
rect 39200 116968 40000 117088
rect 39200 116424 40000 116544
rect 0 115880 800 116000
rect 39200 115880 40000 116000
rect 39200 115336 40000 115456
rect 0 114792 800 114912
rect 39200 114792 40000 114912
rect 39200 114248 40000 114368
rect 0 113704 800 113824
rect 39200 113704 40000 113824
rect 39200 113160 40000 113280
rect 0 112616 800 112736
rect 39200 112616 40000 112736
rect 39200 112072 40000 112192
rect 0 111528 800 111648
rect 39200 111528 40000 111648
rect 39200 110984 40000 111104
rect 0 110440 800 110560
rect 39200 110440 40000 110560
rect 39200 109896 40000 110016
rect 0 109352 800 109472
rect 39200 109352 40000 109472
rect 39200 108808 40000 108928
rect 0 108264 800 108384
rect 39200 108264 40000 108384
rect 39200 107720 40000 107840
rect 0 107176 800 107296
rect 39200 107176 40000 107296
rect 39200 106632 40000 106752
rect 0 106088 800 106208
rect 39200 106088 40000 106208
rect 39200 105544 40000 105664
rect 0 105000 800 105120
rect 39200 105000 40000 105120
rect 39200 104456 40000 104576
rect 0 103912 800 104032
rect 39200 103912 40000 104032
rect 39200 103368 40000 103488
rect 0 102824 800 102944
rect 39200 102824 40000 102944
rect 39200 102280 40000 102400
rect 0 101736 800 101856
rect 39200 101736 40000 101856
rect 39200 101192 40000 101312
rect 0 100648 800 100768
rect 39200 100648 40000 100768
rect 39200 100104 40000 100224
rect 0 99560 800 99680
rect 39200 99560 40000 99680
rect 39200 99016 40000 99136
rect 0 98472 800 98592
rect 39200 98472 40000 98592
rect 39200 97928 40000 98048
rect 0 97384 800 97504
rect 39200 97384 40000 97504
rect 39200 96840 40000 96960
rect 0 96296 800 96416
rect 39200 96296 40000 96416
rect 39200 95752 40000 95872
rect 0 95208 800 95328
rect 39200 95208 40000 95328
rect 39200 94664 40000 94784
rect 0 94120 800 94240
rect 39200 94120 40000 94240
rect 39200 93576 40000 93696
rect 0 93032 800 93152
rect 39200 93032 40000 93152
rect 39200 92488 40000 92608
rect 0 91944 800 92064
rect 39200 91944 40000 92064
rect 39200 91400 40000 91520
rect 0 90856 800 90976
rect 39200 90856 40000 90976
rect 39200 90312 40000 90432
rect 0 89768 800 89888
rect 39200 89768 40000 89888
rect 39200 89224 40000 89344
rect 0 88680 800 88800
rect 39200 88680 40000 88800
rect 39200 88136 40000 88256
rect 0 87592 800 87712
rect 39200 87592 40000 87712
rect 39200 87048 40000 87168
rect 0 86504 800 86624
rect 39200 86504 40000 86624
rect 39200 85960 40000 86080
rect 0 85416 800 85536
rect 39200 85416 40000 85536
rect 39200 84872 40000 84992
rect 0 84328 800 84448
rect 39200 84328 40000 84448
rect 39200 83784 40000 83904
rect 0 83240 800 83360
rect 39200 83240 40000 83360
rect 39200 82696 40000 82816
rect 0 82152 800 82272
rect 39200 82152 40000 82272
rect 39200 81608 40000 81728
rect 0 81064 800 81184
rect 39200 81064 40000 81184
rect 39200 80520 40000 80640
rect 0 79976 800 80096
rect 39200 79976 40000 80096
rect 39200 79432 40000 79552
rect 0 78888 800 79008
rect 39200 78888 40000 79008
rect 39200 78344 40000 78464
rect 0 77800 800 77920
rect 39200 77800 40000 77920
rect 39200 77256 40000 77376
rect 0 76712 800 76832
rect 39200 76712 40000 76832
rect 39200 76168 40000 76288
rect 0 75624 800 75744
rect 39200 75624 40000 75744
rect 39200 75080 40000 75200
rect 0 74536 800 74656
rect 39200 74536 40000 74656
rect 39200 73992 40000 74112
rect 0 73448 800 73568
rect 39200 73448 40000 73568
rect 39200 72904 40000 73024
rect 0 72360 800 72480
rect 39200 72360 40000 72480
rect 39200 71816 40000 71936
rect 0 71272 800 71392
rect 39200 71272 40000 71392
rect 39200 70728 40000 70848
rect 0 70184 800 70304
rect 39200 70184 40000 70304
rect 39200 69640 40000 69760
rect 0 69096 800 69216
rect 39200 69096 40000 69216
rect 39200 68552 40000 68672
rect 0 68008 800 68128
rect 39200 68008 40000 68128
rect 39200 67464 40000 67584
rect 0 66920 800 67040
rect 39200 66920 40000 67040
rect 39200 66376 40000 66496
rect 0 65832 800 65952
rect 39200 65832 40000 65952
rect 39200 65288 40000 65408
rect 0 64744 800 64864
rect 39200 64744 40000 64864
rect 39200 64200 40000 64320
rect 0 63656 800 63776
rect 39200 63656 40000 63776
rect 39200 63112 40000 63232
rect 0 62568 800 62688
rect 39200 62568 40000 62688
rect 39200 62024 40000 62144
rect 0 61480 800 61600
rect 39200 61480 40000 61600
rect 39200 60936 40000 61056
rect 0 60392 800 60512
rect 39200 60392 40000 60512
rect 39200 59848 40000 59968
rect 0 59304 800 59424
rect 39200 59304 40000 59424
rect 39200 58760 40000 58880
rect 0 58216 800 58336
rect 39200 58216 40000 58336
rect 39200 57672 40000 57792
rect 0 57128 800 57248
rect 39200 57128 40000 57248
rect 39200 56584 40000 56704
rect 0 56040 800 56160
rect 39200 56040 40000 56160
rect 39200 55496 40000 55616
rect 0 54952 800 55072
rect 39200 54952 40000 55072
rect 39200 54408 40000 54528
rect 0 53864 800 53984
rect 39200 53864 40000 53984
rect 39200 53320 40000 53440
rect 0 52776 800 52896
rect 39200 52776 40000 52896
rect 39200 52232 40000 52352
rect 0 51688 800 51808
rect 39200 51688 40000 51808
rect 39200 51144 40000 51264
rect 0 50600 800 50720
rect 39200 50600 40000 50720
rect 39200 50056 40000 50176
rect 0 49512 800 49632
rect 39200 49512 40000 49632
rect 39200 48968 40000 49088
rect 0 48424 800 48544
rect 39200 48424 40000 48544
rect 39200 47880 40000 48000
rect 0 47336 800 47456
rect 39200 47336 40000 47456
rect 39200 46792 40000 46912
rect 0 46248 800 46368
rect 39200 46248 40000 46368
rect 39200 45704 40000 45824
rect 0 45160 800 45280
rect 39200 45160 40000 45280
rect 39200 44616 40000 44736
rect 0 44072 800 44192
rect 39200 44072 40000 44192
rect 39200 43528 40000 43648
rect 0 42984 800 43104
rect 39200 42984 40000 43104
rect 39200 42440 40000 42560
rect 0 41896 800 42016
rect 39200 41896 40000 42016
rect 39200 41352 40000 41472
rect 0 40808 800 40928
rect 39200 40808 40000 40928
rect 39200 40264 40000 40384
rect 0 39720 800 39840
rect 39200 39720 40000 39840
rect 39200 39176 40000 39296
rect 0 38632 800 38752
rect 39200 38632 40000 38752
rect 39200 38088 40000 38208
rect 0 37544 800 37664
rect 39200 37544 40000 37664
rect 39200 37000 40000 37120
rect 0 36456 800 36576
rect 39200 36456 40000 36576
rect 39200 35912 40000 36032
rect 0 35368 800 35488
rect 39200 35368 40000 35488
rect 39200 34824 40000 34944
rect 0 34280 800 34400
rect 39200 34280 40000 34400
rect 39200 33736 40000 33856
rect 0 33192 800 33312
rect 39200 33192 40000 33312
rect 39200 32648 40000 32768
rect 0 32104 800 32224
rect 39200 32104 40000 32224
rect 39200 31560 40000 31680
rect 0 31016 800 31136
rect 39200 31016 40000 31136
rect 39200 30472 40000 30592
rect 0 29928 800 30048
rect 0 28840 800 28960
rect 0 27752 800 27872
rect 0 26664 800 26784
rect 0 25576 800 25696
rect 0 24488 800 24608
rect 0 23400 800 23520
rect 0 22312 800 22432
rect 0 21224 800 21344
rect 0 20136 800 20256
rect 0 19048 800 19168
rect 0 17960 800 18080
rect 0 16872 800 16992
rect 0 15784 800 15904
rect 0 14696 800 14816
rect 0 13608 800 13728
rect 0 12520 800 12640
<< obsm3 >>
rect 105 207472 39915 217633
rect 880 207192 39915 207472
rect 105 206384 39915 207192
rect 880 206104 39915 206384
rect 105 205296 39915 206104
rect 880 205016 39915 205296
rect 105 204208 39915 205016
rect 880 203928 39915 204208
rect 105 203120 39915 203928
rect 880 202840 39915 203120
rect 105 202032 39915 202840
rect 880 201752 39915 202032
rect 105 200944 39915 201752
rect 880 200664 39915 200944
rect 105 199856 39915 200664
rect 880 199576 39915 199856
rect 105 198768 39915 199576
rect 880 198488 39915 198768
rect 105 197680 39915 198488
rect 880 197400 39915 197680
rect 105 196592 39915 197400
rect 880 196312 39915 196592
rect 105 195504 39915 196312
rect 880 195224 39915 195504
rect 105 194416 39915 195224
rect 880 194136 39915 194416
rect 105 193328 39915 194136
rect 880 193048 39915 193328
rect 105 192240 39915 193048
rect 880 191960 39915 192240
rect 105 191152 39915 191960
rect 880 190872 39915 191152
rect 105 190064 39915 190872
rect 880 189784 39915 190064
rect 105 189520 39915 189784
rect 105 189240 39120 189520
rect 105 188976 39915 189240
rect 880 188696 39120 188976
rect 105 188432 39915 188696
rect 105 188152 39120 188432
rect 105 187888 39915 188152
rect 880 187608 39120 187888
rect 105 187344 39915 187608
rect 105 187064 39120 187344
rect 105 186800 39915 187064
rect 880 186520 39120 186800
rect 105 186256 39915 186520
rect 105 185976 39120 186256
rect 105 185712 39915 185976
rect 880 185432 39120 185712
rect 105 185168 39915 185432
rect 105 184888 39120 185168
rect 105 184624 39915 184888
rect 880 184344 39120 184624
rect 105 184080 39915 184344
rect 105 183800 39120 184080
rect 105 183536 39915 183800
rect 880 183256 39120 183536
rect 105 182992 39915 183256
rect 105 182712 39120 182992
rect 105 182448 39915 182712
rect 880 182168 39120 182448
rect 105 181904 39915 182168
rect 105 181624 39120 181904
rect 105 181360 39915 181624
rect 880 181080 39120 181360
rect 105 180816 39915 181080
rect 105 180536 39120 180816
rect 105 180272 39915 180536
rect 880 179992 39120 180272
rect 105 179728 39915 179992
rect 105 179448 39120 179728
rect 105 179184 39915 179448
rect 880 178904 39120 179184
rect 105 178640 39915 178904
rect 105 178360 39120 178640
rect 105 178096 39915 178360
rect 880 177816 39120 178096
rect 105 177552 39915 177816
rect 105 177272 39120 177552
rect 105 177008 39915 177272
rect 880 176728 39120 177008
rect 105 176464 39915 176728
rect 105 176184 39120 176464
rect 105 175920 39915 176184
rect 880 175640 39120 175920
rect 105 175376 39915 175640
rect 105 175096 39120 175376
rect 105 174832 39915 175096
rect 880 174552 39120 174832
rect 105 174288 39915 174552
rect 105 174008 39120 174288
rect 105 173744 39915 174008
rect 880 173464 39120 173744
rect 105 173200 39915 173464
rect 105 172920 39120 173200
rect 105 172656 39915 172920
rect 880 172376 39120 172656
rect 105 172112 39915 172376
rect 105 171832 39120 172112
rect 105 171568 39915 171832
rect 880 171288 39120 171568
rect 105 171024 39915 171288
rect 105 170744 39120 171024
rect 105 170480 39915 170744
rect 880 170200 39120 170480
rect 105 169936 39915 170200
rect 105 169656 39120 169936
rect 105 169392 39915 169656
rect 880 169112 39120 169392
rect 105 168848 39915 169112
rect 105 168568 39120 168848
rect 105 168304 39915 168568
rect 880 168024 39120 168304
rect 105 167760 39915 168024
rect 105 167480 39120 167760
rect 105 167216 39915 167480
rect 880 166936 39120 167216
rect 105 166672 39915 166936
rect 105 166392 39120 166672
rect 105 166128 39915 166392
rect 880 165848 39120 166128
rect 105 165584 39915 165848
rect 105 165304 39120 165584
rect 105 165040 39915 165304
rect 880 164760 39120 165040
rect 105 164496 39915 164760
rect 105 164216 39120 164496
rect 105 163952 39915 164216
rect 880 163672 39120 163952
rect 105 163408 39915 163672
rect 105 163128 39120 163408
rect 105 162864 39915 163128
rect 880 162584 39120 162864
rect 105 162320 39915 162584
rect 105 162040 39120 162320
rect 105 161776 39915 162040
rect 880 161496 39120 161776
rect 105 161232 39915 161496
rect 105 160952 39120 161232
rect 105 160688 39915 160952
rect 880 160408 39120 160688
rect 105 160144 39915 160408
rect 105 159864 39120 160144
rect 105 159600 39915 159864
rect 880 159320 39120 159600
rect 105 159056 39915 159320
rect 105 158776 39120 159056
rect 105 158512 39915 158776
rect 880 158232 39120 158512
rect 105 157968 39915 158232
rect 105 157688 39120 157968
rect 105 157424 39915 157688
rect 880 157144 39120 157424
rect 105 156880 39915 157144
rect 105 156600 39120 156880
rect 105 156336 39915 156600
rect 880 156056 39120 156336
rect 105 155792 39915 156056
rect 105 155512 39120 155792
rect 105 155248 39915 155512
rect 880 154968 39120 155248
rect 105 154704 39915 154968
rect 105 154424 39120 154704
rect 105 154160 39915 154424
rect 880 153880 39120 154160
rect 105 153616 39915 153880
rect 105 153336 39120 153616
rect 105 153072 39915 153336
rect 880 152792 39120 153072
rect 105 152528 39915 152792
rect 105 152248 39120 152528
rect 105 151984 39915 152248
rect 880 151704 39120 151984
rect 105 151440 39915 151704
rect 105 151160 39120 151440
rect 105 150896 39915 151160
rect 880 150616 39120 150896
rect 105 150352 39915 150616
rect 105 150072 39120 150352
rect 105 149808 39915 150072
rect 880 149528 39120 149808
rect 105 149264 39915 149528
rect 105 148984 39120 149264
rect 105 148720 39915 148984
rect 880 148440 39120 148720
rect 105 148176 39915 148440
rect 105 147896 39120 148176
rect 105 147632 39915 147896
rect 880 147352 39120 147632
rect 105 147088 39915 147352
rect 105 146808 39120 147088
rect 105 146544 39915 146808
rect 880 146264 39120 146544
rect 105 146000 39915 146264
rect 105 145720 39120 146000
rect 105 145456 39915 145720
rect 880 145176 39120 145456
rect 105 144912 39915 145176
rect 105 144632 39120 144912
rect 105 144368 39915 144632
rect 880 144088 39120 144368
rect 105 143824 39915 144088
rect 105 143544 39120 143824
rect 105 143280 39915 143544
rect 880 143000 39120 143280
rect 105 142736 39915 143000
rect 105 142456 39120 142736
rect 105 142192 39915 142456
rect 880 141912 39120 142192
rect 105 141648 39915 141912
rect 105 141368 39120 141648
rect 105 141104 39915 141368
rect 880 140824 39120 141104
rect 105 140560 39915 140824
rect 105 140280 39120 140560
rect 105 140016 39915 140280
rect 880 139736 39120 140016
rect 105 139472 39915 139736
rect 105 139192 39120 139472
rect 105 138928 39915 139192
rect 880 138648 39120 138928
rect 105 138384 39915 138648
rect 105 138104 39120 138384
rect 105 137840 39915 138104
rect 880 137560 39120 137840
rect 105 137296 39915 137560
rect 105 137016 39120 137296
rect 105 136752 39915 137016
rect 880 136472 39120 136752
rect 105 136208 39915 136472
rect 105 135928 39120 136208
rect 105 135664 39915 135928
rect 880 135384 39120 135664
rect 105 135120 39915 135384
rect 105 134840 39120 135120
rect 105 134576 39915 134840
rect 880 134296 39120 134576
rect 105 134032 39915 134296
rect 105 133752 39120 134032
rect 105 133488 39915 133752
rect 880 133208 39120 133488
rect 105 132944 39915 133208
rect 105 132664 39120 132944
rect 105 132400 39915 132664
rect 880 132120 39120 132400
rect 105 131856 39915 132120
rect 105 131576 39120 131856
rect 105 131312 39915 131576
rect 880 131032 39120 131312
rect 105 130768 39915 131032
rect 105 130488 39120 130768
rect 105 130224 39915 130488
rect 880 129944 39120 130224
rect 105 129680 39915 129944
rect 105 129400 39120 129680
rect 105 129136 39915 129400
rect 880 128856 39120 129136
rect 105 128592 39915 128856
rect 105 128312 39120 128592
rect 105 128048 39915 128312
rect 880 127768 39120 128048
rect 105 127504 39915 127768
rect 105 127224 39120 127504
rect 105 126960 39915 127224
rect 880 126680 39120 126960
rect 105 126416 39915 126680
rect 105 126136 39120 126416
rect 105 125872 39915 126136
rect 880 125592 39120 125872
rect 105 125328 39915 125592
rect 105 125048 39120 125328
rect 105 124784 39915 125048
rect 880 124504 39120 124784
rect 105 124240 39915 124504
rect 105 123960 39120 124240
rect 105 123696 39915 123960
rect 880 123416 39120 123696
rect 105 123152 39915 123416
rect 105 122872 39120 123152
rect 105 122608 39915 122872
rect 880 122328 39120 122608
rect 105 122064 39915 122328
rect 105 121784 39120 122064
rect 105 121520 39915 121784
rect 880 121240 39120 121520
rect 105 120976 39915 121240
rect 105 120696 39120 120976
rect 105 120432 39915 120696
rect 880 120152 39120 120432
rect 105 119888 39915 120152
rect 105 119608 39120 119888
rect 105 119344 39915 119608
rect 880 119064 39120 119344
rect 105 118800 39915 119064
rect 105 118520 39120 118800
rect 105 118256 39915 118520
rect 880 117976 39120 118256
rect 105 117712 39915 117976
rect 105 117432 39120 117712
rect 105 117168 39915 117432
rect 880 116888 39120 117168
rect 105 116624 39915 116888
rect 105 116344 39120 116624
rect 105 116080 39915 116344
rect 880 115800 39120 116080
rect 105 115536 39915 115800
rect 105 115256 39120 115536
rect 105 114992 39915 115256
rect 880 114712 39120 114992
rect 105 114448 39915 114712
rect 105 114168 39120 114448
rect 105 113904 39915 114168
rect 880 113624 39120 113904
rect 105 113360 39915 113624
rect 105 113080 39120 113360
rect 105 112816 39915 113080
rect 880 112536 39120 112816
rect 105 112272 39915 112536
rect 105 111992 39120 112272
rect 105 111728 39915 111992
rect 880 111448 39120 111728
rect 105 111184 39915 111448
rect 105 110904 39120 111184
rect 105 110640 39915 110904
rect 880 110360 39120 110640
rect 105 110096 39915 110360
rect 105 109816 39120 110096
rect 105 109552 39915 109816
rect 880 109272 39120 109552
rect 105 109008 39915 109272
rect 105 108728 39120 109008
rect 105 108464 39915 108728
rect 880 108184 39120 108464
rect 105 107920 39915 108184
rect 105 107640 39120 107920
rect 105 107376 39915 107640
rect 880 107096 39120 107376
rect 105 106832 39915 107096
rect 105 106552 39120 106832
rect 105 106288 39915 106552
rect 880 106008 39120 106288
rect 105 105744 39915 106008
rect 105 105464 39120 105744
rect 105 105200 39915 105464
rect 880 104920 39120 105200
rect 105 104656 39915 104920
rect 105 104376 39120 104656
rect 105 104112 39915 104376
rect 880 103832 39120 104112
rect 105 103568 39915 103832
rect 105 103288 39120 103568
rect 105 103024 39915 103288
rect 880 102744 39120 103024
rect 105 102480 39915 102744
rect 105 102200 39120 102480
rect 105 101936 39915 102200
rect 880 101656 39120 101936
rect 105 101392 39915 101656
rect 105 101112 39120 101392
rect 105 100848 39915 101112
rect 880 100568 39120 100848
rect 105 100304 39915 100568
rect 105 100024 39120 100304
rect 105 99760 39915 100024
rect 880 99480 39120 99760
rect 105 99216 39915 99480
rect 105 98936 39120 99216
rect 105 98672 39915 98936
rect 880 98392 39120 98672
rect 105 98128 39915 98392
rect 105 97848 39120 98128
rect 105 97584 39915 97848
rect 880 97304 39120 97584
rect 105 97040 39915 97304
rect 105 96760 39120 97040
rect 105 96496 39915 96760
rect 880 96216 39120 96496
rect 105 95952 39915 96216
rect 105 95672 39120 95952
rect 105 95408 39915 95672
rect 880 95128 39120 95408
rect 105 94864 39915 95128
rect 105 94584 39120 94864
rect 105 94320 39915 94584
rect 880 94040 39120 94320
rect 105 93776 39915 94040
rect 105 93496 39120 93776
rect 105 93232 39915 93496
rect 880 92952 39120 93232
rect 105 92688 39915 92952
rect 105 92408 39120 92688
rect 105 92144 39915 92408
rect 880 91864 39120 92144
rect 105 91600 39915 91864
rect 105 91320 39120 91600
rect 105 91056 39915 91320
rect 880 90776 39120 91056
rect 105 90512 39915 90776
rect 105 90232 39120 90512
rect 105 89968 39915 90232
rect 880 89688 39120 89968
rect 105 89424 39915 89688
rect 105 89144 39120 89424
rect 105 88880 39915 89144
rect 880 88600 39120 88880
rect 105 88336 39915 88600
rect 105 88056 39120 88336
rect 105 87792 39915 88056
rect 880 87512 39120 87792
rect 105 87248 39915 87512
rect 105 86968 39120 87248
rect 105 86704 39915 86968
rect 880 86424 39120 86704
rect 105 86160 39915 86424
rect 105 85880 39120 86160
rect 105 85616 39915 85880
rect 880 85336 39120 85616
rect 105 85072 39915 85336
rect 105 84792 39120 85072
rect 105 84528 39915 84792
rect 880 84248 39120 84528
rect 105 83984 39915 84248
rect 105 83704 39120 83984
rect 105 83440 39915 83704
rect 880 83160 39120 83440
rect 105 82896 39915 83160
rect 105 82616 39120 82896
rect 105 82352 39915 82616
rect 880 82072 39120 82352
rect 105 81808 39915 82072
rect 105 81528 39120 81808
rect 105 81264 39915 81528
rect 880 80984 39120 81264
rect 105 80720 39915 80984
rect 105 80440 39120 80720
rect 105 80176 39915 80440
rect 880 79896 39120 80176
rect 105 79632 39915 79896
rect 105 79352 39120 79632
rect 105 79088 39915 79352
rect 880 78808 39120 79088
rect 105 78544 39915 78808
rect 105 78264 39120 78544
rect 105 78000 39915 78264
rect 880 77720 39120 78000
rect 105 77456 39915 77720
rect 105 77176 39120 77456
rect 105 76912 39915 77176
rect 880 76632 39120 76912
rect 105 76368 39915 76632
rect 105 76088 39120 76368
rect 105 75824 39915 76088
rect 880 75544 39120 75824
rect 105 75280 39915 75544
rect 105 75000 39120 75280
rect 105 74736 39915 75000
rect 880 74456 39120 74736
rect 105 74192 39915 74456
rect 105 73912 39120 74192
rect 105 73648 39915 73912
rect 880 73368 39120 73648
rect 105 73104 39915 73368
rect 105 72824 39120 73104
rect 105 72560 39915 72824
rect 880 72280 39120 72560
rect 105 72016 39915 72280
rect 105 71736 39120 72016
rect 105 71472 39915 71736
rect 880 71192 39120 71472
rect 105 70928 39915 71192
rect 105 70648 39120 70928
rect 105 70384 39915 70648
rect 880 70104 39120 70384
rect 105 69840 39915 70104
rect 105 69560 39120 69840
rect 105 69296 39915 69560
rect 880 69016 39120 69296
rect 105 68752 39915 69016
rect 105 68472 39120 68752
rect 105 68208 39915 68472
rect 880 67928 39120 68208
rect 105 67664 39915 67928
rect 105 67384 39120 67664
rect 105 67120 39915 67384
rect 880 66840 39120 67120
rect 105 66576 39915 66840
rect 105 66296 39120 66576
rect 105 66032 39915 66296
rect 880 65752 39120 66032
rect 105 65488 39915 65752
rect 105 65208 39120 65488
rect 105 64944 39915 65208
rect 880 64664 39120 64944
rect 105 64400 39915 64664
rect 105 64120 39120 64400
rect 105 63856 39915 64120
rect 880 63576 39120 63856
rect 105 63312 39915 63576
rect 105 63032 39120 63312
rect 105 62768 39915 63032
rect 880 62488 39120 62768
rect 105 62224 39915 62488
rect 105 61944 39120 62224
rect 105 61680 39915 61944
rect 880 61400 39120 61680
rect 105 61136 39915 61400
rect 105 60856 39120 61136
rect 105 60592 39915 60856
rect 880 60312 39120 60592
rect 105 60048 39915 60312
rect 105 59768 39120 60048
rect 105 59504 39915 59768
rect 880 59224 39120 59504
rect 105 58960 39915 59224
rect 105 58680 39120 58960
rect 105 58416 39915 58680
rect 880 58136 39120 58416
rect 105 57872 39915 58136
rect 105 57592 39120 57872
rect 105 57328 39915 57592
rect 880 57048 39120 57328
rect 105 56784 39915 57048
rect 105 56504 39120 56784
rect 105 56240 39915 56504
rect 880 55960 39120 56240
rect 105 55696 39915 55960
rect 105 55416 39120 55696
rect 105 55152 39915 55416
rect 880 54872 39120 55152
rect 105 54608 39915 54872
rect 105 54328 39120 54608
rect 105 54064 39915 54328
rect 880 53784 39120 54064
rect 105 53520 39915 53784
rect 105 53240 39120 53520
rect 105 52976 39915 53240
rect 880 52696 39120 52976
rect 105 52432 39915 52696
rect 105 52152 39120 52432
rect 105 51888 39915 52152
rect 880 51608 39120 51888
rect 105 51344 39915 51608
rect 105 51064 39120 51344
rect 105 50800 39915 51064
rect 880 50520 39120 50800
rect 105 50256 39915 50520
rect 105 49976 39120 50256
rect 105 49712 39915 49976
rect 880 49432 39120 49712
rect 105 49168 39915 49432
rect 105 48888 39120 49168
rect 105 48624 39915 48888
rect 880 48344 39120 48624
rect 105 48080 39915 48344
rect 105 47800 39120 48080
rect 105 47536 39915 47800
rect 880 47256 39120 47536
rect 105 46992 39915 47256
rect 105 46712 39120 46992
rect 105 46448 39915 46712
rect 880 46168 39120 46448
rect 105 45904 39915 46168
rect 105 45624 39120 45904
rect 105 45360 39915 45624
rect 880 45080 39120 45360
rect 105 44816 39915 45080
rect 105 44536 39120 44816
rect 105 44272 39915 44536
rect 880 43992 39120 44272
rect 105 43728 39915 43992
rect 105 43448 39120 43728
rect 105 43184 39915 43448
rect 880 42904 39120 43184
rect 105 42640 39915 42904
rect 105 42360 39120 42640
rect 105 42096 39915 42360
rect 880 41816 39120 42096
rect 105 41552 39915 41816
rect 105 41272 39120 41552
rect 105 41008 39915 41272
rect 880 40728 39120 41008
rect 105 40464 39915 40728
rect 105 40184 39120 40464
rect 105 39920 39915 40184
rect 880 39640 39120 39920
rect 105 39376 39915 39640
rect 105 39096 39120 39376
rect 105 38832 39915 39096
rect 880 38552 39120 38832
rect 105 38288 39915 38552
rect 105 38008 39120 38288
rect 105 37744 39915 38008
rect 880 37464 39120 37744
rect 105 37200 39915 37464
rect 105 36920 39120 37200
rect 105 36656 39915 36920
rect 880 36376 39120 36656
rect 105 36112 39915 36376
rect 105 35832 39120 36112
rect 105 35568 39915 35832
rect 880 35288 39120 35568
rect 105 35024 39915 35288
rect 105 34744 39120 35024
rect 105 34480 39915 34744
rect 880 34200 39120 34480
rect 105 33936 39915 34200
rect 105 33656 39120 33936
rect 105 33392 39915 33656
rect 880 33112 39120 33392
rect 105 32848 39915 33112
rect 105 32568 39120 32848
rect 105 32304 39915 32568
rect 880 32024 39120 32304
rect 105 31760 39915 32024
rect 105 31480 39120 31760
rect 105 31216 39915 31480
rect 880 30936 39120 31216
rect 105 30672 39915 30936
rect 105 30392 39120 30672
rect 105 30128 39915 30392
rect 880 29848 39915 30128
rect 105 29040 39915 29848
rect 880 28760 39915 29040
rect 105 27952 39915 28760
rect 880 27672 39915 27952
rect 105 26864 39915 27672
rect 880 26584 39915 26864
rect 105 25776 39915 26584
rect 880 25496 39915 25776
rect 105 24688 39915 25496
rect 880 24408 39915 24688
rect 105 23600 39915 24408
rect 880 23320 39915 23600
rect 105 22512 39915 23320
rect 880 22232 39915 22512
rect 105 21424 39915 22232
rect 880 21144 39915 21424
rect 105 20336 39915 21144
rect 880 20056 39915 20336
rect 105 19248 39915 20056
rect 880 18968 39915 19248
rect 105 18160 39915 18968
rect 880 17880 39915 18160
rect 105 17072 39915 17880
rect 880 16792 39915 17072
rect 105 15984 39915 16792
rect 880 15704 39915 15984
rect 105 14896 39915 15704
rect 880 14616 39915 14896
rect 105 13808 39915 14616
rect 880 13528 39915 13808
rect 105 12720 39915 13528
rect 880 12440 39915 12720
rect 105 2143 39915 12440
<< metal4 >>
rect 4208 2128 4528 217648
rect 19568 2128 19888 217648
rect 34928 2128 35248 217648
<< obsm4 >>
rect 427 14587 4128 214573
rect 4608 14587 19488 214573
rect 19968 14587 34848 214573
rect 35328 14587 39133 214573
<< labels >>
rlabel metal3 s 0 95208 800 95328 6 custom_settings[0]
port 1 nsew signal output
rlabel metal3 s 0 106088 800 106208 6 custom_settings[10]
port 2 nsew signal output
rlabel metal3 s 0 107176 800 107296 6 custom_settings[11]
port 3 nsew signal output
rlabel metal3 s 0 108264 800 108384 6 custom_settings[12]
port 4 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 custom_settings[13]
port 5 nsew signal output
rlabel metal3 s 0 110440 800 110560 6 custom_settings[14]
port 6 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 custom_settings[15]
port 7 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 custom_settings[16]
port 8 nsew signal output
rlabel metal3 s 0 113704 800 113824 6 custom_settings[17]
port 9 nsew signal output
rlabel metal3 s 0 114792 800 114912 6 custom_settings[18]
port 10 nsew signal output
rlabel metal3 s 0 115880 800 116000 6 custom_settings[19]
port 11 nsew signal output
rlabel metal3 s 0 96296 800 96416 6 custom_settings[1]
port 12 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 custom_settings[20]
port 13 nsew signal output
rlabel metal3 s 0 118056 800 118176 6 custom_settings[21]
port 14 nsew signal output
rlabel metal3 s 0 119144 800 119264 6 custom_settings[22]
port 15 nsew signal output
rlabel metal3 s 0 120232 800 120352 6 custom_settings[23]
port 16 nsew signal output
rlabel metal3 s 0 121320 800 121440 6 custom_settings[24]
port 17 nsew signal output
rlabel metal3 s 0 122408 800 122528 6 custom_settings[25]
port 18 nsew signal output
rlabel metal3 s 0 123496 800 123616 6 custom_settings[26]
port 19 nsew signal output
rlabel metal3 s 0 124584 800 124704 6 custom_settings[27]
port 20 nsew signal output
rlabel metal3 s 0 125672 800 125792 6 custom_settings[28]
port 21 nsew signal output
rlabel metal3 s 0 126760 800 126880 6 custom_settings[29]
port 22 nsew signal output
rlabel metal3 s 0 97384 800 97504 6 custom_settings[2]
port 23 nsew signal output
rlabel metal3 s 0 127848 800 127968 6 custom_settings[30]
port 24 nsew signal output
rlabel metal3 s 0 128936 800 129056 6 custom_settings[31]
port 25 nsew signal output
rlabel metal3 s 0 98472 800 98592 6 custom_settings[3]
port 26 nsew signal output
rlabel metal3 s 0 99560 800 99680 6 custom_settings[4]
port 27 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 custom_settings[5]
port 28 nsew signal output
rlabel metal3 s 0 101736 800 101856 6 custom_settings[6]
port 29 nsew signal output
rlabel metal3 s 0 102824 800 102944 6 custom_settings[7]
port 30 nsew signal output
rlabel metal3 s 0 103912 800 104032 6 custom_settings[8]
port 31 nsew signal output
rlabel metal3 s 0 105000 800 105120 6 custom_settings[9]
port 32 nsew signal output
rlabel metal2 s 2042 219200 2098 220000 6 io_in_0
port 33 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 io_oeb[0]
port 34 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 io_oeb[10]
port 35 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 io_oeb[11]
port 36 nsew signal output
rlabel metal3 s 0 25576 800 25696 6 io_oeb[12]
port 37 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 io_oeb[13]
port 38 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 io_oeb[14]
port 39 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 io_oeb[15]
port 40 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 io_oeb[16]
port 41 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 io_oeb[17]
port 42 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 io_oeb[18]
port 43 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 io_oeb[19]
port 44 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 io_oeb[1]
port 45 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 io_oeb[20]
port 46 nsew signal output
rlabel metal3 s 0 35368 800 35488 6 io_oeb[21]
port 47 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 io_oeb[22]
port 48 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 io_oeb[23]
port 49 nsew signal output
rlabel metal3 s 0 38632 800 38752 6 io_oeb[24]
port 50 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 io_oeb[25]
port 51 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 io_oeb[26]
port 52 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 io_oeb[27]
port 53 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 io_oeb[28]
port 54 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 io_oeb[29]
port 55 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 io_oeb[2]
port 56 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 io_oeb[30]
port 57 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 io_oeb[31]
port 58 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 io_oeb[32]
port 59 nsew signal output
rlabel metal3 s 0 48424 800 48544 6 io_oeb[33]
port 60 nsew signal output
rlabel metal3 s 0 49512 800 49632 6 io_oeb[34]
port 61 nsew signal output
rlabel metal3 s 0 50600 800 50720 6 io_oeb[35]
port 62 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 io_oeb[36]
port 63 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 io_oeb[37]
port 64 nsew signal output
rlabel metal3 s 0 15784 800 15904 6 io_oeb[3]
port 65 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 io_oeb[4]
port 66 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 io_oeb[5]
port 67 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 io_oeb[6]
port 68 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 io_oeb[7]
port 69 nsew signal output
rlabel metal3 s 0 21224 800 21344 6 io_oeb[8]
port 70 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 io_oeb[9]
port 71 nsew signal output
rlabel metal3 s 39200 70728 40000 70848 6 io_oeb_6502
port 72 nsew signal input
rlabel metal3 s 39200 189320 40000 189440 6 io_oeb_as1802
port 73 nsew signal input
rlabel metal3 s 0 169192 800 169312 6 io_oeb_scrapcpu[0]
port 74 nsew signal input
rlabel metal3 s 0 180072 800 180192 6 io_oeb_scrapcpu[10]
port 75 nsew signal input
rlabel metal3 s 0 181160 800 181280 6 io_oeb_scrapcpu[11]
port 76 nsew signal input
rlabel metal3 s 0 182248 800 182368 6 io_oeb_scrapcpu[12]
port 77 nsew signal input
rlabel metal3 s 0 183336 800 183456 6 io_oeb_scrapcpu[13]
port 78 nsew signal input
rlabel metal3 s 0 184424 800 184544 6 io_oeb_scrapcpu[14]
port 79 nsew signal input
rlabel metal3 s 0 185512 800 185632 6 io_oeb_scrapcpu[15]
port 80 nsew signal input
rlabel metal3 s 0 186600 800 186720 6 io_oeb_scrapcpu[16]
port 81 nsew signal input
rlabel metal3 s 0 187688 800 187808 6 io_oeb_scrapcpu[17]
port 82 nsew signal input
rlabel metal3 s 0 188776 800 188896 6 io_oeb_scrapcpu[18]
port 83 nsew signal input
rlabel metal3 s 0 189864 800 189984 6 io_oeb_scrapcpu[19]
port 84 nsew signal input
rlabel metal3 s 0 170280 800 170400 6 io_oeb_scrapcpu[1]
port 85 nsew signal input
rlabel metal3 s 0 190952 800 191072 6 io_oeb_scrapcpu[20]
port 86 nsew signal input
rlabel metal3 s 0 192040 800 192160 6 io_oeb_scrapcpu[21]
port 87 nsew signal input
rlabel metal3 s 0 193128 800 193248 6 io_oeb_scrapcpu[22]
port 88 nsew signal input
rlabel metal3 s 0 194216 800 194336 6 io_oeb_scrapcpu[23]
port 89 nsew signal input
rlabel metal3 s 0 195304 800 195424 6 io_oeb_scrapcpu[24]
port 90 nsew signal input
rlabel metal3 s 0 196392 800 196512 6 io_oeb_scrapcpu[25]
port 91 nsew signal input
rlabel metal3 s 0 197480 800 197600 6 io_oeb_scrapcpu[26]
port 92 nsew signal input
rlabel metal3 s 0 198568 800 198688 6 io_oeb_scrapcpu[27]
port 93 nsew signal input
rlabel metal3 s 0 199656 800 199776 6 io_oeb_scrapcpu[28]
port 94 nsew signal input
rlabel metal3 s 0 200744 800 200864 6 io_oeb_scrapcpu[29]
port 95 nsew signal input
rlabel metal3 s 0 171368 800 171488 6 io_oeb_scrapcpu[2]
port 96 nsew signal input
rlabel metal3 s 0 201832 800 201952 6 io_oeb_scrapcpu[30]
port 97 nsew signal input
rlabel metal3 s 0 202920 800 203040 6 io_oeb_scrapcpu[31]
port 98 nsew signal input
rlabel metal3 s 0 204008 800 204128 6 io_oeb_scrapcpu[32]
port 99 nsew signal input
rlabel metal3 s 0 205096 800 205216 6 io_oeb_scrapcpu[33]
port 100 nsew signal input
rlabel metal3 s 0 206184 800 206304 6 io_oeb_scrapcpu[34]
port 101 nsew signal input
rlabel metal3 s 0 207272 800 207392 6 io_oeb_scrapcpu[35]
port 102 nsew signal input
rlabel metal3 s 0 172456 800 172576 6 io_oeb_scrapcpu[3]
port 103 nsew signal input
rlabel metal3 s 0 173544 800 173664 6 io_oeb_scrapcpu[4]
port 104 nsew signal input
rlabel metal3 s 0 174632 800 174752 6 io_oeb_scrapcpu[5]
port 105 nsew signal input
rlabel metal3 s 0 175720 800 175840 6 io_oeb_scrapcpu[6]
port 106 nsew signal input
rlabel metal3 s 0 176808 800 176928 6 io_oeb_scrapcpu[7]
port 107 nsew signal input
rlabel metal3 s 0 177896 800 178016 6 io_oeb_scrapcpu[8]
port 108 nsew signal input
rlabel metal3 s 0 178984 800 179104 6 io_oeb_scrapcpu[9]
port 109 nsew signal input
rlabel metal3 s 0 130024 800 130144 6 io_oeb_vliw[0]
port 110 nsew signal input
rlabel metal3 s 0 140904 800 141024 6 io_oeb_vliw[10]
port 111 nsew signal input
rlabel metal3 s 0 141992 800 142112 6 io_oeb_vliw[11]
port 112 nsew signal input
rlabel metal3 s 0 143080 800 143200 6 io_oeb_vliw[12]
port 113 nsew signal input
rlabel metal3 s 0 144168 800 144288 6 io_oeb_vliw[13]
port 114 nsew signal input
rlabel metal3 s 0 145256 800 145376 6 io_oeb_vliw[14]
port 115 nsew signal input
rlabel metal3 s 0 146344 800 146464 6 io_oeb_vliw[15]
port 116 nsew signal input
rlabel metal3 s 0 147432 800 147552 6 io_oeb_vliw[16]
port 117 nsew signal input
rlabel metal3 s 0 148520 800 148640 6 io_oeb_vliw[17]
port 118 nsew signal input
rlabel metal3 s 0 149608 800 149728 6 io_oeb_vliw[18]
port 119 nsew signal input
rlabel metal3 s 0 150696 800 150816 6 io_oeb_vliw[19]
port 120 nsew signal input
rlabel metal3 s 0 131112 800 131232 6 io_oeb_vliw[1]
port 121 nsew signal input
rlabel metal3 s 0 151784 800 151904 6 io_oeb_vliw[20]
port 122 nsew signal input
rlabel metal3 s 0 152872 800 152992 6 io_oeb_vliw[21]
port 123 nsew signal input
rlabel metal3 s 0 153960 800 154080 6 io_oeb_vliw[22]
port 124 nsew signal input
rlabel metal3 s 0 155048 800 155168 6 io_oeb_vliw[23]
port 125 nsew signal input
rlabel metal3 s 0 156136 800 156256 6 io_oeb_vliw[24]
port 126 nsew signal input
rlabel metal3 s 0 157224 800 157344 6 io_oeb_vliw[25]
port 127 nsew signal input
rlabel metal3 s 0 158312 800 158432 6 io_oeb_vliw[26]
port 128 nsew signal input
rlabel metal3 s 0 159400 800 159520 6 io_oeb_vliw[27]
port 129 nsew signal input
rlabel metal3 s 0 160488 800 160608 6 io_oeb_vliw[28]
port 130 nsew signal input
rlabel metal3 s 0 161576 800 161696 6 io_oeb_vliw[29]
port 131 nsew signal input
rlabel metal3 s 0 132200 800 132320 6 io_oeb_vliw[2]
port 132 nsew signal input
rlabel metal3 s 0 162664 800 162784 6 io_oeb_vliw[30]
port 133 nsew signal input
rlabel metal3 s 0 163752 800 163872 6 io_oeb_vliw[31]
port 134 nsew signal input
rlabel metal3 s 0 164840 800 164960 6 io_oeb_vliw[32]
port 135 nsew signal input
rlabel metal3 s 0 165928 800 166048 6 io_oeb_vliw[33]
port 136 nsew signal input
rlabel metal3 s 0 167016 800 167136 6 io_oeb_vliw[34]
port 137 nsew signal input
rlabel metal3 s 0 168104 800 168224 6 io_oeb_vliw[35]
port 138 nsew signal input
rlabel metal3 s 0 133288 800 133408 6 io_oeb_vliw[3]
port 139 nsew signal input
rlabel metal3 s 0 134376 800 134496 6 io_oeb_vliw[4]
port 140 nsew signal input
rlabel metal3 s 0 135464 800 135584 6 io_oeb_vliw[5]
port 141 nsew signal input
rlabel metal3 s 0 136552 800 136672 6 io_oeb_vliw[6]
port 142 nsew signal input
rlabel metal3 s 0 137640 800 137760 6 io_oeb_vliw[7]
port 143 nsew signal input
rlabel metal3 s 0 138728 800 138848 6 io_oeb_vliw[8]
port 144 nsew signal input
rlabel metal3 s 0 139816 800 139936 6 io_oeb_vliw[9]
port 145 nsew signal input
rlabel metal3 s 39200 130568 40000 130688 6 io_oeb_z80[0]
port 146 nsew signal input
rlabel metal3 s 39200 136008 40000 136128 6 io_oeb_z80[10]
port 147 nsew signal input
rlabel metal3 s 39200 136552 40000 136672 6 io_oeb_z80[11]
port 148 nsew signal input
rlabel metal3 s 39200 137096 40000 137216 6 io_oeb_z80[12]
port 149 nsew signal input
rlabel metal3 s 39200 137640 40000 137760 6 io_oeb_z80[13]
port 150 nsew signal input
rlabel metal3 s 39200 138184 40000 138304 6 io_oeb_z80[14]
port 151 nsew signal input
rlabel metal3 s 39200 138728 40000 138848 6 io_oeb_z80[15]
port 152 nsew signal input
rlabel metal3 s 39200 139272 40000 139392 6 io_oeb_z80[16]
port 153 nsew signal input
rlabel metal3 s 39200 139816 40000 139936 6 io_oeb_z80[17]
port 154 nsew signal input
rlabel metal3 s 39200 140360 40000 140480 6 io_oeb_z80[18]
port 155 nsew signal input
rlabel metal3 s 39200 140904 40000 141024 6 io_oeb_z80[19]
port 156 nsew signal input
rlabel metal3 s 39200 131112 40000 131232 6 io_oeb_z80[1]
port 157 nsew signal input
rlabel metal3 s 39200 141448 40000 141568 6 io_oeb_z80[20]
port 158 nsew signal input
rlabel metal3 s 39200 141992 40000 142112 6 io_oeb_z80[21]
port 159 nsew signal input
rlabel metal3 s 39200 142536 40000 142656 6 io_oeb_z80[22]
port 160 nsew signal input
rlabel metal3 s 39200 143080 40000 143200 6 io_oeb_z80[23]
port 161 nsew signal input
rlabel metal3 s 39200 143624 40000 143744 6 io_oeb_z80[24]
port 162 nsew signal input
rlabel metal3 s 39200 144168 40000 144288 6 io_oeb_z80[25]
port 163 nsew signal input
rlabel metal3 s 39200 144712 40000 144832 6 io_oeb_z80[26]
port 164 nsew signal input
rlabel metal3 s 39200 145256 40000 145376 6 io_oeb_z80[27]
port 165 nsew signal input
rlabel metal3 s 39200 145800 40000 145920 6 io_oeb_z80[28]
port 166 nsew signal input
rlabel metal3 s 39200 146344 40000 146464 6 io_oeb_z80[29]
port 167 nsew signal input
rlabel metal3 s 39200 131656 40000 131776 6 io_oeb_z80[2]
port 168 nsew signal input
rlabel metal3 s 39200 146888 40000 147008 6 io_oeb_z80[30]
port 169 nsew signal input
rlabel metal3 s 39200 147432 40000 147552 6 io_oeb_z80[31]
port 170 nsew signal input
rlabel metal3 s 39200 147976 40000 148096 6 io_oeb_z80[32]
port 171 nsew signal input
rlabel metal3 s 39200 148520 40000 148640 6 io_oeb_z80[33]
port 172 nsew signal input
rlabel metal3 s 39200 149064 40000 149184 6 io_oeb_z80[34]
port 173 nsew signal input
rlabel metal3 s 39200 149608 40000 149728 6 io_oeb_z80[35]
port 174 nsew signal input
rlabel metal3 s 39200 132200 40000 132320 6 io_oeb_z80[3]
port 175 nsew signal input
rlabel metal3 s 39200 132744 40000 132864 6 io_oeb_z80[4]
port 176 nsew signal input
rlabel metal3 s 39200 133288 40000 133408 6 io_oeb_z80[5]
port 177 nsew signal input
rlabel metal3 s 39200 133832 40000 133952 6 io_oeb_z80[6]
port 178 nsew signal input
rlabel metal3 s 39200 134376 40000 134496 6 io_oeb_z80[7]
port 179 nsew signal input
rlabel metal3 s 39200 134920 40000 135040 6 io_oeb_z80[8]
port 180 nsew signal input
rlabel metal3 s 39200 135464 40000 135584 6 io_oeb_z80[9]
port 181 nsew signal input
rlabel metal3 s 39200 30472 40000 30592 6 io_out[0]
port 182 nsew signal output
rlabel metal3 s 39200 35912 40000 36032 6 io_out[10]
port 183 nsew signal output
rlabel metal3 s 39200 36456 40000 36576 6 io_out[11]
port 184 nsew signal output
rlabel metal3 s 39200 37000 40000 37120 6 io_out[12]
port 185 nsew signal output
rlabel metal3 s 39200 37544 40000 37664 6 io_out[13]
port 186 nsew signal output
rlabel metal3 s 39200 38088 40000 38208 6 io_out[14]
port 187 nsew signal output
rlabel metal3 s 39200 38632 40000 38752 6 io_out[15]
port 188 nsew signal output
rlabel metal3 s 39200 39176 40000 39296 6 io_out[16]
port 189 nsew signal output
rlabel metal3 s 39200 39720 40000 39840 6 io_out[17]
port 190 nsew signal output
rlabel metal3 s 39200 40264 40000 40384 6 io_out[18]
port 191 nsew signal output
rlabel metal3 s 39200 40808 40000 40928 6 io_out[19]
port 192 nsew signal output
rlabel metal3 s 39200 31016 40000 31136 6 io_out[1]
port 193 nsew signal output
rlabel metal3 s 39200 41352 40000 41472 6 io_out[20]
port 194 nsew signal output
rlabel metal3 s 39200 41896 40000 42016 6 io_out[21]
port 195 nsew signal output
rlabel metal3 s 39200 42440 40000 42560 6 io_out[22]
port 196 nsew signal output
rlabel metal3 s 39200 42984 40000 43104 6 io_out[23]
port 197 nsew signal output
rlabel metal3 s 39200 43528 40000 43648 6 io_out[24]
port 198 nsew signal output
rlabel metal3 s 39200 44072 40000 44192 6 io_out[25]
port 199 nsew signal output
rlabel metal3 s 39200 44616 40000 44736 6 io_out[26]
port 200 nsew signal output
rlabel metal3 s 39200 45160 40000 45280 6 io_out[27]
port 201 nsew signal output
rlabel metal3 s 39200 45704 40000 45824 6 io_out[28]
port 202 nsew signal output
rlabel metal3 s 39200 46248 40000 46368 6 io_out[29]
port 203 nsew signal output
rlabel metal3 s 39200 31560 40000 31680 6 io_out[2]
port 204 nsew signal output
rlabel metal3 s 39200 46792 40000 46912 6 io_out[30]
port 205 nsew signal output
rlabel metal3 s 39200 47336 40000 47456 6 io_out[31]
port 206 nsew signal output
rlabel metal3 s 39200 47880 40000 48000 6 io_out[32]
port 207 nsew signal output
rlabel metal3 s 39200 48424 40000 48544 6 io_out[33]
port 208 nsew signal output
rlabel metal3 s 39200 48968 40000 49088 6 io_out[34]
port 209 nsew signal output
rlabel metal3 s 39200 49512 40000 49632 6 io_out[35]
port 210 nsew signal output
rlabel metal3 s 39200 50056 40000 50176 6 io_out[36]
port 211 nsew signal output
rlabel metal3 s 39200 50600 40000 50720 6 io_out[37]
port 212 nsew signal output
rlabel metal3 s 39200 32104 40000 32224 6 io_out[3]
port 213 nsew signal output
rlabel metal3 s 39200 32648 40000 32768 6 io_out[4]
port 214 nsew signal output
rlabel metal3 s 39200 33192 40000 33312 6 io_out[5]
port 215 nsew signal output
rlabel metal3 s 39200 33736 40000 33856 6 io_out[6]
port 216 nsew signal output
rlabel metal3 s 39200 34280 40000 34400 6 io_out[7]
port 217 nsew signal output
rlabel metal3 s 39200 34824 40000 34944 6 io_out[8]
port 218 nsew signal output
rlabel metal3 s 39200 35368 40000 35488 6 io_out[9]
port 219 nsew signal output
rlabel metal3 s 39200 51144 40000 51264 6 io_out_6502[0]
port 220 nsew signal input
rlabel metal3 s 39200 56584 40000 56704 6 io_out_6502[10]
port 221 nsew signal input
rlabel metal3 s 39200 57128 40000 57248 6 io_out_6502[11]
port 222 nsew signal input
rlabel metal3 s 39200 57672 40000 57792 6 io_out_6502[12]
port 223 nsew signal input
rlabel metal3 s 39200 58216 40000 58336 6 io_out_6502[13]
port 224 nsew signal input
rlabel metal3 s 39200 58760 40000 58880 6 io_out_6502[14]
port 225 nsew signal input
rlabel metal3 s 39200 59304 40000 59424 6 io_out_6502[15]
port 226 nsew signal input
rlabel metal3 s 39200 59848 40000 59968 6 io_out_6502[16]
port 227 nsew signal input
rlabel metal3 s 39200 60392 40000 60512 6 io_out_6502[17]
port 228 nsew signal input
rlabel metal3 s 39200 60936 40000 61056 6 io_out_6502[18]
port 229 nsew signal input
rlabel metal3 s 39200 61480 40000 61600 6 io_out_6502[19]
port 230 nsew signal input
rlabel metal3 s 39200 51688 40000 51808 6 io_out_6502[1]
port 231 nsew signal input
rlabel metal3 s 39200 62024 40000 62144 6 io_out_6502[20]
port 232 nsew signal input
rlabel metal3 s 39200 62568 40000 62688 6 io_out_6502[21]
port 233 nsew signal input
rlabel metal3 s 39200 63112 40000 63232 6 io_out_6502[22]
port 234 nsew signal input
rlabel metal3 s 39200 63656 40000 63776 6 io_out_6502[23]
port 235 nsew signal input
rlabel metal3 s 39200 64200 40000 64320 6 io_out_6502[24]
port 236 nsew signal input
rlabel metal3 s 39200 64744 40000 64864 6 io_out_6502[25]
port 237 nsew signal input
rlabel metal3 s 39200 65288 40000 65408 6 io_out_6502[26]
port 238 nsew signal input
rlabel metal3 s 39200 65832 40000 65952 6 io_out_6502[27]
port 239 nsew signal input
rlabel metal3 s 39200 66376 40000 66496 6 io_out_6502[28]
port 240 nsew signal input
rlabel metal3 s 39200 66920 40000 67040 6 io_out_6502[29]
port 241 nsew signal input
rlabel metal3 s 39200 52232 40000 52352 6 io_out_6502[2]
port 242 nsew signal input
rlabel metal3 s 39200 67464 40000 67584 6 io_out_6502[30]
port 243 nsew signal input
rlabel metal3 s 39200 68008 40000 68128 6 io_out_6502[31]
port 244 nsew signal input
rlabel metal3 s 39200 68552 40000 68672 6 io_out_6502[32]
port 245 nsew signal input
rlabel metal3 s 39200 69096 40000 69216 6 io_out_6502[33]
port 246 nsew signal input
rlabel metal3 s 39200 69640 40000 69760 6 io_out_6502[34]
port 247 nsew signal input
rlabel metal3 s 39200 70184 40000 70304 6 io_out_6502[35]
port 248 nsew signal input
rlabel metal3 s 39200 52776 40000 52896 6 io_out_6502[3]
port 249 nsew signal input
rlabel metal3 s 39200 53320 40000 53440 6 io_out_6502[4]
port 250 nsew signal input
rlabel metal3 s 39200 53864 40000 53984 6 io_out_6502[5]
port 251 nsew signal input
rlabel metal3 s 39200 54408 40000 54528 6 io_out_6502[6]
port 252 nsew signal input
rlabel metal3 s 39200 54952 40000 55072 6 io_out_6502[7]
port 253 nsew signal input
rlabel metal3 s 39200 55496 40000 55616 6 io_out_6502[8]
port 254 nsew signal input
rlabel metal3 s 39200 56040 40000 56160 6 io_out_6502[9]
port 255 nsew signal input
rlabel metal3 s 39200 169736 40000 169856 6 io_out_as1802[0]
port 256 nsew signal input
rlabel metal3 s 39200 175176 40000 175296 6 io_out_as1802[10]
port 257 nsew signal input
rlabel metal3 s 39200 175720 40000 175840 6 io_out_as1802[11]
port 258 nsew signal input
rlabel metal3 s 39200 176264 40000 176384 6 io_out_as1802[12]
port 259 nsew signal input
rlabel metal3 s 39200 176808 40000 176928 6 io_out_as1802[13]
port 260 nsew signal input
rlabel metal3 s 39200 177352 40000 177472 6 io_out_as1802[14]
port 261 nsew signal input
rlabel metal3 s 39200 177896 40000 178016 6 io_out_as1802[15]
port 262 nsew signal input
rlabel metal3 s 39200 178440 40000 178560 6 io_out_as1802[16]
port 263 nsew signal input
rlabel metal3 s 39200 178984 40000 179104 6 io_out_as1802[17]
port 264 nsew signal input
rlabel metal3 s 39200 179528 40000 179648 6 io_out_as1802[18]
port 265 nsew signal input
rlabel metal3 s 39200 180072 40000 180192 6 io_out_as1802[19]
port 266 nsew signal input
rlabel metal3 s 39200 170280 40000 170400 6 io_out_as1802[1]
port 267 nsew signal input
rlabel metal3 s 39200 180616 40000 180736 6 io_out_as1802[20]
port 268 nsew signal input
rlabel metal3 s 39200 181160 40000 181280 6 io_out_as1802[21]
port 269 nsew signal input
rlabel metal3 s 39200 181704 40000 181824 6 io_out_as1802[22]
port 270 nsew signal input
rlabel metal3 s 39200 182248 40000 182368 6 io_out_as1802[23]
port 271 nsew signal input
rlabel metal3 s 39200 182792 40000 182912 6 io_out_as1802[24]
port 272 nsew signal input
rlabel metal3 s 39200 183336 40000 183456 6 io_out_as1802[25]
port 273 nsew signal input
rlabel metal3 s 39200 183880 40000 184000 6 io_out_as1802[26]
port 274 nsew signal input
rlabel metal3 s 39200 184424 40000 184544 6 io_out_as1802[27]
port 275 nsew signal input
rlabel metal3 s 39200 184968 40000 185088 6 io_out_as1802[28]
port 276 nsew signal input
rlabel metal3 s 39200 185512 40000 185632 6 io_out_as1802[29]
port 277 nsew signal input
rlabel metal3 s 39200 170824 40000 170944 6 io_out_as1802[2]
port 278 nsew signal input
rlabel metal3 s 39200 186056 40000 186176 6 io_out_as1802[30]
port 279 nsew signal input
rlabel metal3 s 39200 186600 40000 186720 6 io_out_as1802[31]
port 280 nsew signal input
rlabel metal3 s 39200 187144 40000 187264 6 io_out_as1802[32]
port 281 nsew signal input
rlabel metal3 s 39200 187688 40000 187808 6 io_out_as1802[33]
port 282 nsew signal input
rlabel metal3 s 39200 188232 40000 188352 6 io_out_as1802[34]
port 283 nsew signal input
rlabel metal3 s 39200 188776 40000 188896 6 io_out_as1802[35]
port 284 nsew signal input
rlabel metal3 s 39200 171368 40000 171488 6 io_out_as1802[3]
port 285 nsew signal input
rlabel metal3 s 39200 171912 40000 172032 6 io_out_as1802[4]
port 286 nsew signal input
rlabel metal3 s 39200 172456 40000 172576 6 io_out_as1802[5]
port 287 nsew signal input
rlabel metal3 s 39200 173000 40000 173120 6 io_out_as1802[6]
port 288 nsew signal input
rlabel metal3 s 39200 173544 40000 173664 6 io_out_as1802[7]
port 289 nsew signal input
rlabel metal3 s 39200 174088 40000 174208 6 io_out_as1802[8]
port 290 nsew signal input
rlabel metal3 s 39200 174632 40000 174752 6 io_out_as1802[9]
port 291 nsew signal input
rlabel metal3 s 39200 150152 40000 150272 6 io_out_scrapcpu[0]
port 292 nsew signal input
rlabel metal3 s 39200 155592 40000 155712 6 io_out_scrapcpu[10]
port 293 nsew signal input
rlabel metal3 s 39200 156136 40000 156256 6 io_out_scrapcpu[11]
port 294 nsew signal input
rlabel metal3 s 39200 156680 40000 156800 6 io_out_scrapcpu[12]
port 295 nsew signal input
rlabel metal3 s 39200 157224 40000 157344 6 io_out_scrapcpu[13]
port 296 nsew signal input
rlabel metal3 s 39200 157768 40000 157888 6 io_out_scrapcpu[14]
port 297 nsew signal input
rlabel metal3 s 39200 158312 40000 158432 6 io_out_scrapcpu[15]
port 298 nsew signal input
rlabel metal3 s 39200 158856 40000 158976 6 io_out_scrapcpu[16]
port 299 nsew signal input
rlabel metal3 s 39200 159400 40000 159520 6 io_out_scrapcpu[17]
port 300 nsew signal input
rlabel metal3 s 39200 159944 40000 160064 6 io_out_scrapcpu[18]
port 301 nsew signal input
rlabel metal3 s 39200 160488 40000 160608 6 io_out_scrapcpu[19]
port 302 nsew signal input
rlabel metal3 s 39200 150696 40000 150816 6 io_out_scrapcpu[1]
port 303 nsew signal input
rlabel metal3 s 39200 161032 40000 161152 6 io_out_scrapcpu[20]
port 304 nsew signal input
rlabel metal3 s 39200 161576 40000 161696 6 io_out_scrapcpu[21]
port 305 nsew signal input
rlabel metal3 s 39200 162120 40000 162240 6 io_out_scrapcpu[22]
port 306 nsew signal input
rlabel metal3 s 39200 162664 40000 162784 6 io_out_scrapcpu[23]
port 307 nsew signal input
rlabel metal3 s 39200 163208 40000 163328 6 io_out_scrapcpu[24]
port 308 nsew signal input
rlabel metal3 s 39200 163752 40000 163872 6 io_out_scrapcpu[25]
port 309 nsew signal input
rlabel metal3 s 39200 164296 40000 164416 6 io_out_scrapcpu[26]
port 310 nsew signal input
rlabel metal3 s 39200 164840 40000 164960 6 io_out_scrapcpu[27]
port 311 nsew signal input
rlabel metal3 s 39200 165384 40000 165504 6 io_out_scrapcpu[28]
port 312 nsew signal input
rlabel metal3 s 39200 165928 40000 166048 6 io_out_scrapcpu[29]
port 313 nsew signal input
rlabel metal3 s 39200 151240 40000 151360 6 io_out_scrapcpu[2]
port 314 nsew signal input
rlabel metal3 s 39200 166472 40000 166592 6 io_out_scrapcpu[30]
port 315 nsew signal input
rlabel metal3 s 39200 167016 40000 167136 6 io_out_scrapcpu[31]
port 316 nsew signal input
rlabel metal3 s 39200 167560 40000 167680 6 io_out_scrapcpu[32]
port 317 nsew signal input
rlabel metal3 s 39200 168104 40000 168224 6 io_out_scrapcpu[33]
port 318 nsew signal input
rlabel metal3 s 39200 168648 40000 168768 6 io_out_scrapcpu[34]
port 319 nsew signal input
rlabel metal3 s 39200 169192 40000 169312 6 io_out_scrapcpu[35]
port 320 nsew signal input
rlabel metal3 s 39200 151784 40000 151904 6 io_out_scrapcpu[3]
port 321 nsew signal input
rlabel metal3 s 39200 152328 40000 152448 6 io_out_scrapcpu[4]
port 322 nsew signal input
rlabel metal3 s 39200 152872 40000 152992 6 io_out_scrapcpu[5]
port 323 nsew signal input
rlabel metal3 s 39200 153416 40000 153536 6 io_out_scrapcpu[6]
port 324 nsew signal input
rlabel metal3 s 39200 153960 40000 154080 6 io_out_scrapcpu[7]
port 325 nsew signal input
rlabel metal3 s 39200 154504 40000 154624 6 io_out_scrapcpu[8]
port 326 nsew signal input
rlabel metal3 s 39200 155048 40000 155168 6 io_out_scrapcpu[9]
port 327 nsew signal input
rlabel metal2 s 3882 219200 3938 220000 6 io_out_vliw[0]
port 328 nsew signal input
rlabel metal2 s 13082 219200 13138 220000 6 io_out_vliw[10]
port 329 nsew signal input
rlabel metal2 s 14002 219200 14058 220000 6 io_out_vliw[11]
port 330 nsew signal input
rlabel metal2 s 14922 219200 14978 220000 6 io_out_vliw[12]
port 331 nsew signal input
rlabel metal2 s 15842 219200 15898 220000 6 io_out_vliw[13]
port 332 nsew signal input
rlabel metal2 s 16762 219200 16818 220000 6 io_out_vliw[14]
port 333 nsew signal input
rlabel metal2 s 17682 219200 17738 220000 6 io_out_vliw[15]
port 334 nsew signal input
rlabel metal2 s 18602 219200 18658 220000 6 io_out_vliw[16]
port 335 nsew signal input
rlabel metal2 s 19522 219200 19578 220000 6 io_out_vliw[17]
port 336 nsew signal input
rlabel metal2 s 20442 219200 20498 220000 6 io_out_vliw[18]
port 337 nsew signal input
rlabel metal2 s 21362 219200 21418 220000 6 io_out_vliw[19]
port 338 nsew signal input
rlabel metal2 s 4802 219200 4858 220000 6 io_out_vliw[1]
port 339 nsew signal input
rlabel metal2 s 22282 219200 22338 220000 6 io_out_vliw[20]
port 340 nsew signal input
rlabel metal2 s 23202 219200 23258 220000 6 io_out_vliw[21]
port 341 nsew signal input
rlabel metal2 s 24122 219200 24178 220000 6 io_out_vliw[22]
port 342 nsew signal input
rlabel metal2 s 25042 219200 25098 220000 6 io_out_vliw[23]
port 343 nsew signal input
rlabel metal2 s 25962 219200 26018 220000 6 io_out_vliw[24]
port 344 nsew signal input
rlabel metal2 s 26882 219200 26938 220000 6 io_out_vliw[25]
port 345 nsew signal input
rlabel metal2 s 27802 219200 27858 220000 6 io_out_vliw[26]
port 346 nsew signal input
rlabel metal2 s 28722 219200 28778 220000 6 io_out_vliw[27]
port 347 nsew signal input
rlabel metal2 s 29642 219200 29698 220000 6 io_out_vliw[28]
port 348 nsew signal input
rlabel metal2 s 30562 219200 30618 220000 6 io_out_vliw[29]
port 349 nsew signal input
rlabel metal2 s 5722 219200 5778 220000 6 io_out_vliw[2]
port 350 nsew signal input
rlabel metal2 s 31482 219200 31538 220000 6 io_out_vliw[30]
port 351 nsew signal input
rlabel metal2 s 32402 219200 32458 220000 6 io_out_vliw[31]
port 352 nsew signal input
rlabel metal2 s 33322 219200 33378 220000 6 io_out_vliw[32]
port 353 nsew signal input
rlabel metal2 s 34242 219200 34298 220000 6 io_out_vliw[33]
port 354 nsew signal input
rlabel metal2 s 35162 219200 35218 220000 6 io_out_vliw[34]
port 355 nsew signal input
rlabel metal2 s 36082 219200 36138 220000 6 io_out_vliw[35]
port 356 nsew signal input
rlabel metal2 s 6642 219200 6698 220000 6 io_out_vliw[3]
port 357 nsew signal input
rlabel metal2 s 7562 219200 7618 220000 6 io_out_vliw[4]
port 358 nsew signal input
rlabel metal2 s 8482 219200 8538 220000 6 io_out_vliw[5]
port 359 nsew signal input
rlabel metal2 s 9402 219200 9458 220000 6 io_out_vliw[6]
port 360 nsew signal input
rlabel metal2 s 10322 219200 10378 220000 6 io_out_vliw[7]
port 361 nsew signal input
rlabel metal2 s 11242 219200 11298 220000 6 io_out_vliw[8]
port 362 nsew signal input
rlabel metal2 s 12162 219200 12218 220000 6 io_out_vliw[9]
port 363 nsew signal input
rlabel metal3 s 39200 110440 40000 110560 6 io_out_z80[0]
port 364 nsew signal input
rlabel metal3 s 39200 115880 40000 116000 6 io_out_z80[10]
port 365 nsew signal input
rlabel metal3 s 39200 116424 40000 116544 6 io_out_z80[11]
port 366 nsew signal input
rlabel metal3 s 39200 116968 40000 117088 6 io_out_z80[12]
port 367 nsew signal input
rlabel metal3 s 39200 117512 40000 117632 6 io_out_z80[13]
port 368 nsew signal input
rlabel metal3 s 39200 118056 40000 118176 6 io_out_z80[14]
port 369 nsew signal input
rlabel metal3 s 39200 118600 40000 118720 6 io_out_z80[15]
port 370 nsew signal input
rlabel metal3 s 39200 119144 40000 119264 6 io_out_z80[16]
port 371 nsew signal input
rlabel metal3 s 39200 119688 40000 119808 6 io_out_z80[17]
port 372 nsew signal input
rlabel metal3 s 39200 120232 40000 120352 6 io_out_z80[18]
port 373 nsew signal input
rlabel metal3 s 39200 120776 40000 120896 6 io_out_z80[19]
port 374 nsew signal input
rlabel metal3 s 39200 110984 40000 111104 6 io_out_z80[1]
port 375 nsew signal input
rlabel metal3 s 39200 121320 40000 121440 6 io_out_z80[20]
port 376 nsew signal input
rlabel metal3 s 39200 121864 40000 121984 6 io_out_z80[21]
port 377 nsew signal input
rlabel metal3 s 39200 122408 40000 122528 6 io_out_z80[22]
port 378 nsew signal input
rlabel metal3 s 39200 122952 40000 123072 6 io_out_z80[23]
port 379 nsew signal input
rlabel metal3 s 39200 123496 40000 123616 6 io_out_z80[24]
port 380 nsew signal input
rlabel metal3 s 39200 124040 40000 124160 6 io_out_z80[25]
port 381 nsew signal input
rlabel metal3 s 39200 124584 40000 124704 6 io_out_z80[26]
port 382 nsew signal input
rlabel metal3 s 39200 125128 40000 125248 6 io_out_z80[27]
port 383 nsew signal input
rlabel metal3 s 39200 125672 40000 125792 6 io_out_z80[28]
port 384 nsew signal input
rlabel metal3 s 39200 126216 40000 126336 6 io_out_z80[29]
port 385 nsew signal input
rlabel metal3 s 39200 111528 40000 111648 6 io_out_z80[2]
port 386 nsew signal input
rlabel metal3 s 39200 126760 40000 126880 6 io_out_z80[30]
port 387 nsew signal input
rlabel metal3 s 39200 127304 40000 127424 6 io_out_z80[31]
port 388 nsew signal input
rlabel metal3 s 39200 127848 40000 127968 6 io_out_z80[32]
port 389 nsew signal input
rlabel metal3 s 39200 128392 40000 128512 6 io_out_z80[33]
port 390 nsew signal input
rlabel metal3 s 39200 128936 40000 129056 6 io_out_z80[34]
port 391 nsew signal input
rlabel metal3 s 39200 129480 40000 129600 6 io_out_z80[35]
port 392 nsew signal input
rlabel metal3 s 39200 112072 40000 112192 6 io_out_z80[3]
port 393 nsew signal input
rlabel metal3 s 39200 112616 40000 112736 6 io_out_z80[4]
port 394 nsew signal input
rlabel metal3 s 39200 113160 40000 113280 6 io_out_z80[5]
port 395 nsew signal input
rlabel metal3 s 39200 113704 40000 113824 6 io_out_z80[6]
port 396 nsew signal input
rlabel metal3 s 39200 114248 40000 114368 6 io_out_z80[7]
port 397 nsew signal input
rlabel metal3 s 39200 114792 40000 114912 6 io_out_z80[8]
port 398 nsew signal input
rlabel metal3 s 39200 115336 40000 115456 6 io_out_z80[9]
port 399 nsew signal input
rlabel metal3 s 39200 88680 40000 88800 6 la_data_out[0]
port 400 nsew signal output
rlabel metal3 s 39200 94120 40000 94240 6 la_data_out[10]
port 401 nsew signal output
rlabel metal3 s 39200 94664 40000 94784 6 la_data_out[11]
port 402 nsew signal output
rlabel metal3 s 39200 95208 40000 95328 6 la_data_out[12]
port 403 nsew signal output
rlabel metal3 s 39200 95752 40000 95872 6 la_data_out[13]
port 404 nsew signal output
rlabel metal3 s 39200 96296 40000 96416 6 la_data_out[14]
port 405 nsew signal output
rlabel metal3 s 39200 96840 40000 96960 6 la_data_out[15]
port 406 nsew signal output
rlabel metal3 s 39200 97384 40000 97504 6 la_data_out[16]
port 407 nsew signal output
rlabel metal3 s 39200 97928 40000 98048 6 la_data_out[17]
port 408 nsew signal output
rlabel metal3 s 39200 98472 40000 98592 6 la_data_out[18]
port 409 nsew signal output
rlabel metal3 s 39200 99016 40000 99136 6 la_data_out[19]
port 410 nsew signal output
rlabel metal3 s 39200 89224 40000 89344 6 la_data_out[1]
port 411 nsew signal output
rlabel metal3 s 39200 99560 40000 99680 6 la_data_out[20]
port 412 nsew signal output
rlabel metal3 s 39200 100104 40000 100224 6 la_data_out[21]
port 413 nsew signal output
rlabel metal3 s 39200 100648 40000 100768 6 la_data_out[22]
port 414 nsew signal output
rlabel metal3 s 39200 101192 40000 101312 6 la_data_out[23]
port 415 nsew signal output
rlabel metal3 s 39200 101736 40000 101856 6 la_data_out[24]
port 416 nsew signal output
rlabel metal3 s 39200 102280 40000 102400 6 la_data_out[25]
port 417 nsew signal output
rlabel metal3 s 39200 102824 40000 102944 6 la_data_out[26]
port 418 nsew signal output
rlabel metal3 s 39200 103368 40000 103488 6 la_data_out[27]
port 419 nsew signal output
rlabel metal3 s 39200 103912 40000 104032 6 la_data_out[28]
port 420 nsew signal output
rlabel metal3 s 39200 104456 40000 104576 6 la_data_out[29]
port 421 nsew signal output
rlabel metal3 s 39200 89768 40000 89888 6 la_data_out[2]
port 422 nsew signal output
rlabel metal3 s 39200 105000 40000 105120 6 la_data_out[30]
port 423 nsew signal output
rlabel metal3 s 39200 105544 40000 105664 6 la_data_out[31]
port 424 nsew signal output
rlabel metal3 s 39200 106088 40000 106208 6 la_data_out[32]
port 425 nsew signal output
rlabel metal3 s 39200 106632 40000 106752 6 la_data_out[33]
port 426 nsew signal output
rlabel metal3 s 39200 107176 40000 107296 6 la_data_out[34]
port 427 nsew signal output
rlabel metal3 s 39200 107720 40000 107840 6 la_data_out[35]
port 428 nsew signal output
rlabel metal3 s 39200 108264 40000 108384 6 la_data_out[36]
port 429 nsew signal output
rlabel metal3 s 39200 108808 40000 108928 6 la_data_out[37]
port 430 nsew signal output
rlabel metal3 s 39200 109352 40000 109472 6 la_data_out[38]
port 431 nsew signal output
rlabel metal3 s 39200 109896 40000 110016 6 la_data_out[39]
port 432 nsew signal output
rlabel metal3 s 39200 90312 40000 90432 6 la_data_out[3]
port 433 nsew signal output
rlabel metal3 s 39200 90856 40000 90976 6 la_data_out[4]
port 434 nsew signal output
rlabel metal3 s 39200 91400 40000 91520 6 la_data_out[5]
port 435 nsew signal output
rlabel metal3 s 39200 91944 40000 92064 6 la_data_out[6]
port 436 nsew signal output
rlabel metal3 s 39200 92488 40000 92608 6 la_data_out[7]
port 437 nsew signal output
rlabel metal3 s 39200 93032 40000 93152 6 la_data_out[8]
port 438 nsew signal output
rlabel metal3 s 39200 93576 40000 93696 6 la_data_out[9]
port 439 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 rst_6502
port 440 nsew signal output
rlabel metal2 s 37922 219200 37978 220000 6 rst_as1802
port 441 nsew signal output
rlabel metal2 s 37002 219200 37058 220000 6 rst_scrapcpu
port 442 nsew signal output
rlabel metal2 s 2962 219200 3018 220000 6 rst_vliw
port 443 nsew signal output
rlabel metal3 s 39200 130024 40000 130144 6 rst_z80
port 444 nsew signal output
rlabel metal4 s 4208 2128 4528 217648 6 vccd1
port 445 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 217648 6 vccd1
port 445 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 217648 6 vssd1
port 446 nsew ground bidirectional
rlabel metal3 s 0 53864 800 53984 6 wb_clk_i
port 447 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 wb_rst_i
port 448 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 wbs_ack_o
port 449 nsew signal output
rlabel metal2 s 846 0 902 800 6 wbs_adr_i[0]
port 450 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wbs_adr_i[10]
port 451 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 wbs_adr_i[11]
port 452 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[12]
port 453 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[13]
port 454 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[14]
port 455 nsew signal input
rlabel metal2 s 18786 0 18842 800 6 wbs_adr_i[15]
port 456 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_adr_i[16]
port 457 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[17]
port 458 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_adr_i[18]
port 459 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[19]
port 460 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 wbs_adr_i[1]
port 461 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_adr_i[20]
port 462 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_adr_i[21]
port 463 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_adr_i[22]
port 464 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_adr_i[23]
port 465 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[24]
port 466 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_adr_i[25]
port 467 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_adr_i[26]
port 468 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_adr_i[27]
port 469 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_adr_i[28]
port 470 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_adr_i[29]
port 471 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_adr_i[2]
port 472 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 wbs_adr_i[30]
port 473 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_adr_i[31]
port 474 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_adr_i[3]
port 475 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_adr_i[4]
port 476 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[5]
port 477 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[6]
port 478 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[7]
port 479 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_adr_i[8]
port 480 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 wbs_adr_i[9]
port 481 nsew signal input
rlabel metal3 s 0 91944 800 92064 6 wbs_cyc_i
port 482 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 wbs_dat_i[0]
port 483 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 wbs_dat_i[10]
port 484 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 wbs_dat_i[11]
port 485 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 wbs_dat_i[12]
port 486 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 wbs_dat_i[13]
port 487 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 wbs_dat_i[14]
port 488 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 wbs_dat_i[15]
port 489 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 wbs_dat_i[16]
port 490 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 wbs_dat_i[17]
port 491 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 wbs_dat_i[18]
port 492 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 wbs_dat_i[19]
port 493 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 wbs_dat_i[1]
port 494 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 wbs_dat_i[20]
port 495 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 wbs_dat_i[21]
port 496 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 wbs_dat_i[22]
port 497 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 wbs_dat_i[23]
port 498 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 wbs_dat_i[24]
port 499 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 wbs_dat_i[25]
port 500 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 wbs_dat_i[26]
port 501 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 wbs_dat_i[27]
port 502 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 wbs_dat_i[28]
port 503 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 wbs_dat_i[29]
port 504 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 wbs_dat_i[2]
port 505 nsew signal input
rlabel metal3 s 0 88680 800 88800 6 wbs_dat_i[30]
port 506 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 wbs_dat_i[31]
port 507 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 wbs_dat_i[3]
port 508 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 wbs_dat_i[4]
port 509 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 wbs_dat_i[5]
port 510 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 wbs_dat_i[6]
port 511 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 wbs_dat_i[7]
port 512 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 wbs_dat_i[8]
port 513 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 wbs_dat_i[9]
port 514 nsew signal input
rlabel metal3 s 39200 71272 40000 71392 6 wbs_dat_o[0]
port 515 nsew signal output
rlabel metal3 s 39200 76712 40000 76832 6 wbs_dat_o[10]
port 516 nsew signal output
rlabel metal3 s 39200 77256 40000 77376 6 wbs_dat_o[11]
port 517 nsew signal output
rlabel metal3 s 39200 77800 40000 77920 6 wbs_dat_o[12]
port 518 nsew signal output
rlabel metal3 s 39200 78344 40000 78464 6 wbs_dat_o[13]
port 519 nsew signal output
rlabel metal3 s 39200 78888 40000 79008 6 wbs_dat_o[14]
port 520 nsew signal output
rlabel metal3 s 39200 79432 40000 79552 6 wbs_dat_o[15]
port 521 nsew signal output
rlabel metal3 s 39200 79976 40000 80096 6 wbs_dat_o[16]
port 522 nsew signal output
rlabel metal3 s 39200 80520 40000 80640 6 wbs_dat_o[17]
port 523 nsew signal output
rlabel metal3 s 39200 81064 40000 81184 6 wbs_dat_o[18]
port 524 nsew signal output
rlabel metal3 s 39200 81608 40000 81728 6 wbs_dat_o[19]
port 525 nsew signal output
rlabel metal3 s 39200 71816 40000 71936 6 wbs_dat_o[1]
port 526 nsew signal output
rlabel metal3 s 39200 82152 40000 82272 6 wbs_dat_o[20]
port 527 nsew signal output
rlabel metal3 s 39200 82696 40000 82816 6 wbs_dat_o[21]
port 528 nsew signal output
rlabel metal3 s 39200 83240 40000 83360 6 wbs_dat_o[22]
port 529 nsew signal output
rlabel metal3 s 39200 83784 40000 83904 6 wbs_dat_o[23]
port 530 nsew signal output
rlabel metal3 s 39200 84328 40000 84448 6 wbs_dat_o[24]
port 531 nsew signal output
rlabel metal3 s 39200 84872 40000 84992 6 wbs_dat_o[25]
port 532 nsew signal output
rlabel metal3 s 39200 85416 40000 85536 6 wbs_dat_o[26]
port 533 nsew signal output
rlabel metal3 s 39200 85960 40000 86080 6 wbs_dat_o[27]
port 534 nsew signal output
rlabel metal3 s 39200 86504 40000 86624 6 wbs_dat_o[28]
port 535 nsew signal output
rlabel metal3 s 39200 87048 40000 87168 6 wbs_dat_o[29]
port 536 nsew signal output
rlabel metal3 s 39200 72360 40000 72480 6 wbs_dat_o[2]
port 537 nsew signal output
rlabel metal3 s 39200 87592 40000 87712 6 wbs_dat_o[30]
port 538 nsew signal output
rlabel metal3 s 39200 88136 40000 88256 6 wbs_dat_o[31]
port 539 nsew signal output
rlabel metal3 s 39200 72904 40000 73024 6 wbs_dat_o[3]
port 540 nsew signal output
rlabel metal3 s 39200 73448 40000 73568 6 wbs_dat_o[4]
port 541 nsew signal output
rlabel metal3 s 39200 73992 40000 74112 6 wbs_dat_o[5]
port 542 nsew signal output
rlabel metal3 s 39200 74536 40000 74656 6 wbs_dat_o[6]
port 543 nsew signal output
rlabel metal3 s 39200 75080 40000 75200 6 wbs_dat_o[7]
port 544 nsew signal output
rlabel metal3 s 39200 75624 40000 75744 6 wbs_dat_o[8]
port 545 nsew signal output
rlabel metal3 s 39200 76168 40000 76288 6 wbs_dat_o[9]
port 546 nsew signal output
rlabel metal3 s 0 93032 800 93152 6 wbs_stb_i
port 547 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 wbs_we_i
port 548 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 220000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7639056
string GDS_FILE /home/tholin/Desktop/ci2406-rej-pommedeterrible-tholin/openlane/Multiplexer/runs/24_06_02_17_40/results/signoff/multiplexer.magic.gds
string GDS_START 438344
<< end >>

