magic
tech sky130B
magscale 1 2
timestamp 1717501105
<< obsli1 >>
rect 1104 2159 37812 36465
<< obsm1 >>
rect 934 1300 37982 36496
<< metal2 >>
rect 1122 38200 1178 39000
rect 2870 38200 2926 39000
rect 4618 38200 4674 39000
rect 6366 38200 6422 39000
rect 8114 38200 8170 39000
rect 9862 38200 9918 39000
rect 11610 38200 11666 39000
rect 13358 38200 13414 39000
rect 15106 38200 15162 39000
rect 16854 38200 16910 39000
rect 18602 38200 18658 39000
rect 20350 38200 20406 39000
rect 22098 38200 22154 39000
rect 23846 38200 23902 39000
rect 25594 38200 25650 39000
rect 27342 38200 27398 39000
rect 29090 38200 29146 39000
rect 30838 38200 30894 39000
rect 32586 38200 32642 39000
rect 34334 38200 34390 39000
rect 36082 38200 36138 39000
rect 37830 38200 37886 39000
rect 1766 0 1822 800
rect 3238 0 3294 800
rect 4710 0 4766 800
rect 6182 0 6238 800
rect 7654 0 7710 800
rect 9126 0 9182 800
rect 10598 0 10654 800
rect 12070 0 12126 800
rect 13542 0 13598 800
rect 15014 0 15070 800
rect 16486 0 16542 800
rect 17958 0 18014 800
rect 19430 0 19486 800
rect 20902 0 20958 800
rect 22374 0 22430 800
rect 23846 0 23902 800
rect 25318 0 25374 800
rect 26790 0 26846 800
rect 28262 0 28318 800
rect 29734 0 29790 800
rect 31206 0 31262 800
rect 32678 0 32734 800
rect 34150 0 34206 800
rect 35622 0 35678 800
rect 37094 0 37150 800
<< obsm2 >>
rect 938 38144 1066 38298
rect 1234 38144 2814 38298
rect 2982 38144 4562 38298
rect 4730 38144 6310 38298
rect 6478 38144 8058 38298
rect 8226 38144 9806 38298
rect 9974 38144 11554 38298
rect 11722 38144 13302 38298
rect 13470 38144 15050 38298
rect 15218 38144 16798 38298
rect 16966 38144 18546 38298
rect 18714 38144 20294 38298
rect 20462 38144 22042 38298
rect 22210 38144 23790 38298
rect 23958 38144 25538 38298
rect 25706 38144 27286 38298
rect 27454 38144 29034 38298
rect 29202 38144 30782 38298
rect 30950 38144 32530 38298
rect 32698 38144 34278 38298
rect 34446 38144 36026 38298
rect 36194 38144 37774 38298
rect 37942 38144 37978 38298
rect 938 856 37978 38144
rect 938 575 1710 856
rect 1878 575 3182 856
rect 3350 575 4654 856
rect 4822 575 6126 856
rect 6294 575 7598 856
rect 7766 575 9070 856
rect 9238 575 10542 856
rect 10710 575 12014 856
rect 12182 575 13486 856
rect 13654 575 14958 856
rect 15126 575 16430 856
rect 16598 575 17902 856
rect 18070 575 19374 856
rect 19542 575 20846 856
rect 21014 575 22318 856
rect 22486 575 23790 856
rect 23958 575 25262 856
rect 25430 575 26734 856
rect 26902 575 28206 856
rect 28374 575 29678 856
rect 29846 575 31150 856
rect 31318 575 32622 856
rect 32790 575 34094 856
rect 34262 575 35566 856
rect 35734 575 37038 856
rect 37206 575 37978 856
<< metal3 >>
rect 38200 38088 39000 38208
rect 0 36456 800 36576
rect 38200 36456 39000 36576
rect 0 34824 800 34944
rect 38200 34824 39000 34944
rect 0 33192 800 33312
rect 38200 33192 39000 33312
rect 0 31560 800 31680
rect 38200 31560 39000 31680
rect 0 29928 800 30048
rect 38200 29928 39000 30048
rect 0 28296 800 28416
rect 38200 28296 39000 28416
rect 0 26664 800 26784
rect 38200 26664 39000 26784
rect 0 25032 800 25152
rect 38200 25032 39000 25152
rect 0 23400 800 23520
rect 38200 23400 39000 23520
rect 0 21768 800 21888
rect 38200 21768 39000 21888
rect 0 20136 800 20256
rect 38200 20136 39000 20256
rect 0 18504 800 18624
rect 38200 18504 39000 18624
rect 0 16872 800 16992
rect 38200 16872 39000 16992
rect 0 15240 800 15360
rect 38200 15240 39000 15360
rect 0 13608 800 13728
rect 38200 13608 39000 13728
rect 0 11976 800 12096
rect 38200 11976 39000 12096
rect 0 10344 800 10464
rect 38200 10344 39000 10464
rect 0 8712 800 8832
rect 38200 8712 39000 8832
rect 0 7080 800 7200
rect 38200 7080 39000 7200
rect 0 5448 800 5568
rect 38200 5448 39000 5568
rect 0 3816 800 3936
rect 38200 3816 39000 3936
rect 0 2184 800 2304
rect 38200 2184 39000 2304
rect 38200 552 39000 672
<< obsm3 >>
rect 798 38008 38120 38181
rect 798 36656 38200 38008
rect 880 36376 38120 36656
rect 798 35024 38200 36376
rect 880 34744 38120 35024
rect 798 33392 38200 34744
rect 880 33112 38120 33392
rect 798 31760 38200 33112
rect 880 31480 38120 31760
rect 798 30128 38200 31480
rect 880 29848 38120 30128
rect 798 28496 38200 29848
rect 880 28216 38120 28496
rect 798 26864 38200 28216
rect 880 26584 38120 26864
rect 798 25232 38200 26584
rect 880 24952 38120 25232
rect 798 23600 38200 24952
rect 880 23320 38120 23600
rect 798 21968 38200 23320
rect 880 21688 38120 21968
rect 798 20336 38200 21688
rect 880 20056 38120 20336
rect 798 18704 38200 20056
rect 880 18424 38120 18704
rect 798 17072 38200 18424
rect 880 16792 38120 17072
rect 798 15440 38200 16792
rect 880 15160 38120 15440
rect 798 13808 38200 15160
rect 880 13528 38120 13808
rect 798 12176 38200 13528
rect 880 11896 38120 12176
rect 798 10544 38200 11896
rect 880 10264 38120 10544
rect 798 8912 38200 10264
rect 880 8632 38120 8912
rect 798 7280 38200 8632
rect 880 7000 38120 7280
rect 798 5648 38200 7000
rect 880 5368 38120 5648
rect 798 4016 38200 5368
rect 880 3736 38120 4016
rect 798 2384 38200 3736
rect 880 2104 38120 2384
rect 798 752 38200 2104
rect 798 579 38120 752
<< metal4 >>
rect 4208 2128 4528 36496
rect 19568 2128 19888 36496
rect 34928 2128 35248 36496
<< labels >>
rlabel metal2 s 1766 0 1822 800 6 irq[0]
port 1 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 irq[1]
port 2 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 irq[2]
port 3 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 la_data_out[0]
port 4 nsew signal output
rlabel metal2 s 2870 38200 2926 39000 6 la_data_out[10]
port 5 nsew signal output
rlabel metal2 s 4618 38200 4674 39000 6 la_data_out[11]
port 6 nsew signal output
rlabel metal2 s 6366 38200 6422 39000 6 la_data_out[12]
port 7 nsew signal output
rlabel metal2 s 8114 38200 8170 39000 6 la_data_out[13]
port 8 nsew signal output
rlabel metal2 s 9862 38200 9918 39000 6 la_data_out[14]
port 9 nsew signal output
rlabel metal2 s 11610 38200 11666 39000 6 la_data_out[15]
port 10 nsew signal output
rlabel metal2 s 13358 38200 13414 39000 6 la_data_out[16]
port 11 nsew signal output
rlabel metal2 s 15106 38200 15162 39000 6 la_data_out[17]
port 12 nsew signal output
rlabel metal2 s 16854 38200 16910 39000 6 la_data_out[18]
port 13 nsew signal output
rlabel metal2 s 18602 38200 18658 39000 6 la_data_out[19]
port 14 nsew signal output
rlabel metal2 s 1122 38200 1178 39000 6 la_data_out[1]
port 15 nsew signal output
rlabel metal2 s 22098 38200 22154 39000 6 la_data_out[20]
port 16 nsew signal output
rlabel metal2 s 23846 38200 23902 39000 6 la_data_out[21]
port 17 nsew signal output
rlabel metal2 s 25594 38200 25650 39000 6 la_data_out[22]
port 18 nsew signal output
rlabel metal2 s 27342 38200 27398 39000 6 la_data_out[23]
port 19 nsew signal output
rlabel metal2 s 29090 38200 29146 39000 6 la_data_out[24]
port 20 nsew signal output
rlabel metal2 s 30838 38200 30894 39000 6 la_data_out[25]
port 21 nsew signal output
rlabel metal2 s 32586 38200 32642 39000 6 la_data_out[26]
port 22 nsew signal output
rlabel metal2 s 34334 38200 34390 39000 6 la_data_out[27]
port 23 nsew signal output
rlabel metal2 s 36082 38200 36138 39000 6 la_data_out[28]
port 24 nsew signal output
rlabel metal2 s 37830 38200 37886 39000 6 la_data_out[29]
port 25 nsew signal output
rlabel metal2 s 20350 38200 20406 39000 6 la_data_out[2]
port 26 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 la_data_out[30]
port 27 nsew signal output
rlabel metal2 s 25318 0 25374 800 6 la_data_out[31]
port 28 nsew signal output
rlabel metal2 s 26790 0 26846 800 6 la_data_out[32]
port 29 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 la_data_out[33]
port 30 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 la_data_out[34]
port 31 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 la_data_out[35]
port 32 nsew signal output
rlabel metal2 s 32678 0 32734 800 6 la_data_out[36]
port 33 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 la_data_out[37]
port 34 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 la_data_out[38]
port 35 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 la_data_out[39]
port 36 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 la_data_out[3]
port 37 nsew signal output
rlabel metal3 s 38200 5448 39000 5568 6 la_data_out[40]
port 38 nsew signal output
rlabel metal3 s 38200 7080 39000 7200 6 la_data_out[41]
port 39 nsew signal output
rlabel metal3 s 38200 8712 39000 8832 6 la_data_out[42]
port 40 nsew signal output
rlabel metal3 s 38200 10344 39000 10464 6 la_data_out[43]
port 41 nsew signal output
rlabel metal3 s 38200 11976 39000 12096 6 la_data_out[44]
port 42 nsew signal output
rlabel metal3 s 38200 13608 39000 13728 6 la_data_out[45]
port 43 nsew signal output
rlabel metal3 s 38200 15240 39000 15360 6 la_data_out[46]
port 44 nsew signal output
rlabel metal3 s 38200 16872 39000 16992 6 la_data_out[47]
port 45 nsew signal output
rlabel metal3 s 38200 18504 39000 18624 6 la_data_out[48]
port 46 nsew signal output
rlabel metal3 s 38200 20136 39000 20256 6 la_data_out[49]
port 47 nsew signal output
rlabel metal3 s 38200 3816 39000 3936 6 la_data_out[4]
port 48 nsew signal output
rlabel metal3 s 38200 23400 39000 23520 6 la_data_out[50]
port 49 nsew signal output
rlabel metal3 s 38200 25032 39000 25152 6 la_data_out[51]
port 50 nsew signal output
rlabel metal3 s 38200 26664 39000 26784 6 la_data_out[52]
port 51 nsew signal output
rlabel metal3 s 38200 28296 39000 28416 6 la_data_out[53]
port 52 nsew signal output
rlabel metal3 s 38200 29928 39000 30048 6 la_data_out[54]
port 53 nsew signal output
rlabel metal3 s 38200 31560 39000 31680 6 la_data_out[55]
port 54 nsew signal output
rlabel metal3 s 38200 33192 39000 33312 6 la_data_out[56]
port 55 nsew signal output
rlabel metal3 s 38200 34824 39000 34944 6 la_data_out[57]
port 56 nsew signal output
rlabel metal3 s 38200 36456 39000 36576 6 la_data_out[58]
port 57 nsew signal output
rlabel metal3 s 38200 38088 39000 38208 6 la_data_out[59]
port 58 nsew signal output
rlabel metal3 s 38200 21768 39000 21888 6 la_data_out[5]
port 59 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 la_data_out[60]
port 60 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 la_data_out[61]
port 61 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 la_data_out[62]
port 62 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 la_data_out[63]
port 63 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 la_data_out[64]
port 64 nsew signal output
rlabel metal2 s 15014 0 15070 800 6 la_data_out[65]
port 65 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 la_data_out[66]
port 66 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 la_data_out[67]
port 67 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 la_data_out[68]
port 68 nsew signal output
rlabel metal2 s 20902 0 20958 800 6 la_data_out[69]
port 69 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 la_data_out[6]
port 70 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 la_data_out[70]
port 71 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 la_data_out[71]
port 72 nsew signal output
rlabel metal3 s 0 21768 800 21888 6 la_data_out[72]
port 73 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 la_data_out[73]
port 74 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 la_data_out[74]
port 75 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 la_data_out[75]
port 76 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 la_data_out[76]
port 77 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 la_data_out[77]
port 78 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 la_data_out[78]
port 79 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 la_data_out[79]
port 80 nsew signal output
rlabel metal3 s 0 16872 800 16992 6 la_data_out[7]
port 81 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 la_data_out[80]
port 82 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 la_data_out[81]
port 83 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 la_data_out[82]
port 84 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 la_data_out[83]
port 85 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 la_data_out[84]
port 86 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 la_data_out[85]
port 87 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 la_data_out[86]
port 88 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 la_data_out[87]
port 89 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 la_data_out[8]
port 90 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 la_data_out[9]
port 91 nsew signal output
rlabel metal4 s 4208 2128 4528 36496 6 vccd1
port 92 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 36496 6 vccd1
port 92 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 36496 6 vssd1
port 93 nsew ground bidirectional
rlabel metal3 s 38200 552 39000 672 6 wb_clk_i
port 94 nsew signal input
rlabel metal3 s 38200 2184 39000 2304 6 wb_rst_i
port 95 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 39000 39000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1359912
string GDS_FILE /home/lucah/Desktop/ci2406-rej-pommedeterrible-tholin/openlane/TieUnused/runs/24_06_04_13_35/results/signoff/unused_tie.magic.gds
string GDS_START 108930
<< end >>

