magic
tech sky130B
magscale 1 2
timestamp 1717507627
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 934 348 59970 58200
<< metal2 >>
rect 938 59200 994 60000
rect 2594 59200 2650 60000
rect 4250 59200 4306 60000
rect 5906 59200 5962 60000
rect 7562 59200 7618 60000
rect 9218 59200 9274 60000
rect 10874 59200 10930 60000
rect 12530 59200 12586 60000
rect 14186 59200 14242 60000
rect 15842 59200 15898 60000
rect 17498 59200 17554 60000
rect 19154 59200 19210 60000
rect 20810 59200 20866 60000
rect 22466 59200 22522 60000
rect 24122 59200 24178 60000
rect 25778 59200 25834 60000
rect 27434 59200 27490 60000
rect 29090 59200 29146 60000
rect 30746 59200 30802 60000
rect 32402 59200 32458 60000
rect 34058 59200 34114 60000
rect 35714 59200 35770 60000
rect 37370 59200 37426 60000
rect 39026 59200 39082 60000
rect 40682 59200 40738 60000
rect 42338 59200 42394 60000
rect 43994 59200 44050 60000
rect 45650 59200 45706 60000
rect 47306 59200 47362 60000
rect 48962 59200 49018 60000
rect 50618 59200 50674 60000
rect 52274 59200 52330 60000
rect 53930 59200 53986 60000
rect 55586 59200 55642 60000
rect 57242 59200 57298 60000
rect 58898 59200 58954 60000
rect 938 0 994 800
rect 2594 0 2650 800
rect 4250 0 4306 800
rect 5906 0 5962 800
rect 7562 0 7618 800
rect 9218 0 9274 800
rect 10874 0 10930 800
rect 12530 0 12586 800
rect 14186 0 14242 800
rect 15842 0 15898 800
rect 17498 0 17554 800
rect 19154 0 19210 800
rect 20810 0 20866 800
rect 22466 0 22522 800
rect 24122 0 24178 800
rect 25778 0 25834 800
rect 27434 0 27490 800
rect 29090 0 29146 800
rect 30746 0 30802 800
rect 32402 0 32458 800
rect 34058 0 34114 800
rect 35714 0 35770 800
rect 37370 0 37426 800
rect 39026 0 39082 800
rect 40682 0 40738 800
rect 42338 0 42394 800
rect 43994 0 44050 800
rect 45650 0 45706 800
rect 47306 0 47362 800
rect 48962 0 49018 800
rect 50618 0 50674 800
rect 52274 0 52330 800
rect 53930 0 53986 800
rect 55586 0 55642 800
rect 57242 0 57298 800
rect 58898 0 58954 800
<< obsm2 >>
rect 1050 59144 2538 59242
rect 2706 59144 4194 59242
rect 4362 59144 5850 59242
rect 6018 59144 7506 59242
rect 7674 59144 9162 59242
rect 9330 59144 10818 59242
rect 10986 59144 12474 59242
rect 12642 59144 14130 59242
rect 14298 59144 15786 59242
rect 15954 59144 17442 59242
rect 17610 59144 19098 59242
rect 19266 59144 20754 59242
rect 20922 59144 22410 59242
rect 22578 59144 24066 59242
rect 24234 59144 25722 59242
rect 25890 59144 27378 59242
rect 27546 59144 29034 59242
rect 29202 59144 30690 59242
rect 30858 59144 32346 59242
rect 32514 59144 34002 59242
rect 34170 59144 35658 59242
rect 35826 59144 37314 59242
rect 37482 59144 38970 59242
rect 39138 59144 40626 59242
rect 40794 59144 42282 59242
rect 42450 59144 43938 59242
rect 44106 59144 45594 59242
rect 45762 59144 47250 59242
rect 47418 59144 48906 59242
rect 49074 59144 50562 59242
rect 50730 59144 52218 59242
rect 52386 59144 53874 59242
rect 54042 59144 55530 59242
rect 55698 59144 57186 59242
rect 57354 59144 58842 59242
rect 59010 59144 59966 59242
rect 938 856 59966 59144
rect 1050 303 2538 856
rect 2706 303 4194 856
rect 4362 303 5850 856
rect 6018 303 7506 856
rect 7674 303 9162 856
rect 9330 303 10818 856
rect 10986 303 12474 856
rect 12642 303 14130 856
rect 14298 303 15786 856
rect 15954 303 17442 856
rect 17610 303 19098 856
rect 19266 303 20754 856
rect 20922 303 22410 856
rect 22578 303 24066 856
rect 24234 303 25722 856
rect 25890 303 27378 856
rect 27546 303 29034 856
rect 29202 303 30690 856
rect 30858 303 32346 856
rect 32514 303 34002 856
rect 34170 303 35658 856
rect 35826 303 37314 856
rect 37482 303 38970 856
rect 39138 303 40626 856
rect 40794 303 42282 856
rect 42450 303 43938 856
rect 44106 303 45594 856
rect 45762 303 47250 856
rect 47418 303 48906 856
rect 49074 303 50562 856
rect 50730 303 52218 856
rect 52386 303 53874 856
rect 54042 303 55530 856
rect 55698 303 57186 856
rect 57354 303 58842 856
rect 59010 303 59966 856
<< metal3 >>
rect 59200 58488 60000 58608
rect 59200 56856 60000 56976
rect 59200 55224 60000 55344
rect 59200 53592 60000 53712
rect 59200 51960 60000 52080
rect 59200 50328 60000 50448
rect 59200 48696 60000 48816
rect 59200 47064 60000 47184
rect 59200 45432 60000 45552
rect 0 44888 800 45008
rect 59200 43800 60000 43920
rect 59200 42168 60000 42288
rect 59200 40536 60000 40656
rect 59200 38904 60000 39024
rect 59200 37272 60000 37392
rect 59200 35640 60000 35760
rect 59200 34008 60000 34128
rect 59200 32376 60000 32496
rect 59200 30744 60000 30864
rect 59200 29112 60000 29232
rect 59200 27480 60000 27600
rect 59200 25848 60000 25968
rect 59200 24216 60000 24336
rect 59200 22584 60000 22704
rect 59200 20952 60000 21072
rect 59200 19320 60000 19440
rect 59200 17688 60000 17808
rect 59200 16056 60000 16176
rect 0 14968 800 15088
rect 59200 14424 60000 14544
rect 59200 12792 60000 12912
rect 59200 11160 60000 11280
rect 59200 9528 60000 9648
rect 59200 7896 60000 8016
rect 59200 6264 60000 6384
rect 59200 4632 60000 4752
rect 59200 3000 60000 3120
rect 59200 1368 60000 1488
<< obsm3 >>
rect 800 58408 59120 58581
rect 800 57056 59971 58408
rect 800 56776 59120 57056
rect 800 55424 59971 56776
rect 800 55144 59120 55424
rect 800 53792 59971 55144
rect 800 53512 59120 53792
rect 800 52160 59971 53512
rect 800 51880 59120 52160
rect 800 50528 59971 51880
rect 800 50248 59120 50528
rect 800 48896 59971 50248
rect 800 48616 59120 48896
rect 800 47264 59971 48616
rect 800 46984 59120 47264
rect 800 45632 59971 46984
rect 800 45352 59120 45632
rect 800 45088 59971 45352
rect 880 44808 59971 45088
rect 800 44000 59971 44808
rect 800 43720 59120 44000
rect 800 42368 59971 43720
rect 800 42088 59120 42368
rect 800 40736 59971 42088
rect 800 40456 59120 40736
rect 800 39104 59971 40456
rect 800 38824 59120 39104
rect 800 37472 59971 38824
rect 800 37192 59120 37472
rect 800 35840 59971 37192
rect 800 35560 59120 35840
rect 800 34208 59971 35560
rect 800 33928 59120 34208
rect 800 32576 59971 33928
rect 800 32296 59120 32576
rect 800 30944 59971 32296
rect 800 30664 59120 30944
rect 800 29312 59971 30664
rect 800 29032 59120 29312
rect 800 27680 59971 29032
rect 800 27400 59120 27680
rect 800 26048 59971 27400
rect 800 25768 59120 26048
rect 800 24416 59971 25768
rect 800 24136 59120 24416
rect 800 22784 59971 24136
rect 800 22504 59120 22784
rect 800 21152 59971 22504
rect 800 20872 59120 21152
rect 800 19520 59971 20872
rect 800 19240 59120 19520
rect 800 17888 59971 19240
rect 800 17608 59120 17888
rect 800 16256 59971 17608
rect 800 15976 59120 16256
rect 800 15168 59971 15976
rect 880 14888 59971 15168
rect 800 14624 59971 14888
rect 800 14344 59120 14624
rect 800 12992 59971 14344
rect 800 12712 59120 12992
rect 800 11360 59971 12712
rect 800 11080 59120 11360
rect 800 9728 59971 11080
rect 800 9448 59120 9728
rect 800 8096 59971 9448
rect 800 7816 59120 8096
rect 800 6464 59971 7816
rect 800 6184 59120 6464
rect 800 4832 59971 6184
rect 800 4552 59120 4832
rect 800 3200 59971 4552
rect 800 2920 59120 3200
rect 800 1568 59971 2920
rect 800 1288 59120 1568
rect 800 307 59971 1288
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< obsm4 >>
rect 9811 57792 58453 58309
rect 9811 2048 19488 57792
rect 19968 2048 34848 57792
rect 35328 2048 50208 57792
rect 50688 2048 58453 57792
rect 9811 307 58453 2048
<< labels >>
rlabel metal2 s 938 59200 994 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 17498 59200 17554 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 19154 59200 19210 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 20810 59200 20866 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 22466 59200 22522 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 24122 59200 24178 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 25778 59200 25834 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 27434 59200 27490 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 29090 59200 29146 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 30746 59200 30802 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 32402 59200 32458 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2594 59200 2650 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 34058 59200 34114 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 35714 59200 35770 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 37370 59200 37426 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 39026 59200 39082 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 40682 59200 40738 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 42338 59200 42394 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 43994 59200 44050 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 45650 59200 45706 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 47306 59200 47362 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 48962 59200 49018 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 4250 59200 4306 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 50618 59200 50674 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 52274 59200 52330 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 53930 59200 53986 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 55586 59200 55642 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 57242 59200 57298 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 58898 59200 58954 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 5906 59200 5962 60000 6 io_in[3]
port 30 nsew signal input
rlabel metal2 s 7562 59200 7618 60000 6 io_in[4]
port 31 nsew signal input
rlabel metal2 s 9218 59200 9274 60000 6 io_in[5]
port 32 nsew signal input
rlabel metal2 s 10874 59200 10930 60000 6 io_in[6]
port 33 nsew signal input
rlabel metal2 s 12530 59200 12586 60000 6 io_in[7]
port 34 nsew signal input
rlabel metal2 s 14186 59200 14242 60000 6 io_in[8]
port 35 nsew signal input
rlabel metal2 s 15842 59200 15898 60000 6 io_in[9]
port 36 nsew signal input
rlabel metal2 s 938 0 994 800 6 io_oeb[0]
port 37 nsew signal output
rlabel metal2 s 17498 0 17554 800 6 io_oeb[10]
port 38 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 io_oeb[11]
port 39 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 io_oeb[12]
port 40 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 io_oeb[13]
port 41 nsew signal output
rlabel metal2 s 24122 0 24178 800 6 io_oeb[14]
port 42 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 io_oeb[15]
port 43 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 io_oeb[16]
port 44 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 io_oeb[17]
port 45 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 io_oeb[18]
port 46 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 io_oeb[19]
port 47 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 io_oeb[1]
port 48 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 io_oeb[20]
port 49 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 io_oeb[21]
port 50 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 io_oeb[22]
port 51 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 io_oeb[23]
port 52 nsew signal output
rlabel metal2 s 40682 0 40738 800 6 io_oeb[24]
port 53 nsew signal output
rlabel metal2 s 42338 0 42394 800 6 io_oeb[25]
port 54 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 io_oeb[26]
port 55 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 io_oeb[27]
port 56 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 io_oeb[28]
port 57 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 io_oeb[29]
port 58 nsew signal output
rlabel metal2 s 4250 0 4306 800 6 io_oeb[2]
port 59 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 io_oeb[30]
port 60 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 io_oeb[31]
port 61 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 io_oeb[32]
port 62 nsew signal output
rlabel metal2 s 55586 0 55642 800 6 io_oeb[33]
port 63 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 io_oeb[34]
port 64 nsew signal output
rlabel metal2 s 58898 0 58954 800 6 io_oeb[35]
port 65 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 io_oeb[3]
port 66 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 io_oeb[4]
port 67 nsew signal output
rlabel metal2 s 9218 0 9274 800 6 io_oeb[5]
port 68 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 io_oeb[6]
port 69 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 io_oeb[7]
port 70 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 io_oeb[8]
port 71 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 io_oeb[9]
port 72 nsew signal output
rlabel metal3 s 59200 1368 60000 1488 6 io_out[0]
port 73 nsew signal output
rlabel metal3 s 59200 17688 60000 17808 6 io_out[10]
port 74 nsew signal output
rlabel metal3 s 59200 19320 60000 19440 6 io_out[11]
port 75 nsew signal output
rlabel metal3 s 59200 20952 60000 21072 6 io_out[12]
port 76 nsew signal output
rlabel metal3 s 59200 22584 60000 22704 6 io_out[13]
port 77 nsew signal output
rlabel metal3 s 59200 24216 60000 24336 6 io_out[14]
port 78 nsew signal output
rlabel metal3 s 59200 25848 60000 25968 6 io_out[15]
port 79 nsew signal output
rlabel metal3 s 59200 27480 60000 27600 6 io_out[16]
port 80 nsew signal output
rlabel metal3 s 59200 29112 60000 29232 6 io_out[17]
port 81 nsew signal output
rlabel metal3 s 59200 30744 60000 30864 6 io_out[18]
port 82 nsew signal output
rlabel metal3 s 59200 32376 60000 32496 6 io_out[19]
port 83 nsew signal output
rlabel metal3 s 59200 3000 60000 3120 6 io_out[1]
port 84 nsew signal output
rlabel metal3 s 59200 34008 60000 34128 6 io_out[20]
port 85 nsew signal output
rlabel metal3 s 59200 35640 60000 35760 6 io_out[21]
port 86 nsew signal output
rlabel metal3 s 59200 37272 60000 37392 6 io_out[22]
port 87 nsew signal output
rlabel metal3 s 59200 38904 60000 39024 6 io_out[23]
port 88 nsew signal output
rlabel metal3 s 59200 40536 60000 40656 6 io_out[24]
port 89 nsew signal output
rlabel metal3 s 59200 42168 60000 42288 6 io_out[25]
port 90 nsew signal output
rlabel metal3 s 59200 43800 60000 43920 6 io_out[26]
port 91 nsew signal output
rlabel metal3 s 59200 45432 60000 45552 6 io_out[27]
port 92 nsew signal output
rlabel metal3 s 59200 47064 60000 47184 6 io_out[28]
port 93 nsew signal output
rlabel metal3 s 59200 48696 60000 48816 6 io_out[29]
port 94 nsew signal output
rlabel metal3 s 59200 4632 60000 4752 6 io_out[2]
port 95 nsew signal output
rlabel metal3 s 59200 50328 60000 50448 6 io_out[30]
port 96 nsew signal output
rlabel metal3 s 59200 51960 60000 52080 6 io_out[31]
port 97 nsew signal output
rlabel metal3 s 59200 53592 60000 53712 6 io_out[32]
port 98 nsew signal output
rlabel metal3 s 59200 55224 60000 55344 6 io_out[33]
port 99 nsew signal output
rlabel metal3 s 59200 56856 60000 56976 6 io_out[34]
port 100 nsew signal output
rlabel metal3 s 59200 58488 60000 58608 6 io_out[35]
port 101 nsew signal output
rlabel metal3 s 59200 6264 60000 6384 6 io_out[3]
port 102 nsew signal output
rlabel metal3 s 59200 7896 60000 8016 6 io_out[4]
port 103 nsew signal output
rlabel metal3 s 59200 9528 60000 9648 6 io_out[5]
port 104 nsew signal output
rlabel metal3 s 59200 11160 60000 11280 6 io_out[6]
port 105 nsew signal output
rlabel metal3 s 59200 12792 60000 12912 6 io_out[7]
port 106 nsew signal output
rlabel metal3 s 59200 14424 60000 14544 6 io_out[8]
port 107 nsew signal output
rlabel metal3 s 59200 16056 60000 16176 6 io_out[9]
port 108 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 rst_n
port 109 nsew signal input
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 111 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 111 nsew ground bidirectional
rlabel metal3 s 0 14968 800 15088 6 wb_clk_i
port 112 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 16341350
string GDS_FILE /home/lucah/Desktop/ci2406-rej-pommedeterrible-tholin/openlane/Z80/runs/24_06_04_14_37/results/signoff/ci2406_z80.magic.gds
string GDS_START 1303134
<< end >>

