magic
tech sky130A
magscale 1 2
timestamp 1716587709
<< obsli1 >>
rect 1104 2159 48852 52785
<< obsm1 >>
rect 750 2128 49114 52816
<< metal2 >>
rect 754 54200 810 55000
rect 2134 54200 2190 55000
rect 3514 54200 3570 55000
rect 4894 54200 4950 55000
rect 6274 54200 6330 55000
rect 7654 54200 7710 55000
rect 9034 54200 9090 55000
rect 10414 54200 10470 55000
rect 11794 54200 11850 55000
rect 13174 54200 13230 55000
rect 14554 54200 14610 55000
rect 15934 54200 15990 55000
rect 17314 54200 17370 55000
rect 18694 54200 18750 55000
rect 20074 54200 20130 55000
rect 21454 54200 21510 55000
rect 22834 54200 22890 55000
rect 24214 54200 24270 55000
rect 25594 54200 25650 55000
rect 26974 54200 27030 55000
rect 28354 54200 28410 55000
rect 29734 54200 29790 55000
rect 31114 54200 31170 55000
rect 32494 54200 32550 55000
rect 33874 54200 33930 55000
rect 35254 54200 35310 55000
rect 36634 54200 36690 55000
rect 38014 54200 38070 55000
rect 39394 54200 39450 55000
rect 40774 54200 40830 55000
rect 42154 54200 42210 55000
rect 43534 54200 43590 55000
rect 44914 54200 44970 55000
rect 46294 54200 46350 55000
rect 47674 54200 47730 55000
rect 49054 54200 49110 55000
rect 754 0 810 800
rect 2134 0 2190 800
rect 3514 0 3570 800
rect 4894 0 4950 800
rect 6274 0 6330 800
rect 7654 0 7710 800
rect 9034 0 9090 800
rect 10414 0 10470 800
rect 11794 0 11850 800
rect 13174 0 13230 800
rect 14554 0 14610 800
rect 15934 0 15990 800
rect 17314 0 17370 800
rect 18694 0 18750 800
rect 20074 0 20130 800
rect 21454 0 21510 800
rect 22834 0 22890 800
rect 24214 0 24270 800
rect 25594 0 25650 800
rect 26974 0 27030 800
rect 28354 0 28410 800
rect 29734 0 29790 800
rect 31114 0 31170 800
rect 32494 0 32550 800
rect 33874 0 33930 800
rect 35254 0 35310 800
rect 36634 0 36690 800
rect 38014 0 38070 800
rect 39394 0 39450 800
rect 40774 0 40830 800
rect 42154 0 42210 800
rect 43534 0 43590 800
rect 44914 0 44970 800
rect 46294 0 46350 800
rect 47674 0 47730 800
rect 49054 0 49110 800
<< obsm2 >>
rect 866 54144 2078 54346
rect 2246 54144 3458 54346
rect 3626 54144 4838 54346
rect 5006 54144 6218 54346
rect 6386 54144 7598 54346
rect 7766 54144 8978 54346
rect 9146 54144 10358 54346
rect 10526 54144 11738 54346
rect 11906 54144 13118 54346
rect 13286 54144 14498 54346
rect 14666 54144 15878 54346
rect 16046 54144 17258 54346
rect 17426 54144 18638 54346
rect 18806 54144 20018 54346
rect 20186 54144 21398 54346
rect 21566 54144 22778 54346
rect 22946 54144 24158 54346
rect 24326 54144 25538 54346
rect 25706 54144 26918 54346
rect 27086 54144 28298 54346
rect 28466 54144 29678 54346
rect 29846 54144 31058 54346
rect 31226 54144 32438 54346
rect 32606 54144 33818 54346
rect 33986 54144 35198 54346
rect 35366 54144 36578 54346
rect 36746 54144 37958 54346
rect 38126 54144 39338 54346
rect 39506 54144 40718 54346
rect 40886 54144 42098 54346
rect 42266 54144 43478 54346
rect 43646 54144 44858 54346
rect 45026 54144 46238 54346
rect 46406 54144 47618 54346
rect 47786 54144 48998 54346
rect 756 856 49108 54144
rect 866 734 2078 856
rect 2246 734 3458 856
rect 3626 734 4838 856
rect 5006 734 6218 856
rect 6386 734 7598 856
rect 7766 734 8978 856
rect 9146 734 10358 856
rect 10526 734 11738 856
rect 11906 734 13118 856
rect 13286 734 14498 856
rect 14666 734 15878 856
rect 16046 734 17258 856
rect 17426 734 18638 856
rect 18806 734 20018 856
rect 20186 734 21398 856
rect 21566 734 22778 856
rect 22946 734 24158 856
rect 24326 734 25538 856
rect 25706 734 26918 856
rect 27086 734 28298 856
rect 28466 734 29678 856
rect 29846 734 31058 856
rect 31226 734 32438 856
rect 32606 734 33818 856
rect 33986 734 35198 856
rect 35366 734 36578 856
rect 36746 734 37958 856
rect 38126 734 39338 856
rect 39506 734 40718 856
rect 40886 734 42098 856
rect 42266 734 43478 856
rect 43646 734 44858 856
rect 45026 734 46238 856
rect 46406 734 47618 856
rect 47786 734 48998 856
<< metal3 >>
rect 49200 51144 50000 51264
rect 49200 49784 50000 49904
rect 49200 48424 50000 48544
rect 49200 47064 50000 47184
rect 49200 45704 50000 45824
rect 49200 44344 50000 44464
rect 49200 42984 50000 43104
rect 49200 41624 50000 41744
rect 0 41080 800 41200
rect 49200 40264 50000 40384
rect 49200 38904 50000 39024
rect 49200 37544 50000 37664
rect 49200 36184 50000 36304
rect 49200 34824 50000 34944
rect 49200 33464 50000 33584
rect 49200 32104 50000 32224
rect 49200 30744 50000 30864
rect 49200 29384 50000 29504
rect 49200 28024 50000 28144
rect 49200 26664 50000 26784
rect 49200 25304 50000 25424
rect 49200 23944 50000 24064
rect 49200 22584 50000 22704
rect 49200 21224 50000 21344
rect 49200 19864 50000 19984
rect 49200 18504 50000 18624
rect 49200 17144 50000 17264
rect 49200 15784 50000 15904
rect 49200 14424 50000 14544
rect 0 13608 800 13728
rect 49200 13064 50000 13184
rect 49200 11704 50000 11824
rect 49200 10344 50000 10464
rect 49200 8984 50000 9104
rect 49200 7624 50000 7744
rect 49200 6264 50000 6384
rect 49200 4904 50000 5024
rect 49200 3544 50000 3664
<< obsm3 >>
rect 800 51344 49200 52801
rect 800 51064 49120 51344
rect 800 49984 49200 51064
rect 800 49704 49120 49984
rect 800 48624 49200 49704
rect 800 48344 49120 48624
rect 800 47264 49200 48344
rect 800 46984 49120 47264
rect 800 45904 49200 46984
rect 800 45624 49120 45904
rect 800 44544 49200 45624
rect 800 44264 49120 44544
rect 800 43184 49200 44264
rect 800 42904 49120 43184
rect 800 41824 49200 42904
rect 800 41544 49120 41824
rect 800 41280 49200 41544
rect 880 41000 49200 41280
rect 800 40464 49200 41000
rect 800 40184 49120 40464
rect 800 39104 49200 40184
rect 800 38824 49120 39104
rect 800 37744 49200 38824
rect 800 37464 49120 37744
rect 800 36384 49200 37464
rect 800 36104 49120 36384
rect 800 35024 49200 36104
rect 800 34744 49120 35024
rect 800 33664 49200 34744
rect 800 33384 49120 33664
rect 800 32304 49200 33384
rect 800 32024 49120 32304
rect 800 30944 49200 32024
rect 800 30664 49120 30944
rect 800 29584 49200 30664
rect 800 29304 49120 29584
rect 800 28224 49200 29304
rect 800 27944 49120 28224
rect 800 26864 49200 27944
rect 800 26584 49120 26864
rect 800 25504 49200 26584
rect 800 25224 49120 25504
rect 800 24144 49200 25224
rect 800 23864 49120 24144
rect 800 22784 49200 23864
rect 800 22504 49120 22784
rect 800 21424 49200 22504
rect 800 21144 49120 21424
rect 800 20064 49200 21144
rect 800 19784 49120 20064
rect 800 18704 49200 19784
rect 800 18424 49120 18704
rect 800 17344 49200 18424
rect 800 17064 49120 17344
rect 800 15984 49200 17064
rect 800 15704 49120 15984
rect 800 14624 49200 15704
rect 800 14344 49120 14624
rect 800 13808 49200 14344
rect 880 13528 49200 13808
rect 800 13264 49200 13528
rect 800 12984 49120 13264
rect 800 11904 49200 12984
rect 800 11624 49120 11904
rect 800 10544 49200 11624
rect 800 10264 49120 10544
rect 800 9184 49200 10264
rect 800 8904 49120 9184
rect 800 7824 49200 8904
rect 800 7544 49120 7824
rect 800 6464 49200 7544
rect 800 6184 49120 6464
rect 800 5104 49200 6184
rect 800 4824 49120 5104
rect 800 3744 49200 4824
rect 800 3464 49120 3744
rect 800 2143 49200 3464
<< metal4 >>
rect 4208 2128 4528 52816
rect 19568 2128 19888 52816
rect 34928 2128 35248 52816
<< obsm4 >>
rect 5579 2347 19488 52597
rect 19968 2347 34848 52597
rect 35328 2347 45573 52597
<< labels >>
rlabel metal2 s 754 54200 810 55000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 14554 54200 14610 55000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 15934 54200 15990 55000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 17314 54200 17370 55000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 18694 54200 18750 55000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 20074 54200 20130 55000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 21454 54200 21510 55000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 22834 54200 22890 55000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 24214 54200 24270 55000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 25594 54200 25650 55000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 26974 54200 27030 55000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 2134 54200 2190 55000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 28354 54200 28410 55000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 29734 54200 29790 55000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 31114 54200 31170 55000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 32494 54200 32550 55000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 33874 54200 33930 55000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 35254 54200 35310 55000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 36634 54200 36690 55000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 38014 54200 38070 55000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 39394 54200 39450 55000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 40774 54200 40830 55000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 3514 54200 3570 55000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 42154 54200 42210 55000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 43534 54200 43590 55000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 44914 54200 44970 55000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 46294 54200 46350 55000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 47674 54200 47730 55000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 49054 54200 49110 55000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 4894 54200 4950 55000 6 io_in[3]
port 30 nsew signal input
rlabel metal2 s 6274 54200 6330 55000 6 io_in[4]
port 31 nsew signal input
rlabel metal2 s 7654 54200 7710 55000 6 io_in[5]
port 32 nsew signal input
rlabel metal2 s 9034 54200 9090 55000 6 io_in[6]
port 33 nsew signal input
rlabel metal2 s 10414 54200 10470 55000 6 io_in[7]
port 34 nsew signal input
rlabel metal2 s 11794 54200 11850 55000 6 io_in[8]
port 35 nsew signal input
rlabel metal2 s 13174 54200 13230 55000 6 io_in[9]
port 36 nsew signal input
rlabel metal2 s 754 0 810 800 6 io_oeb[0]
port 37 nsew signal output
rlabel metal2 s 14554 0 14610 800 6 io_oeb[10]
port 38 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 io_oeb[11]
port 39 nsew signal output
rlabel metal2 s 17314 0 17370 800 6 io_oeb[12]
port 40 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 io_oeb[13]
port 41 nsew signal output
rlabel metal2 s 20074 0 20130 800 6 io_oeb[14]
port 42 nsew signal output
rlabel metal2 s 21454 0 21510 800 6 io_oeb[15]
port 43 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 io_oeb[16]
port 44 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 io_oeb[17]
port 45 nsew signal output
rlabel metal2 s 25594 0 25650 800 6 io_oeb[18]
port 46 nsew signal output
rlabel metal2 s 26974 0 27030 800 6 io_oeb[19]
port 47 nsew signal output
rlabel metal2 s 2134 0 2190 800 6 io_oeb[1]
port 48 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 io_oeb[20]
port 49 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 io_oeb[21]
port 50 nsew signal output
rlabel metal2 s 31114 0 31170 800 6 io_oeb[22]
port 51 nsew signal output
rlabel metal2 s 32494 0 32550 800 6 io_oeb[23]
port 52 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 io_oeb[24]
port 53 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 io_oeb[25]
port 54 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 io_oeb[26]
port 55 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 io_oeb[27]
port 56 nsew signal output
rlabel metal2 s 39394 0 39450 800 6 io_oeb[28]
port 57 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 io_oeb[29]
port 58 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 io_oeb[2]
port 59 nsew signal output
rlabel metal2 s 42154 0 42210 800 6 io_oeb[30]
port 60 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 io_oeb[31]
port 61 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 io_oeb[32]
port 62 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 io_oeb[33]
port 63 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 io_oeb[34]
port 64 nsew signal output
rlabel metal2 s 49054 0 49110 800 6 io_oeb[35]
port 65 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 io_oeb[3]
port 66 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 io_oeb[4]
port 67 nsew signal output
rlabel metal2 s 7654 0 7710 800 6 io_oeb[5]
port 68 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 io_oeb[6]
port 69 nsew signal output
rlabel metal2 s 10414 0 10470 800 6 io_oeb[7]
port 70 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 io_oeb[8]
port 71 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 io_oeb[9]
port 72 nsew signal output
rlabel metal3 s 49200 3544 50000 3664 6 io_out[0]
port 73 nsew signal output
rlabel metal3 s 49200 17144 50000 17264 6 io_out[10]
port 74 nsew signal output
rlabel metal3 s 49200 18504 50000 18624 6 io_out[11]
port 75 nsew signal output
rlabel metal3 s 49200 19864 50000 19984 6 io_out[12]
port 76 nsew signal output
rlabel metal3 s 49200 21224 50000 21344 6 io_out[13]
port 77 nsew signal output
rlabel metal3 s 49200 22584 50000 22704 6 io_out[14]
port 78 nsew signal output
rlabel metal3 s 49200 23944 50000 24064 6 io_out[15]
port 79 nsew signal output
rlabel metal3 s 49200 25304 50000 25424 6 io_out[16]
port 80 nsew signal output
rlabel metal3 s 49200 26664 50000 26784 6 io_out[17]
port 81 nsew signal output
rlabel metal3 s 49200 28024 50000 28144 6 io_out[18]
port 82 nsew signal output
rlabel metal3 s 49200 29384 50000 29504 6 io_out[19]
port 83 nsew signal output
rlabel metal3 s 49200 4904 50000 5024 6 io_out[1]
port 84 nsew signal output
rlabel metal3 s 49200 30744 50000 30864 6 io_out[20]
port 85 nsew signal output
rlabel metal3 s 49200 32104 50000 32224 6 io_out[21]
port 86 nsew signal output
rlabel metal3 s 49200 33464 50000 33584 6 io_out[22]
port 87 nsew signal output
rlabel metal3 s 49200 34824 50000 34944 6 io_out[23]
port 88 nsew signal output
rlabel metal3 s 49200 36184 50000 36304 6 io_out[24]
port 89 nsew signal output
rlabel metal3 s 49200 37544 50000 37664 6 io_out[25]
port 90 nsew signal output
rlabel metal3 s 49200 38904 50000 39024 6 io_out[26]
port 91 nsew signal output
rlabel metal3 s 49200 40264 50000 40384 6 io_out[27]
port 92 nsew signal output
rlabel metal3 s 49200 41624 50000 41744 6 io_out[28]
port 93 nsew signal output
rlabel metal3 s 49200 42984 50000 43104 6 io_out[29]
port 94 nsew signal output
rlabel metal3 s 49200 6264 50000 6384 6 io_out[2]
port 95 nsew signal output
rlabel metal3 s 49200 44344 50000 44464 6 io_out[30]
port 96 nsew signal output
rlabel metal3 s 49200 45704 50000 45824 6 io_out[31]
port 97 nsew signal output
rlabel metal3 s 49200 47064 50000 47184 6 io_out[32]
port 98 nsew signal output
rlabel metal3 s 49200 48424 50000 48544 6 io_out[33]
port 99 nsew signal output
rlabel metal3 s 49200 49784 50000 49904 6 io_out[34]
port 100 nsew signal output
rlabel metal3 s 49200 51144 50000 51264 6 io_out[35]
port 101 nsew signal output
rlabel metal3 s 49200 7624 50000 7744 6 io_out[3]
port 102 nsew signal output
rlabel metal3 s 49200 8984 50000 9104 6 io_out[4]
port 103 nsew signal output
rlabel metal3 s 49200 10344 50000 10464 6 io_out[5]
port 104 nsew signal output
rlabel metal3 s 49200 11704 50000 11824 6 io_out[6]
port 105 nsew signal output
rlabel metal3 s 49200 13064 50000 13184 6 io_out[7]
port 106 nsew signal output
rlabel metal3 s 49200 14424 50000 14544 6 io_out[8]
port 107 nsew signal output
rlabel metal3 s 49200 15784 50000 15904 6 io_out[9]
port 108 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 rst_n
port 109 nsew signal input
rlabel metal4 s 4208 2128 4528 52816 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 52816 6 vccd1
port 110 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 52816 6 vssd1
port 111 nsew ground bidirectional
rlabel metal3 s 0 13608 800 13728 6 wb_clk_i
port 112 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 55000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9216114
string GDS_FILE /run/media/tholin/8a6b8802-051e-45a8-8492-771202e4c08a/caravel_user_project/openlane/ScrapCPU/runs/24_05_24_23_48/results/signoff/scrapcpu.magic.gds
string GDS_START 925012
<< end >>

