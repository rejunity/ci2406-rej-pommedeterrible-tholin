// This is the unpowered netlist.
module execution_unit (busy,
    dest_pred_val,
    is_load,
    is_store,
    pred_val,
    rst,
    sign_extend,
    take_branch,
    wb_clk_i,
    curr_PC,
    dest_idx,
    dest_mask,
    dest_pred,
    dest_val,
    instruction,
    loadstore_address,
    loadstore_dest,
    loadstore_size,
    new_PC,
    pred_idx,
    reg1_idx,
    reg1_val,
    reg2_idx,
    reg2_val);
 output busy;
 output dest_pred_val;
 output is_load;
 output is_store;
 input pred_val;
 input rst;
 output sign_extend;
 output take_branch;
 input wb_clk_i;
 input [27:0] curr_PC;
 output [4:0] dest_idx;
 output [1:0] dest_mask;
 output [2:0] dest_pred;
 output [31:0] dest_val;
 input [41:0] instruction;
 output [31:0] loadstore_address;
 output [4:0] loadstore_dest;
 output [1:0] loadstore_size;
 output [27:0] new_PC;
 output [2:0] pred_idx;
 output [4:0] reg1_idx;
 input [31:0] reg1_val;
 output [4:0] reg2_idx;
 input [31:0] reg2_val;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire _06471_;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire busy_l;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire div_complete;
 wire \div_counter[0] ;
 wire \div_counter[1] ;
 wire \div_counter[2] ;
 wire \div_counter[3] ;
 wire \div_counter[4] ;
 wire \div_res[0] ;
 wire \div_res[10] ;
 wire \div_res[11] ;
 wire \div_res[12] ;
 wire \div_res[13] ;
 wire \div_res[14] ;
 wire \div_res[15] ;
 wire \div_res[16] ;
 wire \div_res[17] ;
 wire \div_res[18] ;
 wire \div_res[19] ;
 wire \div_res[1] ;
 wire \div_res[20] ;
 wire \div_res[21] ;
 wire \div_res[22] ;
 wire \div_res[23] ;
 wire \div_res[24] ;
 wire \div_res[25] ;
 wire \div_res[26] ;
 wire \div_res[27] ;
 wire \div_res[28] ;
 wire \div_res[29] ;
 wire \div_res[2] ;
 wire \div_res[30] ;
 wire \div_res[31] ;
 wire \div_res[3] ;
 wire \div_res[4] ;
 wire \div_res[5] ;
 wire \div_res[6] ;
 wire \div_res[7] ;
 wire \div_res[8] ;
 wire \div_res[9] ;
 wire \div_shifter[0] ;
 wire \div_shifter[10] ;
 wire \div_shifter[11] ;
 wire \div_shifter[12] ;
 wire \div_shifter[13] ;
 wire \div_shifter[14] ;
 wire \div_shifter[15] ;
 wire \div_shifter[16] ;
 wire \div_shifter[17] ;
 wire \div_shifter[18] ;
 wire \div_shifter[19] ;
 wire \div_shifter[1] ;
 wire \div_shifter[20] ;
 wire \div_shifter[21] ;
 wire \div_shifter[22] ;
 wire \div_shifter[23] ;
 wire \div_shifter[24] ;
 wire \div_shifter[25] ;
 wire \div_shifter[26] ;
 wire \div_shifter[27] ;
 wire \div_shifter[28] ;
 wire \div_shifter[29] ;
 wire \div_shifter[2] ;
 wire \div_shifter[30] ;
 wire \div_shifter[31] ;
 wire \div_shifter[32] ;
 wire \div_shifter[33] ;
 wire \div_shifter[34] ;
 wire \div_shifter[35] ;
 wire \div_shifter[36] ;
 wire \div_shifter[37] ;
 wire \div_shifter[38] ;
 wire \div_shifter[39] ;
 wire \div_shifter[3] ;
 wire \div_shifter[40] ;
 wire \div_shifter[41] ;
 wire \div_shifter[42] ;
 wire \div_shifter[43] ;
 wire \div_shifter[44] ;
 wire \div_shifter[45] ;
 wire \div_shifter[46] ;
 wire \div_shifter[47] ;
 wire \div_shifter[48] ;
 wire \div_shifter[49] ;
 wire \div_shifter[4] ;
 wire \div_shifter[50] ;
 wire \div_shifter[51] ;
 wire \div_shifter[52] ;
 wire \div_shifter[53] ;
 wire \div_shifter[54] ;
 wire \div_shifter[55] ;
 wire \div_shifter[56] ;
 wire \div_shifter[57] ;
 wire \div_shifter[58] ;
 wire \div_shifter[59] ;
 wire \div_shifter[5] ;
 wire \div_shifter[60] ;
 wire \div_shifter[61] ;
 wire \div_shifter[62] ;
 wire \div_shifter[63] ;
 wire \div_shifter[6] ;
 wire \div_shifter[7] ;
 wire \div_shifter[8] ;
 wire \div_shifter[9] ;
 wire divi1_sign;
 wire \divi2_l[0] ;
 wire \divi2_l[10] ;
 wire \divi2_l[11] ;
 wire \divi2_l[12] ;
 wire \divi2_l[13] ;
 wire \divi2_l[14] ;
 wire \divi2_l[15] ;
 wire \divi2_l[16] ;
 wire \divi2_l[17] ;
 wire \divi2_l[18] ;
 wire \divi2_l[19] ;
 wire \divi2_l[1] ;
 wire \divi2_l[20] ;
 wire \divi2_l[21] ;
 wire \divi2_l[22] ;
 wire \divi2_l[23] ;
 wire \divi2_l[24] ;
 wire \divi2_l[25] ;
 wire \divi2_l[26] ;
 wire \divi2_l[27] ;
 wire \divi2_l[28] ;
 wire \divi2_l[29] ;
 wire \divi2_l[2] ;
 wire \divi2_l[30] ;
 wire \divi2_l[31] ;
 wire \divi2_l[3] ;
 wire \divi2_l[4] ;
 wire \divi2_l[5] ;
 wire \divi2_l[6] ;
 wire \divi2_l[7] ;
 wire \divi2_l[8] ;
 wire \divi2_l[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(curr_PC[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(curr_PC[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(curr_PC[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(instruction[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(instruction[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(instruction[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(instruction[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(instruction[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(instruction[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(reg1_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(reg1_val[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(curr_PC[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(reg1_val[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(reg1_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(reg1_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(reg1_val[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(reg1_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(reg1_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(reg1_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(reg1_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(reg1_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(reg1_val[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(curr_PC[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(reg1_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(reg1_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(reg2_val[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(reg2_val[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(reg2_val[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(reg2_val[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(reg2_val[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(reg2_val[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(reg2_val[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(reg2_val[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(reg2_val[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(reg2_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(reg2_val[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(reg2_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(reg2_val[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(reg2_val[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(reg2_val[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(reg2_val[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(reg2_val[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(reg2_val[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(curr_PC[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(reg2_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(reg2_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(reg2_val[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(reg2_val[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(reg2_val[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(reg2_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(reg2_val[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(reg2_val[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(reg2_val[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(curr_PC[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(pred_val));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(reg1_val[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(reg1_val[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(instruction[41]));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(instruction[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(curr_PC[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(curr_PC[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(curr_PC[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(curr_PC[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA__06509__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__06511__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__06519__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__06522__C_N (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06526__B_N (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06527__B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06529__A3 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06531__B_N (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06532__B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06533__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06534__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06535__A2 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06538__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06541__A1 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06542__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06548__B (.DIODE(_04807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06554__B (.DIODE(_04872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06562__B (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06567__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06568__B (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06570__B (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06571__B (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06574__B (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__B (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06588__B (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06590__A (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06591__B (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06592__B (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06598__B (.DIODE(_05350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06601__B (.DIODE(_05371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06606__B (.DIODE(_05436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06608__B (.DIODE(_05458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06609__B (.DIODE(_05458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06610__B (.DIODE(_05458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06612__A3 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06613__B (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06617__B (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06618__B (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06621__B (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06630__B (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06632__A (.DIODE(_05696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06634__B (.DIODE(_05696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06635__B (.DIODE(_05696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06638__B (.DIODE(_05750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06642__B (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06643__B (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06645__A3 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06646__B (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06654__A3 (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06655__B (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06658__A (.DIODE(_05911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06659__A (.DIODE(_04460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06659__B (.DIODE(_05911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06660__A (.DIODE(_04460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06661__B (.DIODE(_05911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06665__A2 (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__B (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06671__A3 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__A_N (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06673__B (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06674__B (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__A3 (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__A_N (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__B (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__B (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__B (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06683__A3 (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06684__A_N (.DIODE(_06127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06685__B (.DIODE(_06127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06686__B (.DIODE(_06127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__A3 (.DIODE(_04872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06690__A_N (.DIODE(_06181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06691__B (.DIODE(_06181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06692__B (.DIODE(_06181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06695__A3 (.DIODE(_04807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06696__A_N (.DIODE(_06233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06697__B (.DIODE(_06233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06698__B (.DIODE(_06233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06701__A3 (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__A3 (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06703__B (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06704__B (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06705__B (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06708__A3 (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06709__A_N (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06710__B (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06711__B (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__A3 (.DIODE(_05350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06715__A_N (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06716__B (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06718__B (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06721__A3 (.DIODE(_05436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06722__A_N (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06723__B (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06724__B (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06726__C1 (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06727__C_N (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06728__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06729__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__A3 (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06737__A3 (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06738__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__06740__B (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__06743__A3 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06744__A_N (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__B (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06746__B (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06749__A3 (.DIODE(_05750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06750__A_N (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__06751__B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__C1 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06757__B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06759__A3 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__A3 (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__C1 (.DIODE(_05893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06766__B1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__06766__B2 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__B (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__C1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__06828__A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__06828__B (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06847__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06848__A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06849__B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06850__B (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__A2 (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__B1 (.DIODE(_06390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06854__B1 (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06855__B1 (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06856__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__B (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__06859__A_N (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA__06860__B (.DIODE(_06400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06861__B (.DIODE(_06400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06862__B (.DIODE(_06400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06869__B (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06870__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06871__B (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06872__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06873__B (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06874__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06875__B (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06876__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06877__B (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06878__C1 (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__B (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06881__B (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06883__B (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__B (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06887__B (.DIODE(_06392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__A2 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__A2 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__06899__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__A1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__06901__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__06906__B1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__06908__B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__06909__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__B (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__06916__B1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__B1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__B (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__B (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06923__A1 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06924__A1 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__B (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__B (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__D (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__B (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__D (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__06930__A (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06931__A (.DIODE(_06233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06931__B (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06932__A (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__A1 (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__A2 (.DIODE(_06127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__A3 (.DIODE(_06181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__B (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__C (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__B1 (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__A (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06937__A (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06937__B (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__A (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__B (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__B (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__C (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__D (.DIODE(_06127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__A (.DIODE(_06181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__B (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__B2 (.DIODE(_05911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__A1_N (.DIODE(_05911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__B1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__A2 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__A3 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__C (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06955__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__06955__B (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__B (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__C (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__A1 (.DIODE(_06181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06959__A1 (.DIODE(_06127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06959__A2 (.DIODE(_06181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__A (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__B (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__A (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__A (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__B1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__06969__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__06972__B1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__06975__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__06976__S (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06977__A (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__06978__B (.DIODE(_05911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__A (.DIODE(_05696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__B (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__A (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__06995__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__06996__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__S (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__A1 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07005__B1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__B1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__07009__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07010__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07011__S (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__A (.DIODE(_05458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__A1 (.DIODE(_05458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__07027__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07028__B (.DIODE(_05458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__C (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__A1 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__B1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__07040__S (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__A1 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07050__A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__S (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07057__A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__A1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__B2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07061__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07062__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__07063__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__B1 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07069__A (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07069__B (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__A (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__B (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__B (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__C (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__A1 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__A (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__B (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07075__A (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07075__B (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__A1 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__A2 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__B1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__B1 (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07078__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__B (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__A2 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__B1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__C1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__A3 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__B1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__C1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07098__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__A2 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07103__B (.DIODE(_00246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07104__A_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07104__B (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07105__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07105__C_N (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07107__B1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__B (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__C (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07113__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__07113__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__07113__B1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07113__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07115__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__07115__A2 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__A2 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__A1 (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__A3 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__A (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__C (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07133__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__S (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__A (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07140__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A1 (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__C (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__B (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07151__B1 (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__B (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07153__S (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__S (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__A (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__A1 (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__A2 (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__B1 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__B2 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07168__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07168__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07168__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07168__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__A2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07172__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__A2 (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__B1_N (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A2 (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__B1_N (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__B (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__C (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__07187__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07187__B (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__B1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__B2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07189__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07192__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__B1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__A1 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07208__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__B1 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07221__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__B2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07229__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__A1 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__A2 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__B1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__A3 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__B1 (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA__07233__A (.DIODE(_04460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__A_N (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__B (.DIODE(_00386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__C (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__B (.DIODE(_00386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__C_N (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__B (.DIODE(_00386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07253__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__A2 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07255__A (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__B2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__B (.DIODE(_00418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__B (.DIODE(_00418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__B (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__B2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__A (.DIODE(_06127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__A (.DIODE(_06127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__A2 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__B (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__B (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07287__S (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A1 (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__A1_N (.DIODE(_06245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__B2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07293__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__A (.DIODE(_06233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__A2 (.DIODE(_06433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__B (.DIODE(_00451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__B (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__C (.DIODE(_00451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__B (.DIODE(_00451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__A (.DIODE(_06181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__B2 (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__A1 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__B1 (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__B2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__A (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__A1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__B2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A1 (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A2 (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__B1 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__B2 (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07324__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__A1 (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07348__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__A (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07355__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07355__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07355__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07355__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07356__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__A2 (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__B1 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__B2 (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07371__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07373__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__B2 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07385__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07387__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07387__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07387__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07387__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07388__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__B (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__A1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__B1 (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07419__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07422__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07426__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__A2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__B2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__B2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__A2 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__B2 (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07450__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07450__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07450__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07450__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07451__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07452__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__07452__A2 (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07452__B1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07452__B2 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__07453__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__A1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07462__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07464__A (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__A2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__B2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07486__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07492__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__B1 (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07493__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__07494__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__B1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07512__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__B (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__A1 (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__B2 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07525__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__A1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07527__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A2 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__B2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07556__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07556__A2 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07556__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07556__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__A2 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__B1 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__B2 (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__A1 (.DIODE(_04504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__A1 (.DIODE(_04504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__S (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__B2 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A2 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__B2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__A (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__A2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__A2 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__A1 (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__A3 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__B1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__A1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__B2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__A1 (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07628__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07628__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07628__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07628__B2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__A1 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__B2 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07677__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__B1 (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__A2 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__B2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__A1 (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07687__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__B1 (.DIODE(_00137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__A (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__A1 (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__B2 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07706__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07706__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07706__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07706__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A2 (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07716__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__A2 (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__B1 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07721__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__B1 (.DIODE(_00152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__B (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__B1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__B2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07770__A (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07776__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__A2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__A (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__B (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__A2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__B2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__B1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__07842__A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__A2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__B2 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__07844__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__A2 (.DIODE(_00193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__B1 (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__07847__A (.DIODE(_00179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__B2 (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__07866__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__B2 (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__B2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__A1 (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__A2 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__B1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__07907__B1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__A1 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__07923__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07923__A2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__07923__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07923__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07924__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__07937__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__07939__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__B2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__07951__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__B (.DIODE(_01100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__B1 (.DIODE(_01100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__B (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__07995__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08003__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08008__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__A2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08068__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08081__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08081__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08081__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08081__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__B2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08108__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__A2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__B2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__B2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__B (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__B2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__A (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__A1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__B2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__B2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08179__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__A2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__B1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__B2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__B (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__A1 (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__A2 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__B1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__B1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__B2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__B (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08235__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__B2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A1 (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A2 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__B (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__B1 (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__A (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08285__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__08285__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__08285__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08285__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__B1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08296__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08297__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08297__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08297__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__08297__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08300__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08300__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08300__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08300__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08301__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08333__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08333__B (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__A_N (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__B2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08346__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__A2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__B1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08380__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08383__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__A (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__A1 (.DIODE(_06456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__A2 (.DIODE(_06457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__B1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__08386__A1 (.DIODE(_01537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08386__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__B (.DIODE(_01537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__A2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08390__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08396__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08428__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08430__B (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08434__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08436__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08438__B2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08444__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08446__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08480__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08480__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08480__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08480__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08484__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__B1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__B2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08486__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08488__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08492__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08494__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08523__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__B2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08531__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08535__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08541__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08543__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08565__B (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__B2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08567__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08568__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__A2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__B2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08571__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08573__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08594__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08596__B2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08600__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08606__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08606__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08606__B1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08606__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08608__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08610__B2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08631__B2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08635__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__B (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08645__A1 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08659__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__A2 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__B1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__B2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08661__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__A1 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08663__B2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__A2 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__B1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08672__B2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08687__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08687__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08687__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08687__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08688__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__B1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__B2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08690__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08692__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__A1 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08698__A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__A2 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__08699__B1 (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08700__A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__08700__B (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08701__A2 (.DIODE(_01853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08713__A (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08714__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__A1 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__A2 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08715__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08716__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__A2 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08718__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08730__C (.DIODE(_01853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__08733__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__A2 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__B2 (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA__08736__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08738__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__A2 (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__B1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08755__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08755__B (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__A2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08756__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08758__A1 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__08766__B1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A1 (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A2 (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__B1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__08768__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__08768__B (.DIODE(_01918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08768__C (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__A1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08770__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__A_N (.DIODE(_01924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08780__A (.DIODE(_01924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08782__A1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__08782__A2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__08782__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__08782__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08784__A (.DIODE(_01924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08786__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__A1 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__B1 (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__B2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__08788__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08788__B (.DIODE(_01940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08791__A1 (.DIODE(_01924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08798__B (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__08801__A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__B2 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08806__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__A1 (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__A2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__B1 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__B2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08808__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08813__A1 (.DIODE(net252));
 sky130_fd_sc_hd__diode_2 ANTENNA__08813__A2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08813__B1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08813__B2 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__08814__A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__B (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__08816__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08822__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__08824__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A1 (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A1 (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__B (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08856__B (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08858__B (.DIODE(_02008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08874__A2 (.DIODE(_02024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__A2 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08878__A2 (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__A2 (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08882__A2 (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__08886__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08888__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__08888__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__08888__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__08888__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__08889__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__A2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__08905__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__B2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__A1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__B1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__B2 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__08910__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__08915__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__08915__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08915__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__08915__B2 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__08916__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__08917__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08917__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__08917__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08917__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__B2 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__08922__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__A2 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__A3 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08928__B2 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__A1 (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__A2 (.DIODE(_00756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08930__B1 (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08936__A (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08936__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__B2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__B1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08950__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__A2 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__08954__B2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__08982__A (.DIODE(_02035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__B (.DIODE(_02031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__B (.DIODE(_02027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__A_N (.DIODE(_02024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__A1 (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__A (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09036__A1 (.DIODE(_01993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__A (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__D (.DIODE(_02211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09060__B (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09061__B (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09062__B1 (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__A1 (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__B1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09065__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09066__A0 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__S (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09083__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__A0 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09087__S (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__S (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09105__A0 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09109__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__A0 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__S (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__09135__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09143__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__09143__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__09145__B (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__B (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09149__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__09149__A2 (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__B (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__B (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__A (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09153__A (.DIODE(_06395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09156__B (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__S (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__A1 (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__09173__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__A1 (.DIODE(_02326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__S (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09179__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__A2 (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__B2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__09181__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__B1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__09185__B2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09201__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09203__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09204__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__09206__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09212__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09213__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09214__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09218__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__09222__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__09223__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__B (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09224__C (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__A1 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__A2 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__B1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09226__B1 (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09228__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__B1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__B1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09250__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__B2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__09284__A1 (.DIODE(_02035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A1 (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__A1 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__B1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09288__A1 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__09294__S (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__S (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__09296__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__S (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__S (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09304__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09308__S (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__S (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__S (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA__09321__S (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09322__S (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__B1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__09330__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__09330__B (.DIODE(_02481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__A3 (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__09336__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09336__C (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09338__A2 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A2 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__A2 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__B (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__B1 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09345__B2 (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__A2 (.DIODE(_02481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09347__A2 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__B2 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09350__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__09353__B1 (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09357__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__09359__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__A2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__B1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__B2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09397__B2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09400__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__09400__A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09400__B1 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09400__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09403__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09409__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__B2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__09419__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09420__A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__B2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__09430__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09462__A1 (.DIODE(_02035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__A (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__C_N (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__A1 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09467__A1 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__09475__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09476__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__S (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__09482__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09486__S (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__A (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__B (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09504__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__A3 (.DIODE(_02300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09510__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__B1 (.DIODE(_06390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__B1 (.DIODE(_02663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__B2 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__A2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__A_N (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__B (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__C (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__A1 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__A2 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__B1 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__B2 (.DIODE(_00209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__09564__A (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09568__A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__09568__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09570__B2 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09580__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A2 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09582__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09586__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__A_N (.DIODE(_02135_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__B (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__C (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09619__B1 (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__A2 (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09620__C1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09622__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09624__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09626__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09630__S (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__09634__A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__B1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09650__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09660__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09662__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__A2 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__B1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09664__B (.DIODE(_02811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09666__A1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__09670__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__A2 (.DIODE(_02817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__09676__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__A1_N (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__A2_N (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__B1 (.DIODE(_00430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09678__B2 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09682__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__A1 (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09700__B2 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__B2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09706__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A2 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A3 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__B1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09708__A (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09716__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09718__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09722__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__B1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__B2 (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA__09726__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__09728__A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09740__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09742__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__A (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__A1 (.DIODE(_02035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__A1 (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__A1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__A1 (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__B1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09796__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__A1 (.DIODE(_06281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__A2 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__B1 (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09812__A2 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09812__B1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09816__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__B (.DIODE(_02937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__B1 (.DIODE(_02967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__B2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__09832__A1_N (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__09832__A2_N (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__09832__B1 (.DIODE(_00430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09832__B2 (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__09846__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09846__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09846__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09846__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__A1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__B2 (.DIODE(_00168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__A2 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__09861__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__B (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09863__A_N (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__09867__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__A2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__09873__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__B2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__09881__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__09883__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__09885__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__A (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__C (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__B1 (.DIODE(_03064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__B (.DIODE(_03064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09921__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__09948__B1 (.DIODE(_02300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__B1 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__A1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__A2 (.DIODE(_03103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__B1 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__09964__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__B2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__09966__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__B1 (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__B2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__B2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__09979__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09980__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__B1 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__C1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__A1 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__A2 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__A3 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__B1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09996__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__A2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__B1 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__B2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__10002__A (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__A2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10010__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__B1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__B2 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__A1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__B2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10020__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__A (.DIODE(_03064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10054__B1 (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__A2 (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__C1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10056__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__B1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__10076__S (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__A1_N (.DIODE(_06265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10083__A2_N (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__10084__A2 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10084__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__10085__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10089__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__C (.DIODE(_03209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__D (.DIODE(_03237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__B2 (.DIODE(_03238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10099__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__10099__A2 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__10099__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10099__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10100__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__B2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__A2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__B2 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__10113__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10120__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__10120__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10120__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__10120__B2 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__10121__A (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__B (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__C (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__A1 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__A2 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__10124__B1 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10125__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__B1 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__A3 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__B2 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__A1 (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__A2 (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__B1 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__B2 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10137__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__A2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__B2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__B2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__A2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__A1 (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__A1 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10185__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__A1 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10191__B1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__B1 (.DIODE(_06258_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__B2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__A2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__A2 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__B1 (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__A1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__B1 (.DIODE(_03366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__A2 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__A3 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__B1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__A2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__B1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__B2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__A1 (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__A2 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__B2 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__10238__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__A1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__B2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10241__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__B (.DIODE(_00756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10252__A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__A2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__B1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__B2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10264__A1 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10264__A2 (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10264__B1 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10264__B2 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__A (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10317__A1 (.DIODE(_02035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10317__B1_N (.DIODE(_03460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10320__B (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__A (.DIODE(_02766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__C (.DIODE(_03064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10322__A1 (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10322__A2 (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10322__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10323__A1 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10323__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__A1 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__10332__C1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__S (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__10344__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__A1_N (.DIODE(_06252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__A2_N (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__A2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__B2 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__A3 (.DIODE(_03477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__A4 (.DIODE(_03497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A1_N (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A2_N (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__B2 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__A (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__B (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__A2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__B1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__B2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__B2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__10391__B2 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__10392__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10393__B (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10393__C (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10394__A1 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10394__A2 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10394__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__10395__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__10396__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__10397__B1 (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__A (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10411__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__B1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10413__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__A (.DIODE(_03199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__B (.DIODE(_03329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__D_N (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10448__B1 (.DIODE(_03590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__B (.DIODE(_03590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10450__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__B1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__B1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__S (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__10464__S (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__A1 (.DIODE(_06246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__A2 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__C1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__B1 (.DIODE(_03614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__B2 (.DIODE(_03615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__A1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__A3 (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__B2 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__B2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__A2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__B2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10498__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__B1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10503__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__10515__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10515__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10515__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10515__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__A2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__A1 (.DIODE(_03590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A1 (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__B1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__A1 (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__C1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A0 (.DIODE(_02300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A1 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10587__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A1_N (.DIODE(_06233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__A2_N (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__C1 (.DIODE(_03734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__B1 (.DIODE(_03738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10599__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__A2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__B2 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__10609__A (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10623__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10623__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10623__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10623__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10625__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__10625__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10625__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10625__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__A2 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__B1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10635__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10641__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__A (.DIODE(_03590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__B (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__A (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10685__A1 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10685__B1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__C1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10702__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10702__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__A0 (.DIODE(_02300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__A1 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__10710__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__A1 (.DIODE(_06181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__B1 (.DIODE(_03852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__C1 (.DIODE(_03853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10714__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__C1 (.DIODE(_03857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10719__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__10720__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__B2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10725__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__A1 (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__A2 (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__B2 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10729__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10731__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10735__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__10739__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10739__A2 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10739__B1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10739__B2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10740__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10741__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10741__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10741__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10741__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10745__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10745__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10745__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10745__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__B1 (.DIODE(_00430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__C1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10751__A1 (.DIODE(_00430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10751__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__A2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__B1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10759__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10760__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__B (.DIODE(_00756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__A2 (.DIODE(_00756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__B2 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10796__B (.DIODE(_03936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__A1 (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__A (.DIODE(_04504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10804__B1 (.DIODE(_04504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10806__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__C1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__10825__A1 (.DIODE(_06127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10825__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__10826__B (.DIODE(_03963_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__10830__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__B1 (.DIODE(_03971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10833__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10834__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10835__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10835__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10835__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10835__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10836__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10838__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__10842__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10845__A (.DIODE(_00219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10845__B (.DIODE(_00221_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__A1 (.DIODE(_00225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__A2 (.DIODE(_00226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10846__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10847__C_N (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__B1_N (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__B1 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10850__A (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__10852__B2 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__10853__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__10858__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10858__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10858__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10858__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__10865__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10865__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10865__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10865__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10866__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__B2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10875__A_N (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10875__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__10876__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__10876__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__A2 (.DIODE(_03936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10908__B (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10910__B1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10914__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__10916__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__C1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__S (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__S (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__C1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__10933__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__C1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__A1 (.DIODE(_06082_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__B1 (.DIODE(_04075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__C1 (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__B1 (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__B1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__B2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__10954__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__10963__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__10965__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__10970__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__10973__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__A1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__10975__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__B1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__A2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__B1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__10982__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__A1 (.DIODE(_03936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11023__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__11025__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__11027__C1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__S (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__C1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11042__C1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__C1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__A1 (.DIODE(_06046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__11048__D1 (.DIODE(_04178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11049__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__11049__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__A3 (.DIODE(_04166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__A4 (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11054__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11056__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11060__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11067__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11067__A2 (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__11067__B1 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__11067__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__A_N (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__11070__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__A1 (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__A2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__B2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__11072__A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__11077__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__11077__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11077__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11077__B2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__11079__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11079__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11079__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11079__B2 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__11080__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11082__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__A (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11091__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11120__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__11124__A (.DIODE(_04504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11126__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__B1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11136__S (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__C1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__A0 (.DIODE(_02300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__A1 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__A1 (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__A2 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__C1 (.DIODE(_04284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__A1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__B1 (.DIODE(_04287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__11157__B (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11161__B1 (.DIODE(_04293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__A1 (.DIODE(_03460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__B1 (.DIODE(_04297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11163__A (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11163__D_N (.DIODE(_02035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__A (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__B (.DIODE(_04300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__B (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__A2 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11173__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__B2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__B (.DIODE(_00386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__C (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__A2_N (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__B2 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11198__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__A1 (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__A2 (.DIODE(_04300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__A (.DIODE(_03822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__B (.DIODE(_04371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__A (.DIODE(_02137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__A1 (.DIODE(_04504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11254__C1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__A2 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__B1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__A1 (.DIODE(_05911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__B1 (.DIODE(_02300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__C1 (.DIODE(_04400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__B2 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11267__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11269__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__A1 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__A2 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__B1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__B2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11273__A (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11281__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11281__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11281__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11281__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11282__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__B2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__A2 (.DIODE(_04371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11333__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__11336__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__B1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11347__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__A2 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11351__B1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__B1 (.DIODE(_02300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__C1 (.DIODE(_06390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11353__C1 (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11356__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11358__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11363__B2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11364__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__11366__A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11368__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11374__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__A2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__B1 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11376__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11380__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__B (.DIODE(_00756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__A2 (.DIODE(_00756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11386__B2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__B (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__A1 (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__A2 (.DIODE(_04300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__A2 (.DIODE(_04371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__B1 (.DIODE(_02137_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__B1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11432__C1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11439__A0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__11439__A1 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__A2_N (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__B1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11441__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11450__B (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11452__B2 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11453__A1 (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11453__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__11456__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__B2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11462__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11463__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__11463__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11466__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__A (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11469__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11469__A2 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA__11469__B1 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__11469__B2 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__B1 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__A2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__A (.DIODE(_04371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11514__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11515__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__B1 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11520__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__11522__C1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11534__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11535__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__C1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A1 (.DIODE(_05696_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__B1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11548__A1 (.DIODE(_04299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11548__A2 (.DIODE(_04300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__A1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__B2 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__A2 (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__B1 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__B2 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__A1 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__A2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__B1 (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11558__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__A2 (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__B2 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__B2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__A (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__A1 (.DIODE(_00436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__A1 (.DIODE(_04371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11605__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__B1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__B (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__11626__A2 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11626__C1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11627__A2 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11628__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11628__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__11629__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__11632__A1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__S (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__B2 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__B2 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__11640__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__B2 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11642__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11649__A (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11649__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__A1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__A2 (.DIODE(_00307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__B1 (.DIODE(_00308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__B2 (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11652__A (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__A_N (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11654__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__A1 (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11656__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__11663__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__A1 (.DIODE(_04371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__11686__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11690__C1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11697__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11697__C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__11700__C1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__A0 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__A1 (.DIODE(_05544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__11713__A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11714__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__11715__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11715__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11715__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11715__B2 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11717__B2 (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__A1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__A2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__B1 (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11727__B (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A2 (.DIODE(_00756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__A1 (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__A1 (.DIODE(_04371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__B1 (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__C1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__11774__A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11775__A1 (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__11775__C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__11778__C1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__A0 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__11783__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11787__C1 (.DIODE(_04974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__A1 (.DIODE(_05458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__A2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__B1 (.DIODE(_06390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__B1 (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__B2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__11794__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__11795__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__B2 (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__11799__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__A1 (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__B2 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__11809__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__B1 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__A_N (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__A2 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__A1 (.DIODE(_04371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__B1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__S (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__11853__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11858__A0 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11858__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__B1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__11862__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__B2 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__C1 (.DIODE(_05056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11864__A1 (.DIODE(_05371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11864__A2 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__11868__A1 (.DIODE(_06390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11874__A2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11874__B1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__A3 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__11876__A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA__11876__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__A1 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__B1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__A1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__B2 (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11885__A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__A2 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__B1 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11887__A (.DIODE(_00248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11910__A (.DIODE(_04371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11919__B1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11925__A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11926__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11926__C1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__11936__A2 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11936__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__11937__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__B1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__11943__A1 (.DIODE(_06390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11945__A1 (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA__11945__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__11945__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__11945__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__11946__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11950__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__11950__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__11954__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__11956__A (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__B1 (.DIODE(_00757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__B2 (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__B1 (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__A1 (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__B1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__B1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__B1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__C1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__12003__C1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A2 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__12007__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__12010__B2 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12012__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__12013__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__A2 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__B1 (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__12017__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12017__A3 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12017__B1 (.DIODE(_00248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__A2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__B2 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__B (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__B1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__S (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__B1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12070__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12070__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__A2_N (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__B1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12080__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__12081__B1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__A2 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12084__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12085__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__A2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__B1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__B2 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__12096__A0 (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12110__A (.DIODE(_04371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12119__B1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12127__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12128__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__A2 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__B1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__A2 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__B1 (.DIODE(_02300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12133__C1 (.DIODE(_06390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__A1 (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12138__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12139__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__A1_N (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12142__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__A2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12144__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__12148__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12148__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__A1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__A2 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12176__C1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__12182__A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__12183__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__12183__C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12186__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__A2 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__B1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12192__A2 (.DIODE(_02300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12192__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__12193__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__A1 (.DIODE(_05263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__A2 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__C1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__12198__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__12198__A2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__12198__B1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12198__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__A1 (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__A2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__12200__B1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__C_N (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__12222__C1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__12224__A1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__12228__B1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__12229__C1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__12231__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12237__A2 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12237__B1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12238__A2 (.DIODE(_02300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12238__C1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__B (.DIODE(_05459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12241__A1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__A2 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__C1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__B (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__C (.DIODE(_00757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__A2 (.DIODE(_00757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__12247__A0 (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__A_N (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__B (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__B1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__C1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__12266__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__A (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12271__S (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__A2 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__A0 (.DIODE(_02295_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__A1 (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__A1 (.DIODE(_02291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__A1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__12284__A1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__A1 (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__A2 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__C1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__A2 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__12294__C1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__12298__A1 (.DIODE(_02138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12298__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A (.DIODE(_02211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__A1 (.DIODE(_02211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__B1 (.DIODE(_02298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__12304__B1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__A2 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__B1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__12310__A2 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12310__A3 (.DIODE(_02300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12310__C1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__A2 (.DIODE(_02294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__A1 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__B1 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__A1 (.DIODE(_02293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__A1 (.DIODE(_04752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__A2 (.DIODE(_06426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__C1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__A0 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__A (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__A (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12322__A (.DIODE(_05893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__A (.DIODE(_05893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__A (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12330__A (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12336__A (.DIODE(_05750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__A (.DIODE(_05750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12344__A (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12350__A (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__A (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__A (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12358__A (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__A (.DIODE(_05436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12365__A (.DIODE(_05436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12371__A (.DIODE(_05350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__A (.DIODE(_05350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__A (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12379__A (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12385__A (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__A (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__A (.DIODE(_04807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12393__A (.DIODE(_04807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12399__A (.DIODE(_04872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__A (.DIODE(_04872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12405__A0 (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__A (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12407__A (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12413__A (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12414__A (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__A (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12421__A (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__C (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__12499__B (.DIODE(_04654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__B (.DIODE(_05893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12506__B (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__B (.DIODE(_05823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__B (.DIODE(_05750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12512__B (.DIODE(_05750_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12516__B (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12517__B (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__B (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12522__B (.DIODE(_05591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12526__B (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12527__B (.DIODE(_05512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__B (.DIODE(_05436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12532__B (.DIODE(_05436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__B (.DIODE(_05350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__B (.DIODE(_05350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__B (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12542__B (.DIODE(_05089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__B (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12546__B (.DIODE(_04959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12552__B (.DIODE(_04807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__B (.DIODE(_04807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12558__B (.DIODE(_04872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__B (.DIODE(_04872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12564__B (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__B (.DIODE(_05241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12570__B (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12571__B (.DIODE(_05165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12576__B (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__A2 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12663__B (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12667__A1 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12667__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12669__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12675__C1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__12676__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12677__A1 (.DIODE(_00263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12677__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12677__C1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__12678__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__A1 (.DIODE(_00300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12680__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12681__A1 (.DIODE(_00310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12681__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12683__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12684__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__12686__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__12688__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__12688__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12690__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__12690__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12692__B (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__A1 (.DIODE(_00430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12694__A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__12694__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12695__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12696__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__A1 (.DIODE(_06483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12698__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__A1 (.DIODE(_06459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12700__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__A1 (.DIODE(_06467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__C1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__12702__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__12702__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12703__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12704__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__12706__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__12708__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12709__A1 (.DIODE(_06503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12709__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12710__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__12716__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__A1 (.DIODE(_00197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12723__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12725__A1 (.DIODE(_00222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12725__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12727__A1 (.DIODE(_00228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12727__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__A (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__A2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12729__C1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__B (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__A1 (.DIODE(_00756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__A2 (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA__12731__C1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__12835__B1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__12836__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__12837__A2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__12838__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__12840__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12842__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12844__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12846__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12848__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12850__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12852__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12854__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12856__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12858__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12874__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12880__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12882__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12886__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__12892__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__12894__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__12896__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__12898__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12899__B2 (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__A1 (.DIODE(_00187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12902__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__A1 (.DIODE(_00180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12906__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12910__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__12914__A1 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__12914__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12918__A1 (.DIODE(_06490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12918__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12922__A1 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__12924__A1 (.DIODE(_06440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12926__A1 (.DIODE(_06435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12926__A2 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__12928__A1 (.DIODE(_06474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12928__A2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__12930__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__12932__A1 (.DIODE(_00386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12934__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__12936__A1 (.DIODE(_00451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12938__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__12940__A1 (.DIODE(_00437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12942__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__12944__A1 (.DIODE(_00284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12946__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__12948__A1 (.DIODE(_00301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12950__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__12954__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__12956__A1 (.DIODE(_00333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__12957__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12958__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__12959__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12960__A1 (.DIODE(_00418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12961__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__12962__B1 (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12963__C (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__12964__A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__A1 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__12965__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12968__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12969__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__12973__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12974__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__12975__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__12978__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__12979__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__12979__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__12980__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__12982__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__12983__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__12984__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__12986__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__12987__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__12987__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12992__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__12997__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__13001__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13002__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13006__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13007__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13007__B2 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__13011__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13012__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13016__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13017__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13022__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13023__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__13026__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13027__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13031__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13032__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13036__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13038__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__13041__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13043__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__13046__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13048__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__13051__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13056__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13060__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13065__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13067__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__13069__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13071__A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__13074__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13078__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13083__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13085__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__13087__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13088__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13088__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13092__S (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13093__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13096__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13097__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13101__S (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13102__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13102__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13105__B (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13106__A2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__13107__A2 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13107__B2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13108__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__13110__A2 (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA__13110__B1 (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA__13111__A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__13113__A2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__13114__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13114__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13116__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13119__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA__13122__A2 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__13122__B2 (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_wb_clk_i_A (.DIODE(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout103_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout106_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout10_A (.DIODE(_00408_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(_00255_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout111_A (.DIODE(_00248_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout112_A (.DIODE(_00248_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(_00248_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout114_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(_00152_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout11_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(_06484_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(_06482_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout126_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(_06460_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout13_A (.DIODE(_00306_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(_00290_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(_00275_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(_00275_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout14_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(_00137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout158_A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(_00209_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(_00194_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(_00193_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(_00168_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(_00164_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout18_A (.DIODE(_00223_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(_06489_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout195_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout19_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout207_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(_00179_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(_06413_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout223_A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout225_A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout226_A (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout22_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout231_A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(_06287_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(_06281_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(_02494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(_02494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout246_A (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(_02494_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(_02299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout252_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout254_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout255_A (.DIODE(_00188_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout258_A (.DIODE(_06391_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout259_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout260_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(_06391_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout262_A (.DIODE(_06390_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout263_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout26_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout273_A (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout28_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout293_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout29_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(_04504_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout30_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout31_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout33_A (.DIODE(_00728_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout34_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout35_A (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout36_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout38_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout3_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout40_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout42_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout44_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout45_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout47_A (.DIODE(_00309_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout48_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout4_A (.DIODE(_00757_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout50_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout52_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout53_A (.DIODE(_00265_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout54_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout55_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout57_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout58_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout5_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout60_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout62_A (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout63_A (.DIODE(_00185_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout64_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout65_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout67_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout68_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout70_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout71_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout73_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout74_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout76_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout77_A (.DIODE(_00136_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout78_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout7_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout80_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout82_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout84_A (.DIODE(_02137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout85_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(_02137_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(_00457_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout8_A (.DIODE(_00421_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout94_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(_00391_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout96_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout9_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap256_A (.DIODE(_00187_));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_676 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_170 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_366 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_395 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_539 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_20 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_532 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_622 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_618 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_359 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_104 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_562 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_24 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_738 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_38 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_776 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_280 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_14 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_646 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_420 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _06504_ (.A(net553),
    .Y(_04340_));
 sky130_fd_sc_hd__inv_2 _06505_ (.A(net559),
    .Y(_04351_));
 sky130_fd_sc_hd__inv_2 _06506_ (.A(net367),
    .Y(_04362_));
 sky130_fd_sc_hd__inv_2 _06507_ (.A(net363),
    .Y(_04373_));
 sky130_fd_sc_hd__inv_2 _06508_ (.A(\div_shifter[28] ),
    .Y(_04384_));
 sky130_fd_sc_hd__inv_2 _06509_ (.A(net272),
    .Y(_04395_));
 sky130_fd_sc_hd__inv_2 _06510_ (.A(instruction[3]),
    .Y(_04406_));
 sky130_fd_sc_hd__clkinv_4 _06511_ (.A(net304),
    .Y(_04416_));
 sky130_fd_sc_hd__inv_2 _06512_ (.A(instruction[41]),
    .Y(_04427_));
 sky130_fd_sc_hd__inv_2 _06513_ (.A(reg1_val[1]),
    .Y(_04438_));
 sky130_fd_sc_hd__inv_2 _06514_ (.A(reg1_val[4]),
    .Y(_04449_));
 sky130_fd_sc_hd__inv_2 _06515_ (.A(reg1_val[16]),
    .Y(_04460_));
 sky130_fd_sc_hd__inv_2 _06516_ (.A(reg1_val[22]),
    .Y(_04471_));
 sky130_fd_sc_hd__inv_2 _06517_ (.A(reg1_val[26]),
    .Y(_04482_));
 sky130_fd_sc_hd__inv_2 _06518_ (.A(reg1_val[30]),
    .Y(_04493_));
 sky130_fd_sc_hd__inv_2 _06519_ (.A(net307),
    .Y(_04504_));
 sky130_fd_sc_hd__inv_2 _06520_ (.A(curr_PC[0]),
    .Y(_04514_));
 sky130_fd_sc_hd__inv_2 _06521_ (.A(rst),
    .Y(_04525_));
 sky130_fd_sc_hd__or4bb_4 _06522_ (.A(instruction[0]),
    .B(instruction[1]),
    .C_N(net308),
    .D_N(pred_val),
    .X(_04536_));
 sky130_fd_sc_hd__nor2_8 _06523_ (.A(instruction[3]),
    .B(_04536_),
    .Y(is_load));
 sky130_fd_sc_hd__nor2_8 _06524_ (.A(_04406_),
    .B(_04536_),
    .Y(is_store));
 sky130_fd_sc_hd__and3b_1 _06525_ (.A_N(instruction[0]),
    .B(pred_val),
    .C(instruction[1]),
    .X(_04567_));
 sky130_fd_sc_hd__and4bb_1 _06526_ (.A_N(instruction[0]),
    .B_N(net308),
    .C(instruction[1]),
    .D(pred_val),
    .X(_04578_));
 sky130_fd_sc_hd__or4bb_2 _06527_ (.A(instruction[0]),
    .B(net308),
    .C_N(instruction[1]),
    .D_N(pred_val),
    .X(_04589_));
 sky130_fd_sc_hd__and2_1 _06528_ (.A(reg2_val[31]),
    .B(net284),
    .X(_04600_));
 sky130_fd_sc_hd__o31a_1 _06529_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(net308),
    .B1(pred_val),
    .X(_04611_));
 sky130_fd_sc_hd__o311a_1 _06530_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(instruction[2]),
    .B1(instruction[41]),
    .C1(pred_val),
    .X(_04621_));
 sky130_fd_sc_hd__and4bb_1 _06531_ (.A_N(instruction[1]),
    .B_N(net308),
    .C(instruction[0]),
    .D(pred_val),
    .X(_04632_));
 sky130_fd_sc_hd__or4bb_4 _06532_ (.A(instruction[1]),
    .B(net308),
    .C_N(instruction[0]),
    .D_N(pred_val),
    .X(_04643_));
 sky130_fd_sc_hd__and2_2 _06533_ (.A(instruction[25]),
    .B(net282),
    .X(_04654_));
 sky130_fd_sc_hd__o211a_1 _06534_ (.A1(instruction[1]),
    .A2(net308),
    .B1(instruction[25]),
    .C1(pred_val),
    .X(_04665_));
 sky130_fd_sc_hd__o211ai_4 _06535_ (.A1(instruction[1]),
    .A2(net308),
    .B1(instruction[25]),
    .C1(pred_val),
    .Y(_04676_));
 sky130_fd_sc_hd__a21o_1 _06536_ (.A1(instruction[41]),
    .A2(_04632_),
    .B1(_04665_),
    .X(_04687_));
 sky130_fd_sc_hd__a21oi_2 _06537_ (.A1(instruction[41]),
    .A2(_04632_),
    .B1(_04665_),
    .Y(_04698_));
 sky130_fd_sc_hd__a221o_1 _06538_ (.A1(instruction[24]),
    .A2(net280),
    .B1(_04632_),
    .B2(instruction[41]),
    .C1(_04665_),
    .X(_04709_));
 sky130_fd_sc_hd__and2_2 _06539_ (.A(net287),
    .B(_04709_),
    .X(_04719_));
 sky130_fd_sc_hd__nand2_1 _06540_ (.A(net287),
    .B(_04709_),
    .Y(_04730_));
 sky130_fd_sc_hd__a21oi_4 _06541_ (.A1(net280),
    .A2(net243),
    .B1(_04600_),
    .Y(_04741_));
 sky130_fd_sc_hd__a31o_4 _06542_ (.A1(net287),
    .A2(net280),
    .A3(_04709_),
    .B1(_04600_),
    .X(_04752_));
 sky130_fd_sc_hd__and2_1 _06543_ (.A(reg1_val[31]),
    .B(_04741_),
    .X(_04763_));
 sky130_fd_sc_hd__nor2_1 _06544_ (.A(reg1_val[31]),
    .B(_04741_),
    .Y(_04774_));
 sky130_fd_sc_hd__or2_4 _06545_ (.A(_04763_),
    .B(_04774_),
    .X(_04785_));
 sky130_fd_sc_hd__inv_2 _06546_ (.A(_04785_),
    .Y(_04796_));
 sky130_fd_sc_hd__and2_4 _06547_ (.A(instruction[36]),
    .B(net281),
    .X(_04807_));
 sky130_fd_sc_hd__or2_1 _06548_ (.A(net266),
    .B(_04807_),
    .X(_04817_));
 sky130_fd_sc_hd__a22o_2 _06549_ (.A1(reg2_val[26]),
    .A2(net285),
    .B1(_04719_),
    .B2(_04817_),
    .X(_04828_));
 sky130_fd_sc_hd__nand2_1 _06550_ (.A(reg1_val[26]),
    .B(_04828_),
    .Y(_04839_));
 sky130_fd_sc_hd__or2_1 _06551_ (.A(reg1_val[26]),
    .B(_04828_),
    .X(_04850_));
 sky130_fd_sc_hd__and2_1 _06552_ (.A(_04839_),
    .B(_04850_),
    .X(_04861_));
 sky130_fd_sc_hd__and2_4 _06553_ (.A(instruction[37]),
    .B(net281),
    .X(_04872_));
 sky130_fd_sc_hd__or2_1 _06554_ (.A(net266),
    .B(_04872_),
    .X(_04883_));
 sky130_fd_sc_hd__a22o_2 _06555_ (.A1(reg2_val[27]),
    .A2(net285),
    .B1(net243),
    .B2(_04883_),
    .X(_04894_));
 sky130_fd_sc_hd__inv_2 _06556_ (.A(_04894_),
    .Y(_04904_));
 sky130_fd_sc_hd__and2_1 _06557_ (.A(reg1_val[27]),
    .B(_04894_),
    .X(_04915_));
 sky130_fd_sc_hd__nor2_1 _06558_ (.A(reg1_val[27]),
    .B(_04894_),
    .Y(_04926_));
 sky130_fd_sc_hd__inv_2 _06559_ (.A(_04926_),
    .Y(_04937_));
 sky130_fd_sc_hd__nor2_1 _06560_ (.A(_04915_),
    .B(_04926_),
    .Y(_04948_));
 sky130_fd_sc_hd__and2_4 _06561_ (.A(instruction[35]),
    .B(net281),
    .X(_04959_));
 sky130_fd_sc_hd__nor2_1 _06562_ (.A(net266),
    .B(_04959_),
    .Y(_04970_));
 sky130_fd_sc_hd__o2bb2a_2 _06563_ (.A1_N(reg2_val[25]),
    .A2_N(net285),
    .B1(_04730_),
    .B2(_04970_),
    .X(_04980_));
 sky130_fd_sc_hd__nand2b_1 _06564_ (.A_N(_04980_),
    .B(reg1_val[25]),
    .Y(_04991_));
 sky130_fd_sc_hd__nand2b_1 _06565_ (.A_N(reg1_val[25]),
    .B(_04980_),
    .Y(_05002_));
 sky130_fd_sc_hd__and2_1 _06566_ (.A(_04991_),
    .B(_05002_),
    .X(_05013_));
 sky130_fd_sc_hd__and2_4 _06567_ (.A(instruction[40]),
    .B(net282),
    .X(_05024_));
 sky130_fd_sc_hd__or2_1 _06568_ (.A(net266),
    .B(_05024_),
    .X(_05035_));
 sky130_fd_sc_hd__a22o_4 _06569_ (.A1(reg2_val[30]),
    .A2(net283),
    .B1(net243),
    .B2(_05035_),
    .X(_05046_));
 sky130_fd_sc_hd__and2_1 _06570_ (.A(reg1_val[30]),
    .B(_05046_),
    .X(_05057_));
 sky130_fd_sc_hd__nor2_1 _06571_ (.A(reg1_val[30]),
    .B(_05046_),
    .Y(_05067_));
 sky130_fd_sc_hd__nor2_2 _06572_ (.A(_05057_),
    .B(_05067_),
    .Y(_05078_));
 sky130_fd_sc_hd__and2_4 _06573_ (.A(instruction[34]),
    .B(net281),
    .X(_05089_));
 sky130_fd_sc_hd__or2_1 _06574_ (.A(net266),
    .B(_05089_),
    .X(_05100_));
 sky130_fd_sc_hd__a22oi_4 _06575_ (.A1(reg2_val[24]),
    .A2(net285),
    .B1(net243),
    .B2(_05100_),
    .Y(_05111_));
 sky130_fd_sc_hd__a22o_1 _06576_ (.A1(reg2_val[24]),
    .A2(net285),
    .B1(net243),
    .B2(_05100_),
    .X(_05122_));
 sky130_fd_sc_hd__nand2_1 _06577_ (.A(reg1_val[24]),
    .B(_05122_),
    .Y(_05133_));
 sky130_fd_sc_hd__or2_1 _06578_ (.A(reg1_val[24]),
    .B(_05122_),
    .X(_05144_));
 sky130_fd_sc_hd__and2_1 _06579_ (.A(_05133_),
    .B(_05144_),
    .X(_05154_));
 sky130_fd_sc_hd__and2_4 _06580_ (.A(instruction[39]),
    .B(net281),
    .X(_05165_));
 sky130_fd_sc_hd__or2_1 _06581_ (.A(net265),
    .B(_05165_),
    .X(_05176_));
 sky130_fd_sc_hd__a22oi_4 _06582_ (.A1(reg2_val[29]),
    .A2(net284),
    .B1(net243),
    .B2(_05176_),
    .Y(_05187_));
 sky130_fd_sc_hd__a22o_2 _06583_ (.A1(reg2_val[29]),
    .A2(net283),
    .B1(net243),
    .B2(_05176_),
    .X(_05198_));
 sky130_fd_sc_hd__and2_1 _06584_ (.A(reg1_val[29]),
    .B(_05198_),
    .X(_05209_));
 sky130_fd_sc_hd__or2_1 _06585_ (.A(reg1_val[29]),
    .B(_05198_),
    .X(_05220_));
 sky130_fd_sc_hd__and2b_1 _06586_ (.A_N(_05209_),
    .B(_05220_),
    .X(_05230_));
 sky130_fd_sc_hd__and2_4 _06587_ (.A(instruction[38]),
    .B(net281),
    .X(_05241_));
 sky130_fd_sc_hd__or2_1 _06588_ (.A(net266),
    .B(_05241_),
    .X(_05252_));
 sky130_fd_sc_hd__a22o_4 _06589_ (.A1(reg2_val[28]),
    .A2(net283),
    .B1(_04719_),
    .B2(_05252_),
    .X(_05263_));
 sky130_fd_sc_hd__inv_2 _06590_ (.A(_05263_),
    .Y(_05274_));
 sky130_fd_sc_hd__and2_1 _06591_ (.A(reg1_val[28]),
    .B(_05263_),
    .X(_05285_));
 sky130_fd_sc_hd__or2_1 _06592_ (.A(reg1_val[28]),
    .B(_05263_),
    .X(_05295_));
 sky130_fd_sc_hd__and2b_1 _06593_ (.A_N(_05285_),
    .B(_05295_),
    .X(_05306_));
 sky130_fd_sc_hd__or4_1 _06594_ (.A(_04861_),
    .B(_04948_),
    .C(_05013_),
    .D(_05154_),
    .X(_05317_));
 sky130_fd_sc_hd__or4_1 _06595_ (.A(_04785_),
    .B(_05078_),
    .C(_05230_),
    .D(_05306_),
    .X(_05328_));
 sky130_fd_sc_hd__nor2_1 _06596_ (.A(_05317_),
    .B(_05328_),
    .Y(_05339_));
 sky130_fd_sc_hd__and2_4 _06597_ (.A(instruction[33]),
    .B(net281),
    .X(_05350_));
 sky130_fd_sc_hd__or2_1 _06598_ (.A(net266),
    .B(_05350_),
    .X(_05360_));
 sky130_fd_sc_hd__a22oi_4 _06599_ (.A1(reg2_val[23]),
    .A2(net285),
    .B1(net243),
    .B2(_05360_),
    .Y(_05371_));
 sky130_fd_sc_hd__a22o_2 _06600_ (.A1(reg2_val[23]),
    .A2(net285),
    .B1(net243),
    .B2(_05360_),
    .X(_05382_));
 sky130_fd_sc_hd__nand2_1 _06601_ (.A(reg1_val[23]),
    .B(_05371_),
    .Y(_05393_));
 sky130_fd_sc_hd__and2_1 _06602_ (.A(reg1_val[23]),
    .B(_05382_),
    .X(_05404_));
 sky130_fd_sc_hd__nor2_1 _06603_ (.A(reg1_val[23]),
    .B(_05382_),
    .Y(_05415_));
 sky130_fd_sc_hd__nor2_1 _06604_ (.A(_05404_),
    .B(_05415_),
    .Y(_05425_));
 sky130_fd_sc_hd__and2_4 _06605_ (.A(instruction[32]),
    .B(net281),
    .X(_05436_));
 sky130_fd_sc_hd__or2_1 _06606_ (.A(net266),
    .B(_05436_),
    .X(_05447_));
 sky130_fd_sc_hd__a22o_4 _06607_ (.A1(reg2_val[22]),
    .A2(net285),
    .B1(_04719_),
    .B2(_05447_),
    .X(_05458_));
 sky130_fd_sc_hd__or2_1 _06608_ (.A(_04471_),
    .B(_05458_),
    .X(_05469_));
 sky130_fd_sc_hd__and2_1 _06609_ (.A(reg1_val[22]),
    .B(_05458_),
    .X(_05479_));
 sky130_fd_sc_hd__nor2_1 _06610_ (.A(reg1_val[22]),
    .B(_05458_),
    .Y(_05490_));
 sky130_fd_sc_hd__nor2_1 _06611_ (.A(_05479_),
    .B(_05490_),
    .Y(_05501_));
 sky130_fd_sc_hd__o311a_4 _06612_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(net308),
    .B1(instruction[31]),
    .C1(pred_val),
    .X(_05512_));
 sky130_fd_sc_hd__nor2_1 _06613_ (.A(net266),
    .B(_05512_),
    .Y(_05522_));
 sky130_fd_sc_hd__o2bb2a_1 _06614_ (.A1_N(reg2_val[21]),
    .A2_N(net285),
    .B1(_04730_),
    .B2(_05522_),
    .X(_05533_));
 sky130_fd_sc_hd__a2bb2o_2 _06615_ (.A1_N(_05522_),
    .A2_N(_04730_),
    .B1(net285),
    .B2(reg2_val[21]),
    .X(_05544_));
 sky130_fd_sc_hd__nand2_1 _06616_ (.A(reg1_val[21]),
    .B(_05533_),
    .Y(_05553_));
 sky130_fd_sc_hd__and2_1 _06617_ (.A(reg1_val[21]),
    .B(_05544_),
    .X(_05563_));
 sky130_fd_sc_hd__nor2_1 _06618_ (.A(reg1_val[21]),
    .B(_05544_),
    .Y(_05572_));
 sky130_fd_sc_hd__nor2_1 _06619_ (.A(_05563_),
    .B(_05572_),
    .Y(_05582_));
 sky130_fd_sc_hd__and2_4 _06620_ (.A(instruction[30]),
    .B(net281),
    .X(_05591_));
 sky130_fd_sc_hd__or2_1 _06621_ (.A(net265),
    .B(_05591_),
    .X(_05601_));
 sky130_fd_sc_hd__a22oi_4 _06622_ (.A1(reg2_val[20]),
    .A2(net284),
    .B1(net243),
    .B2(_05601_),
    .Y(_05611_));
 sky130_fd_sc_hd__a22o_2 _06623_ (.A1(reg2_val[20]),
    .A2(net284),
    .B1(net243),
    .B2(_05601_),
    .X(_05620_));
 sky130_fd_sc_hd__nand2_1 _06624_ (.A(reg1_val[20]),
    .B(_05611_),
    .Y(_05630_));
 sky130_fd_sc_hd__nand2_1 _06625_ (.A(reg1_val[20]),
    .B(_05620_),
    .Y(_05639_));
 sky130_fd_sc_hd__inv_2 _06626_ (.A(_05639_),
    .Y(_05649_));
 sky130_fd_sc_hd__nor2_1 _06627_ (.A(reg1_val[20]),
    .B(_05620_),
    .Y(_05658_));
 sky130_fd_sc_hd__nor2_1 _06628_ (.A(_05649_),
    .B(_05658_),
    .Y(_05668_));
 sky130_fd_sc_hd__and2_4 _06629_ (.A(instruction[29]),
    .B(net281),
    .X(_05677_));
 sky130_fd_sc_hd__or2_1 _06630_ (.A(net265),
    .B(_05677_),
    .X(_05686_));
 sky130_fd_sc_hd__a22o_2 _06631_ (.A1(reg2_val[19]),
    .A2(net283),
    .B1(net243),
    .B2(_05686_),
    .X(_05696_));
 sky130_fd_sc_hd__inv_2 _06632_ (.A(_05696_),
    .Y(_05705_));
 sky130_fd_sc_hd__nand2_1 _06633_ (.A(reg1_val[19]),
    .B(_05705_),
    .Y(_05715_));
 sky130_fd_sc_hd__nand2_1 _06634_ (.A(reg1_val[19]),
    .B(_05696_),
    .Y(_05723_));
 sky130_fd_sc_hd__or2_1 _06635_ (.A(reg1_val[19]),
    .B(_05696_),
    .X(_05732_));
 sky130_fd_sc_hd__and2_1 _06636_ (.A(_05723_),
    .B(_05732_),
    .X(_05741_));
 sky130_fd_sc_hd__and2_4 _06637_ (.A(instruction[28]),
    .B(net281),
    .X(_05750_));
 sky130_fd_sc_hd__or2_1 _06638_ (.A(net265),
    .B(_05750_),
    .X(_05759_));
 sky130_fd_sc_hd__a22oi_2 _06639_ (.A1(reg2_val[18]),
    .A2(net284),
    .B1(net243),
    .B2(_05759_),
    .Y(_05768_));
 sky130_fd_sc_hd__a22o_2 _06640_ (.A1(reg2_val[18]),
    .A2(net284),
    .B1(net243),
    .B2(_05759_),
    .X(_05778_));
 sky130_fd_sc_hd__nand2_1 _06641_ (.A(reg1_val[18]),
    .B(_05768_),
    .Y(_05787_));
 sky130_fd_sc_hd__nand2_1 _06642_ (.A(reg1_val[18]),
    .B(_05778_),
    .Y(_05796_));
 sky130_fd_sc_hd__or2_1 _06643_ (.A(reg1_val[18]),
    .B(_05778_),
    .X(_05805_));
 sky130_fd_sc_hd__and2_1 _06644_ (.A(_05796_),
    .B(_05805_),
    .X(_05814_));
 sky130_fd_sc_hd__o311a_4 _06645_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(net308),
    .B1(instruction[27]),
    .C1(pred_val),
    .X(_05823_));
 sky130_fd_sc_hd__or2_1 _06646_ (.A(net265),
    .B(_05823_),
    .X(_05832_));
 sky130_fd_sc_hd__a22o_2 _06647_ (.A1(reg2_val[17]),
    .A2(net284),
    .B1(net243),
    .B2(_05832_),
    .X(_05840_));
 sky130_fd_sc_hd__inv_2 _06648_ (.A(_05840_),
    .Y(_05850_));
 sky130_fd_sc_hd__nand2_1 _06649_ (.A(reg1_val[17]),
    .B(_05850_),
    .Y(_05859_));
 sky130_fd_sc_hd__and2_1 _06650_ (.A(reg1_val[17]),
    .B(_05840_),
    .X(_05868_));
 sky130_fd_sc_hd__nor2_1 _06651_ (.A(reg1_val[17]),
    .B(_05840_),
    .Y(_05875_));
 sky130_fd_sc_hd__inv_2 _06652_ (.A(_05875_),
    .Y(_05881_));
 sky130_fd_sc_hd__nor2_1 _06653_ (.A(_05868_),
    .B(_05875_),
    .Y(_05887_));
 sky130_fd_sc_hd__o311a_2 _06654_ (.A1(instruction[0]),
    .A2(instruction[1]),
    .A3(net308),
    .B1(instruction[26]),
    .C1(pred_val),
    .X(_05893_));
 sky130_fd_sc_hd__nand2_1 _06655_ (.A(instruction[26]),
    .B(net282),
    .Y(_05899_));
 sky130_fd_sc_hd__nand2_1 _06656_ (.A(_04687_),
    .B(_05899_),
    .Y(_05905_));
 sky130_fd_sc_hd__a22o_2 _06657_ (.A1(reg2_val[16]),
    .A2(net284),
    .B1(net243),
    .B2(_05905_),
    .X(_05911_));
 sky130_fd_sc_hd__inv_2 _06658_ (.A(_05911_),
    .Y(_05922_));
 sky130_fd_sc_hd__nor2_1 _06659_ (.A(_04460_),
    .B(_05911_),
    .Y(_05933_));
 sky130_fd_sc_hd__nor2_1 _06660_ (.A(_04460_),
    .B(_05922_),
    .Y(_05944_));
 sky130_fd_sc_hd__or2_1 _06661_ (.A(reg1_val[16]),
    .B(_05911_),
    .X(_05955_));
 sky130_fd_sc_hd__nand2b_1 _06662_ (.A_N(_05944_),
    .B(_05955_),
    .Y(_05966_));
 sky130_fd_sc_hd__and2_1 _06663_ (.A(reg2_val[15]),
    .B(net283),
    .X(_05977_));
 sky130_fd_sc_hd__a31o_1 _06664_ (.A1(net286),
    .A2(net280),
    .A3(net265),
    .B1(_05977_),
    .X(_05988_));
 sky130_fd_sc_hd__a31oi_4 _06665_ (.A1(net286),
    .A2(net280),
    .A3(net265),
    .B1(_05977_),
    .Y(_05999_));
 sky130_fd_sc_hd__nand2_1 _06666_ (.A(reg1_val[15]),
    .B(_05999_),
    .Y(_06010_));
 sky130_fd_sc_hd__nand2_1 _06667_ (.A(reg1_val[15]),
    .B(_05988_),
    .Y(_06021_));
 sky130_fd_sc_hd__or2_1 _06668_ (.A(reg1_val[15]),
    .B(_05988_),
    .X(_06028_));
 sky130_fd_sc_hd__nand2_2 _06669_ (.A(_06021_),
    .B(_06028_),
    .Y(_06034_));
 sky130_fd_sc_hd__and2_1 _06670_ (.A(reg2_val[14]),
    .B(net283),
    .X(_06040_));
 sky130_fd_sc_hd__a31o_4 _06671_ (.A1(net286),
    .A2(net266),
    .A3(_05024_),
    .B1(_06040_),
    .X(_06046_));
 sky130_fd_sc_hd__and2b_1 _06672_ (.A_N(_06046_),
    .B(reg1_val[14]),
    .X(_06052_));
 sky130_fd_sc_hd__nand2_1 _06673_ (.A(reg1_val[14]),
    .B(_06046_),
    .Y(_06058_));
 sky130_fd_sc_hd__or2_1 _06674_ (.A(reg1_val[14]),
    .B(_06046_),
    .X(_06064_));
 sky130_fd_sc_hd__nand2_2 _06675_ (.A(_06058_),
    .B(_06064_),
    .Y(_06070_));
 sky130_fd_sc_hd__and2_1 _06676_ (.A(reg2_val[13]),
    .B(net283),
    .X(_06076_));
 sky130_fd_sc_hd__a31o_4 _06677_ (.A1(net286),
    .A2(net266),
    .A3(_05165_),
    .B1(_06076_),
    .X(_06082_));
 sky130_fd_sc_hd__nand2b_1 _06678_ (.A_N(_06082_),
    .B(net303),
    .Y(_06088_));
 sky130_fd_sc_hd__nand2_1 _06679_ (.A(net303),
    .B(_06082_),
    .Y(_06094_));
 sky130_fd_sc_hd__or2_1 _06680_ (.A(net303),
    .B(_06082_),
    .X(_06100_));
 sky130_fd_sc_hd__nand2_1 _06681_ (.A(_06094_),
    .B(_06100_),
    .Y(_06109_));
 sky130_fd_sc_hd__and2_1 _06682_ (.A(reg2_val[12]),
    .B(net283),
    .X(_06118_));
 sky130_fd_sc_hd__a31o_4 _06683_ (.A1(net286),
    .A2(net266),
    .A3(_05241_),
    .B1(_06118_),
    .X(_06127_));
 sky130_fd_sc_hd__nand2b_1 _06684_ (.A_N(_06127_),
    .B(reg1_val[12]),
    .Y(_06136_));
 sky130_fd_sc_hd__nand2_1 _06685_ (.A(reg1_val[12]),
    .B(_06127_),
    .Y(_06145_));
 sky130_fd_sc_hd__or2_1 _06686_ (.A(reg1_val[12]),
    .B(_06127_),
    .X(_06154_));
 sky130_fd_sc_hd__nand2_1 _06687_ (.A(_06145_),
    .B(_06154_),
    .Y(_06163_));
 sky130_fd_sc_hd__and2_1 _06688_ (.A(reg2_val[11]),
    .B(net283),
    .X(_06172_));
 sky130_fd_sc_hd__a31o_4 _06689_ (.A1(net286),
    .A2(net266),
    .A3(_04872_),
    .B1(_06172_),
    .X(_06181_));
 sky130_fd_sc_hd__nand2b_1 _06690_ (.A_N(_06181_),
    .B(reg1_val[11]),
    .Y(_06189_));
 sky130_fd_sc_hd__nand2_1 _06691_ (.A(reg1_val[11]),
    .B(_06181_),
    .Y(_06198_));
 sky130_fd_sc_hd__or2_1 _06692_ (.A(reg1_val[11]),
    .B(_06181_),
    .X(_06207_));
 sky130_fd_sc_hd__nand2_2 _06693_ (.A(_06198_),
    .B(_06207_),
    .Y(_06216_));
 sky130_fd_sc_hd__and2_1 _06694_ (.A(reg2_val[10]),
    .B(net283),
    .X(_06225_));
 sky130_fd_sc_hd__a31o_2 _06695_ (.A1(net286),
    .A2(net266),
    .A3(_04807_),
    .B1(_06225_),
    .X(_06233_));
 sky130_fd_sc_hd__nand2b_1 _06696_ (.A_N(_06233_),
    .B(reg1_val[10]),
    .Y(_06240_));
 sky130_fd_sc_hd__nand2_1 _06697_ (.A(reg1_val[10]),
    .B(_06233_),
    .Y(_06241_));
 sky130_fd_sc_hd__or2_1 _06698_ (.A(reg1_val[10]),
    .B(_06233_),
    .X(_06242_));
 sky130_fd_sc_hd__nand2_1 _06699_ (.A(_06241_),
    .B(_06242_),
    .Y(_06243_));
 sky130_fd_sc_hd__and2_1 _06700_ (.A(reg2_val[9]),
    .B(net284),
    .X(_06244_));
 sky130_fd_sc_hd__a31o_1 _06701_ (.A1(net286),
    .A2(net265),
    .A3(_04959_),
    .B1(_06244_),
    .X(_06245_));
 sky130_fd_sc_hd__a31oi_4 _06702_ (.A1(net286),
    .A2(net265),
    .A3(_04959_),
    .B1(_06244_),
    .Y(_06246_));
 sky130_fd_sc_hd__nand2_1 _06703_ (.A(reg1_val[9]),
    .B(_06246_),
    .Y(_06247_));
 sky130_fd_sc_hd__nor2_1 _06704_ (.A(reg1_val[9]),
    .B(_06245_),
    .Y(_06248_));
 sky130_fd_sc_hd__nand2_1 _06705_ (.A(reg1_val[9]),
    .B(_06245_),
    .Y(_06249_));
 sky130_fd_sc_hd__nand2b_1 _06706_ (.A_N(_06248_),
    .B(_06249_),
    .Y(_06250_));
 sky130_fd_sc_hd__and2_1 _06707_ (.A(reg2_val[8]),
    .B(net283),
    .X(_06251_));
 sky130_fd_sc_hd__a31o_4 _06708_ (.A1(net286),
    .A2(net265),
    .A3(_05089_),
    .B1(_06251_),
    .X(_06252_));
 sky130_fd_sc_hd__nand2b_1 _06709_ (.A_N(_06252_),
    .B(reg1_val[8]),
    .Y(_06253_));
 sky130_fd_sc_hd__nor2_1 _06710_ (.A(reg1_val[8]),
    .B(_06252_),
    .Y(_06254_));
 sky130_fd_sc_hd__nand2_1 _06711_ (.A(reg1_val[8]),
    .B(_06252_),
    .Y(_06255_));
 sky130_fd_sc_hd__nand2b_1 _06712_ (.A_N(_06254_),
    .B(_06255_),
    .Y(_06256_));
 sky130_fd_sc_hd__and2_1 _06713_ (.A(reg2_val[7]),
    .B(net283),
    .X(_06257_));
 sky130_fd_sc_hd__a31o_4 _06714_ (.A1(net286),
    .A2(net265),
    .A3(_05350_),
    .B1(_06257_),
    .X(_06258_));
 sky130_fd_sc_hd__and2b_1 _06715_ (.A_N(_06258_),
    .B(reg1_val[7]),
    .X(_06259_));
 sky130_fd_sc_hd__nor2_1 _06716_ (.A(reg1_val[7]),
    .B(_06258_),
    .Y(_06260_));
 sky130_fd_sc_hd__inv_2 _06717_ (.A(_06260_),
    .Y(_06261_));
 sky130_fd_sc_hd__nand2_1 _06718_ (.A(reg1_val[7]),
    .B(_06258_),
    .Y(_06262_));
 sky130_fd_sc_hd__nand2_1 _06719_ (.A(_06261_),
    .B(_06262_),
    .Y(_06263_));
 sky130_fd_sc_hd__and2_1 _06720_ (.A(reg2_val[6]),
    .B(net283),
    .X(_06264_));
 sky130_fd_sc_hd__a31o_4 _06721_ (.A1(net287),
    .A2(net265),
    .A3(_05436_),
    .B1(_06264_),
    .X(_06265_));
 sky130_fd_sc_hd__nand2b_1 _06722_ (.A_N(_06265_),
    .B(reg1_val[6]),
    .Y(_06266_));
 sky130_fd_sc_hd__nor2_1 _06723_ (.A(reg1_val[6]),
    .B(_06265_),
    .Y(_06267_));
 sky130_fd_sc_hd__nand2_1 _06724_ (.A(reg1_val[6]),
    .B(_06265_),
    .Y(_06268_));
 sky130_fd_sc_hd__and2b_1 _06725_ (.A_N(_06267_),
    .B(_06268_),
    .X(_06269_));
 sky130_fd_sc_hd__o2111a_1 _06726_ (.A1(_04427_),
    .A2(_04643_),
    .B1(_04676_),
    .C1(_05512_),
    .D1(net287),
    .X(_06270_));
 sky130_fd_sc_hd__or3b_1 _06727_ (.A(net285),
    .B(_04687_),
    .C_N(_05512_),
    .X(_06271_));
 sky130_fd_sc_hd__a21oi_2 _06728_ (.A1(reg2_val[5]),
    .A2(net284),
    .B1(net264),
    .Y(_06272_));
 sky130_fd_sc_hd__a21o_2 _06729_ (.A1(reg2_val[5]),
    .A2(net284),
    .B1(net264),
    .X(_06273_));
 sky130_fd_sc_hd__nand2_1 _06730_ (.A(reg1_val[5]),
    .B(_06272_),
    .Y(_06274_));
 sky130_fd_sc_hd__nor2_1 _06731_ (.A(reg1_val[5]),
    .B(_06273_),
    .Y(_06275_));
 sky130_fd_sc_hd__or2_1 _06732_ (.A(reg1_val[5]),
    .B(_06273_),
    .X(_06276_));
 sky130_fd_sc_hd__and2_1 _06733_ (.A(reg1_val[5]),
    .B(_06273_),
    .X(_06277_));
 sky130_fd_sc_hd__nor2_1 _06734_ (.A(_06275_),
    .B(_06277_),
    .Y(_06278_));
 sky130_fd_sc_hd__and2_1 _06735_ (.A(reg2_val[4]),
    .B(net283),
    .X(_06279_));
 sky130_fd_sc_hd__a31o_1 _06736_ (.A1(net286),
    .A2(net265),
    .A3(_05591_),
    .B1(_06279_),
    .X(_06280_));
 sky130_fd_sc_hd__a31oi_4 _06737_ (.A1(net286),
    .A2(net265),
    .A3(_05591_),
    .B1(_06279_),
    .Y(_06281_));
 sky130_fd_sc_hd__nor2_1 _06738_ (.A(_04449_),
    .B(net240),
    .Y(_06282_));
 sky130_fd_sc_hd__nor2_1 _06739_ (.A(reg1_val[4]),
    .B(net240),
    .Y(_06283_));
 sky130_fd_sc_hd__nand2_1 _06740_ (.A(reg1_val[4]),
    .B(net240),
    .Y(_06284_));
 sky130_fd_sc_hd__nand2b_2 _06741_ (.A_N(_06283_),
    .B(_06284_),
    .Y(_06285_));
 sky130_fd_sc_hd__and2_1 _06742_ (.A(reg2_val[3]),
    .B(net283),
    .X(_06286_));
 sky130_fd_sc_hd__a31o_4 _06743_ (.A1(net286),
    .A2(net265),
    .A3(_05677_),
    .B1(_06286_),
    .X(_06287_));
 sky130_fd_sc_hd__and2b_1 _06744_ (.A_N(_06287_),
    .B(reg1_val[3]),
    .X(_06288_));
 sky130_fd_sc_hd__nor2_1 _06745_ (.A(reg1_val[3]),
    .B(_06287_),
    .Y(_06289_));
 sky130_fd_sc_hd__nand2_1 _06746_ (.A(reg1_val[3]),
    .B(_06287_),
    .Y(_06290_));
 sky130_fd_sc_hd__nand2b_2 _06747_ (.A_N(_06289_),
    .B(_06290_),
    .Y(_06291_));
 sky130_fd_sc_hd__and2_1 _06748_ (.A(reg2_val[2]),
    .B(net283),
    .X(_06292_));
 sky130_fd_sc_hd__a31o_1 _06749_ (.A1(net286),
    .A2(net265),
    .A3(_05750_),
    .B1(_06292_),
    .X(_06293_));
 sky130_fd_sc_hd__and2b_1 _06750_ (.A_N(net233),
    .B(reg1_val[2]),
    .X(_06294_));
 sky130_fd_sc_hd__xnor2_2 _06751_ (.A(reg1_val[2]),
    .B(net233),
    .Y(_06295_));
 sky130_fd_sc_hd__o211ai_4 _06752_ (.A1(_04427_),
    .A2(_04643_),
    .B1(_04676_),
    .C1(_05823_),
    .Y(_06296_));
 sky130_fd_sc_hd__nor2_1 _06753_ (.A(reg2_val[1]),
    .B(net287),
    .Y(_06297_));
 sky130_fd_sc_hd__and2_1 _06754_ (.A(reg2_val[1]),
    .B(net285),
    .X(_06298_));
 sky130_fd_sc_hd__a21oi_4 _06755_ (.A1(net287),
    .A2(_06296_),
    .B1(_06297_),
    .Y(_06299_));
 sky130_fd_sc_hd__a21o_1 _06756_ (.A1(net287),
    .A2(_06296_),
    .B1(_06297_),
    .X(_06300_));
 sky130_fd_sc_hd__nand2_1 _06757_ (.A(reg1_val[1]),
    .B(net229),
    .Y(_06301_));
 sky130_fd_sc_hd__a211o_1 _06758_ (.A1(net287),
    .A2(_06296_),
    .B1(_06297_),
    .C1(_04438_),
    .X(_06302_));
 sky130_fd_sc_hd__a311oi_2 _06759_ (.A1(net287),
    .A2(_04698_),
    .A3(_05823_),
    .B1(_06298_),
    .C1(reg1_val[1]),
    .Y(_06303_));
 sky130_fd_sc_hd__a311o_1 _06760_ (.A1(net287),
    .A2(_04698_),
    .A3(_05823_),
    .B1(_06298_),
    .C1(reg1_val[1]),
    .X(_06304_));
 sky130_fd_sc_hd__nand2_1 _06761_ (.A(_06302_),
    .B(_06304_),
    .Y(_06305_));
 sky130_fd_sc_hd__o211a_2 _06762_ (.A1(_04427_),
    .A2(_04643_),
    .B1(_04676_),
    .C1(_05893_),
    .X(_06306_));
 sky130_fd_sc_hd__or2_2 _06763_ (.A(reg2_val[0]),
    .B(net286),
    .X(_06307_));
 sky130_fd_sc_hd__o21a_1 _06764_ (.A1(net284),
    .A2(_06306_),
    .B1(_06307_),
    .X(_06308_));
 sky130_fd_sc_hd__o21ai_4 _06765_ (.A1(net284),
    .A2(_06306_),
    .B1(_06307_),
    .Y(_06309_));
 sky130_fd_sc_hd__a22o_1 _06766_ (.A1(_06302_),
    .A2(_06304_),
    .B1(net227),
    .B2(_04416_),
    .X(_06310_));
 sky130_fd_sc_hd__a21boi_1 _06767_ (.A1(_06301_),
    .A2(_06310_),
    .B1_N(_06295_),
    .Y(_06311_));
 sky130_fd_sc_hd__o21a_1 _06768_ (.A1(_06294_),
    .A2(_06311_),
    .B1(_06291_),
    .X(_06312_));
 sky130_fd_sc_hd__o21a_1 _06769_ (.A1(_06288_),
    .A2(_06312_),
    .B1(_06285_),
    .X(_06313_));
 sky130_fd_sc_hd__o21bai_1 _06770_ (.A1(_06282_),
    .A2(_06313_),
    .B1_N(_06278_),
    .Y(_06314_));
 sky130_fd_sc_hd__a21o_1 _06771_ (.A1(_06274_),
    .A2(_06314_),
    .B1(_06269_),
    .X(_06315_));
 sky130_fd_sc_hd__nand2_1 _06772_ (.A(_06266_),
    .B(_06315_),
    .Y(_06316_));
 sky130_fd_sc_hd__a21boi_1 _06773_ (.A1(_06266_),
    .A2(_06315_),
    .B1_N(_06263_),
    .Y(_06317_));
 sky130_fd_sc_hd__o21ai_1 _06774_ (.A1(_06259_),
    .A2(_06317_),
    .B1(_06256_),
    .Y(_06318_));
 sky130_fd_sc_hd__nand2_1 _06775_ (.A(_06253_),
    .B(_06318_),
    .Y(_06319_));
 sky130_fd_sc_hd__a21bo_1 _06776_ (.A1(_06253_),
    .A2(_06318_),
    .B1_N(_06250_),
    .X(_06320_));
 sky130_fd_sc_hd__nand2_1 _06777_ (.A(_06247_),
    .B(_06320_),
    .Y(_06321_));
 sky130_fd_sc_hd__a21bo_1 _06778_ (.A1(_06247_),
    .A2(_06320_),
    .B1_N(_06243_),
    .X(_06322_));
 sky130_fd_sc_hd__a21bo_1 _06779_ (.A1(_06240_),
    .A2(_06322_),
    .B1_N(_06216_),
    .X(_06323_));
 sky130_fd_sc_hd__a21bo_1 _06780_ (.A1(_06189_),
    .A2(_06323_),
    .B1_N(_06163_),
    .X(_06324_));
 sky130_fd_sc_hd__a21bo_1 _06781_ (.A1(_06136_),
    .A2(_06324_),
    .B1_N(_06109_),
    .X(_06325_));
 sky130_fd_sc_hd__a21boi_1 _06782_ (.A1(_06088_),
    .A2(_06325_),
    .B1_N(_06070_),
    .Y(_06326_));
 sky130_fd_sc_hd__o21ai_1 _06783_ (.A1(_06052_),
    .A2(_06326_),
    .B1(_06034_),
    .Y(_06327_));
 sky130_fd_sc_hd__a21boi_1 _06784_ (.A1(_06010_),
    .A2(_06327_),
    .B1_N(_05966_),
    .Y(_06328_));
 sky130_fd_sc_hd__nor2_1 _06785_ (.A(_05933_),
    .B(_06328_),
    .Y(_06329_));
 sky130_fd_sc_hd__o21bai_1 _06786_ (.A1(_05933_),
    .A2(_06328_),
    .B1_N(_05887_),
    .Y(_06330_));
 sky130_fd_sc_hd__and2_1 _06787_ (.A(_05859_),
    .B(_06330_),
    .X(_06331_));
 sky130_fd_sc_hd__a21o_1 _06788_ (.A1(_05859_),
    .A2(_06330_),
    .B1(_05814_),
    .X(_06332_));
 sky130_fd_sc_hd__a21o_1 _06789_ (.A1(_05787_),
    .A2(_06332_),
    .B1(_05741_),
    .X(_06333_));
 sky130_fd_sc_hd__and2_1 _06790_ (.A(_05715_),
    .B(_06333_),
    .X(_06334_));
 sky130_fd_sc_hd__a21o_1 _06791_ (.A1(_05715_),
    .A2(_06333_),
    .B1(_05668_),
    .X(_06335_));
 sky130_fd_sc_hd__and2_1 _06792_ (.A(_05630_),
    .B(_06335_),
    .X(_06336_));
 sky130_fd_sc_hd__a21o_1 _06793_ (.A1(_05630_),
    .A2(_06335_),
    .B1(_05582_),
    .X(_06337_));
 sky130_fd_sc_hd__and2_1 _06794_ (.A(_05553_),
    .B(_06337_),
    .X(_06338_));
 sky130_fd_sc_hd__a21o_1 _06795_ (.A1(_05553_),
    .A2(_06337_),
    .B1(_05501_),
    .X(_06339_));
 sky130_fd_sc_hd__and2_1 _06796_ (.A(_05469_),
    .B(_06339_),
    .X(_06340_));
 sky130_fd_sc_hd__a21o_1 _06797_ (.A1(_05469_),
    .A2(_06339_),
    .B1(_05425_),
    .X(_06341_));
 sky130_fd_sc_hd__and2_1 _06798_ (.A(_05393_),
    .B(_06341_),
    .X(_06342_));
 sky130_fd_sc_hd__and2b_1 _06799_ (.A_N(_06342_),
    .B(_05339_),
    .X(_06343_));
 sky130_fd_sc_hd__or2_1 _06800_ (.A(_04493_),
    .B(_05046_),
    .X(_06344_));
 sky130_fd_sc_hd__nand2_1 _06801_ (.A(reg1_val[29]),
    .B(_05187_),
    .Y(_06345_));
 sky130_fd_sc_hd__nand2_1 _06802_ (.A(reg1_val[28]),
    .B(_05274_),
    .Y(_06346_));
 sky130_fd_sc_hd__nand2_1 _06803_ (.A(reg1_val[27]),
    .B(_04904_),
    .Y(_06347_));
 sky130_fd_sc_hd__or2_1 _06804_ (.A(_04482_),
    .B(_04828_),
    .X(_06348_));
 sky130_fd_sc_hd__nand2_1 _06805_ (.A(reg1_val[25]),
    .B(_04980_),
    .Y(_06349_));
 sky130_fd_sc_hd__nand2_1 _06806_ (.A(reg1_val[24]),
    .B(_05111_),
    .Y(_06350_));
 sky130_fd_sc_hd__o21a_1 _06807_ (.A1(_05013_),
    .A2(_06350_),
    .B1(_06349_),
    .X(_06351_));
 sky130_fd_sc_hd__o21a_1 _06808_ (.A1(_04861_),
    .A2(_06351_),
    .B1(_06348_),
    .X(_06352_));
 sky130_fd_sc_hd__o21a_1 _06809_ (.A1(_04948_),
    .A2(_06352_),
    .B1(_06347_),
    .X(_06353_));
 sky130_fd_sc_hd__o21a_1 _06810_ (.A1(_05306_),
    .A2(_06353_),
    .B1(_06346_),
    .X(_06354_));
 sky130_fd_sc_hd__o21a_1 _06811_ (.A1(_05230_),
    .A2(_06354_),
    .B1(_06345_),
    .X(_06355_));
 sky130_fd_sc_hd__o21ai_1 _06812_ (.A1(_05078_),
    .A2(_06355_),
    .B1(_06344_),
    .Y(_06356_));
 sky130_fd_sc_hd__a2111o_1 _06813_ (.A1(_04796_),
    .A2(_06356_),
    .B1(_06343_),
    .C1(instruction[6]),
    .D1(_04763_),
    .X(_06357_));
 sky130_fd_sc_hd__a21o_1 _06814_ (.A1(_05393_),
    .A2(_06341_),
    .B1(_05154_),
    .X(_06358_));
 sky130_fd_sc_hd__a21o_1 _06815_ (.A1(_06350_),
    .A2(_06358_),
    .B1(_05013_),
    .X(_06359_));
 sky130_fd_sc_hd__a21o_1 _06816_ (.A1(_06349_),
    .A2(_06359_),
    .B1(_04861_),
    .X(_06360_));
 sky130_fd_sc_hd__a21o_1 _06817_ (.A1(_06348_),
    .A2(_06360_),
    .B1(_04948_),
    .X(_06361_));
 sky130_fd_sc_hd__a21o_1 _06818_ (.A1(_06347_),
    .A2(_06361_),
    .B1(_05306_),
    .X(_06362_));
 sky130_fd_sc_hd__and2_1 _06819_ (.A(_06346_),
    .B(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__a21o_1 _06820_ (.A1(_06346_),
    .A2(_06362_),
    .B1(_05230_),
    .X(_06364_));
 sky130_fd_sc_hd__and2_1 _06821_ (.A(_06345_),
    .B(_06364_),
    .X(_06365_));
 sky130_fd_sc_hd__a21o_1 _06822_ (.A1(_06345_),
    .A2(_06364_),
    .B1(_05078_),
    .X(_06366_));
 sky130_fd_sc_hd__nand2_1 _06823_ (.A(_06344_),
    .B(_06366_),
    .Y(_06367_));
 sky130_fd_sc_hd__a31o_1 _06824_ (.A1(_04796_),
    .A2(_06344_),
    .A3(_06366_),
    .B1(_04763_),
    .X(_06368_));
 sky130_fd_sc_hd__a21bo_1 _06825_ (.A1(instruction[6]),
    .A2(_06368_),
    .B1_N(_06357_),
    .X(_06369_));
 sky130_fd_sc_hd__or2_4 _06826_ (.A(instruction[3]),
    .B(instruction[4]),
    .X(_06370_));
 sky130_fd_sc_hd__o211ai_4 _06827_ (.A1(net284),
    .A2(_06306_),
    .B1(_06307_),
    .C1(net304),
    .Y(_06371_));
 sky130_fd_sc_hd__nand2_1 _06828_ (.A(net302),
    .B(net226),
    .Y(_06372_));
 sky130_fd_sc_hd__nand2_1 _06829_ (.A(_06371_),
    .B(_06372_),
    .Y(_06373_));
 sky130_fd_sc_hd__and4_1 _06830_ (.A(_06216_),
    .B(_06243_),
    .C(_06250_),
    .D(_06263_),
    .X(_06374_));
 sky130_fd_sc_hd__and4_1 _06831_ (.A(_06034_),
    .B(_06070_),
    .C(_06109_),
    .D(_06163_),
    .X(_06375_));
 sky130_fd_sc_hd__nor2_1 _06832_ (.A(_06269_),
    .B(_06278_),
    .Y(_06376_));
 sky130_fd_sc_hd__and4_1 _06833_ (.A(_06256_),
    .B(_06295_),
    .C(_06305_),
    .D(_06373_),
    .X(_06377_));
 sky130_fd_sc_hd__and4_1 _06834_ (.A(_06285_),
    .B(_06291_),
    .C(_06376_),
    .D(_06377_),
    .X(_06378_));
 sky130_fd_sc_hd__and3_1 _06835_ (.A(_06374_),
    .B(_06375_),
    .C(_06378_),
    .X(_06379_));
 sky130_fd_sc_hd__or4b_1 _06836_ (.A(_05741_),
    .B(_05814_),
    .C(_05887_),
    .D_N(_05966_),
    .X(_06380_));
 sky130_fd_sc_hd__or4_1 _06837_ (.A(_05425_),
    .B(_05501_),
    .C(_05582_),
    .D(_05668_),
    .X(_06381_));
 sky130_fd_sc_hd__nor2_1 _06838_ (.A(_06380_),
    .B(_06381_),
    .Y(_06382_));
 sky130_fd_sc_hd__and3_1 _06839_ (.A(_05339_),
    .B(_06379_),
    .C(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__a21oi_1 _06840_ (.A1(instruction[6]),
    .A2(_04785_),
    .B1(_06370_),
    .Y(_06384_));
 sky130_fd_sc_hd__o21a_1 _06841_ (.A1(instruction[6]),
    .A2(_06383_),
    .B1(_06384_),
    .X(_06385_));
 sky130_fd_sc_hd__nand2_4 _06842_ (.A(instruction[3]),
    .B(instruction[4]),
    .Y(_06386_));
 sky130_fd_sc_hd__inv_2 _06843_ (.A(_06386_),
    .Y(_06387_));
 sky130_fd_sc_hd__or2_2 _06844_ (.A(_04406_),
    .B(instruction[4]),
    .X(_06388_));
 sky130_fd_sc_hd__a221o_2 _06845_ (.A1(instruction[3]),
    .A2(_06369_),
    .B1(_06383_),
    .B2(_06387_),
    .C1(_06385_),
    .X(_06389_));
 sky130_fd_sc_hd__xor2_4 _06846_ (.A(instruction[5]),
    .B(_06389_),
    .X(dest_pred_val));
 sky130_fd_sc_hd__and2_4 _06847_ (.A(net308),
    .B(_04567_),
    .X(_06390_));
 sky130_fd_sc_hd__nand2_2 _06848_ (.A(net308),
    .B(_04567_),
    .Y(_06391_));
 sky130_fd_sc_hd__and4b_4 _06849_ (.A_N(instruction[1]),
    .B(net308),
    .C(instruction[0]),
    .D(pred_val),
    .X(_06392_));
 sky130_fd_sc_hd__nand4b_4 _06850_ (.A_N(instruction[1]),
    .B(net308),
    .C(instruction[0]),
    .D(pred_val),
    .Y(_06393_));
 sky130_fd_sc_hd__a21o_4 _06851_ (.A1(dest_pred_val),
    .A2(_06392_),
    .B1(_06390_),
    .X(take_branch));
 sky130_fd_sc_hd__a21oi_1 _06852_ (.A1(instruction[6]),
    .A2(instruction[5]),
    .B1(instruction[4]),
    .Y(_06394_));
 sky130_fd_sc_hd__nand2b_4 _06853_ (.A_N(instruction[5]),
    .B(instruction[6]),
    .Y(_06395_));
 sky130_fd_sc_hd__a221oi_2 _06854_ (.A1(net285),
    .A2(_04643_),
    .B1(_06395_),
    .B2(instruction[4]),
    .C1(_06394_),
    .Y(_06396_));
 sky130_fd_sc_hd__a221o_1 _06855_ (.A1(net285),
    .A2(_04643_),
    .B1(_06395_),
    .B2(instruction[4]),
    .C1(_06394_),
    .X(_06397_));
 sky130_fd_sc_hd__nor2_1 _06856_ (.A(net272),
    .B(_06396_),
    .Y(_06398_));
 sky130_fd_sc_hd__nand2_1 _06857_ (.A(net267),
    .B(_06397_),
    .Y(_06399_));
 sky130_fd_sc_hd__nor2_8 _06858_ (.A(div_complete),
    .B(net222),
    .Y(busy));
 sky130_fd_sc_hd__and4b_4 _06859_ (.A_N(net308),
    .B(instruction[1]),
    .C(pred_val),
    .D(instruction[0]),
    .X(_06400_));
 sky130_fd_sc_hd__and2_4 _06860_ (.A(instruction[11]),
    .B(_06400_),
    .X(dest_pred[0]));
 sky130_fd_sc_hd__and2_4 _06861_ (.A(instruction[12]),
    .B(_06400_),
    .X(dest_pred[1]));
 sky130_fd_sc_hd__and2_4 _06862_ (.A(instruction[13]),
    .B(_06400_),
    .X(dest_pred[2]));
 sky130_fd_sc_hd__or2_2 _06863_ (.A(_04567_),
    .B(_04632_),
    .X(_06401_));
 sky130_fd_sc_hd__and2_4 _06864_ (.A(instruction[11]),
    .B(_06401_),
    .X(dest_idx[0]));
 sky130_fd_sc_hd__and2_4 _06865_ (.A(instruction[12]),
    .B(_06401_),
    .X(dest_idx[1]));
 sky130_fd_sc_hd__and2_4 _06866_ (.A(instruction[13]),
    .B(_06401_),
    .X(dest_idx[2]));
 sky130_fd_sc_hd__and2_4 _06867_ (.A(instruction[14]),
    .B(_06401_),
    .X(dest_idx[3]));
 sky130_fd_sc_hd__and2_4 _06868_ (.A(instruction[15]),
    .B(_06401_),
    .X(dest_idx[4]));
 sky130_fd_sc_hd__or2_1 _06869_ (.A(instruction[18]),
    .B(_06392_),
    .X(_06402_));
 sky130_fd_sc_hd__o211a_4 _06870_ (.A1(instruction[11]),
    .A2(_06393_),
    .B1(_06402_),
    .C1(net282),
    .X(reg1_idx[0]));
 sky130_fd_sc_hd__or2_1 _06871_ (.A(instruction[19]),
    .B(_06392_),
    .X(_06403_));
 sky130_fd_sc_hd__o211a_4 _06872_ (.A1(instruction[12]),
    .A2(_06393_),
    .B1(_06403_),
    .C1(net282),
    .X(reg1_idx[1]));
 sky130_fd_sc_hd__or2_1 _06873_ (.A(instruction[20]),
    .B(_06392_),
    .X(_06404_));
 sky130_fd_sc_hd__o211a_4 _06874_ (.A1(instruction[13]),
    .A2(_06393_),
    .B1(_06404_),
    .C1(net282),
    .X(reg1_idx[2]));
 sky130_fd_sc_hd__or2_1 _06875_ (.A(instruction[21]),
    .B(_06392_),
    .X(_06405_));
 sky130_fd_sc_hd__o211a_4 _06876_ (.A1(instruction[14]),
    .A2(_06393_),
    .B1(_06405_),
    .C1(net282),
    .X(reg1_idx[3]));
 sky130_fd_sc_hd__or2_1 _06877_ (.A(instruction[22]),
    .B(_06392_),
    .X(_06406_));
 sky130_fd_sc_hd__o211a_4 _06878_ (.A1(instruction[15]),
    .A2(_06393_),
    .B1(_06406_),
    .C1(net282),
    .X(reg1_idx[4]));
 sky130_fd_sc_hd__or2_1 _06879_ (.A(instruction[25]),
    .B(_06392_),
    .X(_06407_));
 sky130_fd_sc_hd__o211a_4 _06880_ (.A1(instruction[18]),
    .A2(_06393_),
    .B1(_06407_),
    .C1(net281),
    .X(reg2_idx[0]));
 sky130_fd_sc_hd__or2_1 _06881_ (.A(instruction[26]),
    .B(_06392_),
    .X(_06408_));
 sky130_fd_sc_hd__o211a_4 _06882_ (.A1(instruction[19]),
    .A2(_06393_),
    .B1(_06408_),
    .C1(net281),
    .X(reg2_idx[1]));
 sky130_fd_sc_hd__or2_1 _06883_ (.A(instruction[27]),
    .B(_06392_),
    .X(_06409_));
 sky130_fd_sc_hd__o211a_4 _06884_ (.A1(instruction[20]),
    .A2(_06393_),
    .B1(_06409_),
    .C1(net281),
    .X(reg2_idx[2]));
 sky130_fd_sc_hd__or2_1 _06885_ (.A(instruction[28]),
    .B(_06392_),
    .X(_06410_));
 sky130_fd_sc_hd__o211a_4 _06886_ (.A1(instruction[21]),
    .A2(_06393_),
    .B1(_06410_),
    .C1(net281),
    .X(reg2_idx[3]));
 sky130_fd_sc_hd__or2_1 _06887_ (.A(instruction[29]),
    .B(_06392_),
    .X(_06411_));
 sky130_fd_sc_hd__o211a_4 _06888_ (.A1(instruction[22]),
    .A2(_06393_),
    .B1(_06411_),
    .C1(net281),
    .X(reg2_idx[4]));
 sky130_fd_sc_hd__nor3_4 _06889_ (.A(instruction[6]),
    .B(instruction[5]),
    .C(_06388_),
    .Y(_06412_));
 sky130_fd_sc_hd__or3_4 _06890_ (.A(instruction[6]),
    .B(instruction[5]),
    .C(_06388_),
    .X(_06413_));
 sky130_fd_sc_hd__or2_1 _06891_ (.A(instruction[6]),
    .B(instruction[5]),
    .X(_06414_));
 sky130_fd_sc_hd__nand2_2 _06892_ (.A(_04406_),
    .B(instruction[4]),
    .Y(_06415_));
 sky130_fd_sc_hd__nor2_1 _06893_ (.A(_06414_),
    .B(_06415_),
    .Y(_06416_));
 sky130_fd_sc_hd__or2_2 _06894_ (.A(_06414_),
    .B(_06415_),
    .X(_06417_));
 sky130_fd_sc_hd__a31o_1 _06895_ (.A1(instruction[17]),
    .A2(_06413_),
    .A3(_06417_),
    .B1(_04589_),
    .X(_06418_));
 sky130_fd_sc_hd__nor2_1 _06896_ (.A(instruction[6]),
    .B(is_load),
    .Y(_06419_));
 sky130_fd_sc_hd__o211a_1 _06897_ (.A1(instruction[40]),
    .A2(_04643_),
    .B1(_06418_),
    .C1(_06419_),
    .X(_06420_));
 sky130_fd_sc_hd__a32o_2 _06898_ (.A1(instruction[24]),
    .A2(net307),
    .A3(is_load),
    .B1(_04687_),
    .B2(_06420_),
    .X(_06421_));
 sky130_fd_sc_hd__nand2_8 _06899_ (.A(net261),
    .B(_06421_),
    .Y(dest_mask[0]));
 sky130_fd_sc_hd__a22o_2 _06900_ (.A1(net307),
    .A2(is_load),
    .B1(net266),
    .B2(_06420_),
    .X(_06422_));
 sky130_fd_sc_hd__nand2_8 _06901_ (.A(net261),
    .B(_06422_),
    .Y(dest_mask[1]));
 sky130_fd_sc_hd__nand2b_4 _06902_ (.A_N(instruction[6]),
    .B(instruction[5]),
    .Y(_06423_));
 sky130_fd_sc_hd__nor2_2 _06903_ (.A(_06370_),
    .B(_06423_),
    .Y(_06424_));
 sky130_fd_sc_hd__and2_1 _06904_ (.A(net305),
    .B(_06424_),
    .X(_06425_));
 sky130_fd_sc_hd__nand2_8 _06905_ (.A(net306),
    .B(_06424_),
    .Y(_06426_));
 sky130_fd_sc_hd__a21oi_4 _06906_ (.A1(instruction[6]),
    .A2(instruction[5]),
    .B1(net212),
    .Y(_06427_));
 sky130_fd_sc_hd__inv_2 _06907_ (.A(_06427_),
    .Y(_06428_));
 sky130_fd_sc_hd__and2_1 _06908_ (.A(reg1_val[31]),
    .B(net307),
    .X(_06429_));
 sky130_fd_sc_hd__or4_2 _06909_ (.A(net304),
    .B(reg1_val[1]),
    .C(reg1_val[2]),
    .D(reg1_val[3]),
    .X(_06430_));
 sky130_fd_sc_hd__or4_2 _06910_ (.A(reg1_val[4]),
    .B(reg1_val[5]),
    .C(reg1_val[6]),
    .D(_06430_),
    .X(_06431_));
 sky130_fd_sc_hd__or4_2 _06911_ (.A(reg1_val[7]),
    .B(reg1_val[8]),
    .C(reg1_val[9]),
    .D(_06431_),
    .X(_06432_));
 sky130_fd_sc_hd__or4_4 _06912_ (.A(reg1_val[10]),
    .B(reg1_val[11]),
    .C(reg1_val[12]),
    .D(_06432_),
    .X(_06433_));
 sky130_fd_sc_hd__and2_2 _06913_ (.A(net274),
    .B(_06433_),
    .X(_06434_));
 sky130_fd_sc_hd__xor2_4 _06914_ (.A(net303),
    .B(_06434_),
    .X(_06435_));
 sky130_fd_sc_hd__xnor2_1 _06915_ (.A(net303),
    .B(_06434_),
    .Y(_06436_));
 sky130_fd_sc_hd__o21a_1 _06916_ (.A1(reg1_val[10]),
    .A2(_06432_),
    .B1(net275),
    .X(_06437_));
 sky130_fd_sc_hd__xnor2_2 _06917_ (.A(reg1_val[11]),
    .B(_06437_),
    .Y(_06438_));
 sky130_fd_sc_hd__o31a_2 _06918_ (.A1(reg1_val[10]),
    .A2(reg1_val[11]),
    .A3(_06432_),
    .B1(net275),
    .X(_06439_));
 sky130_fd_sc_hd__xnor2_4 _06919_ (.A(reg1_val[12]),
    .B(_06439_),
    .Y(_06440_));
 sky130_fd_sc_hd__nor2_1 _06920_ (.A(net179),
    .B(_06440_),
    .Y(_06441_));
 sky130_fd_sc_hd__and2_1 _06921_ (.A(net157),
    .B(_06441_),
    .X(_06442_));
 sky130_fd_sc_hd__and2_1 _06922_ (.A(net179),
    .B(_06440_),
    .X(_06443_));
 sky130_fd_sc_hd__a21oi_1 _06923_ (.A1(_06435_),
    .A2(_06443_),
    .B1(_06442_),
    .Y(_06444_));
 sky130_fd_sc_hd__a21o_1 _06924_ (.A1(_06435_),
    .A2(_06443_),
    .B1(_06442_),
    .X(_06445_));
 sky130_fd_sc_hd__and2_1 _06925_ (.A(net307),
    .B(_04752_),
    .X(_06446_));
 sky130_fd_sc_hd__nand2_2 _06926_ (.A(net307),
    .B(_04752_),
    .Y(_06447_));
 sky130_fd_sc_hd__or4_4 _06927_ (.A(_06287_),
    .B(net233),
    .C(_06299_),
    .D(net227),
    .X(_06448_));
 sky130_fd_sc_hd__or4_2 _06928_ (.A(_06258_),
    .B(_06265_),
    .C(_06273_),
    .D(net240),
    .X(_06449_));
 sky130_fd_sc_hd__nor2_2 _06929_ (.A(_06448_),
    .B(_06449_),
    .Y(_06450_));
 sky130_fd_sc_hd__or3_1 _06930_ (.A(_06252_),
    .B(_06448_),
    .C(_06449_),
    .X(_06451_));
 sky130_fd_sc_hd__or2_1 _06931_ (.A(_06233_),
    .B(_06245_),
    .X(_06452_));
 sky130_fd_sc_hd__or4_2 _06932_ (.A(_06252_),
    .B(_06448_),
    .C(_06449_),
    .D(_06452_),
    .X(_06453_));
 sky130_fd_sc_hd__o41a_4 _06933_ (.A1(_06082_),
    .A2(_06127_),
    .A3(_06181_),
    .A4(_06453_),
    .B1(net193),
    .X(_06454_));
 sky130_fd_sc_hd__and3_1 _06934_ (.A(net306),
    .B(_04752_),
    .C(_06046_),
    .X(_06455_));
 sky130_fd_sc_hd__o21ai_4 _06935_ (.A1(_06454_),
    .A2(_06455_),
    .B1(_05999_),
    .Y(_06456_));
 sky130_fd_sc_hd__or3_4 _06936_ (.A(_05999_),
    .B(_06454_),
    .C(_06455_),
    .X(_06457_));
 sky130_fd_sc_hd__and2_1 _06937_ (.A(_06456_),
    .B(_06457_),
    .X(_06458_));
 sky130_fd_sc_hd__nand2_4 _06938_ (.A(_06456_),
    .B(_06457_),
    .Y(_06459_));
 sky130_fd_sc_hd__or2_2 _06939_ (.A(_06441_),
    .B(_06443_),
    .X(_06460_));
 sky130_fd_sc_hd__inv_2 _06940_ (.A(net130),
    .Y(_06461_));
 sky130_fd_sc_hd__or4_1 _06941_ (.A(_05988_),
    .B(_06046_),
    .C(_06082_),
    .D(_06127_),
    .X(_06462_));
 sky130_fd_sc_hd__nor4_2 _06942_ (.A(_06181_),
    .B(_06252_),
    .C(_06452_),
    .D(_06462_),
    .Y(_06463_));
 sky130_fd_sc_hd__nand2_1 _06943_ (.A(_06450_),
    .B(_06463_),
    .Y(_06464_));
 sky130_fd_sc_hd__a21oi_1 _06944_ (.A1(_06450_),
    .A2(_06463_),
    .B1(_06447_),
    .Y(_06465_));
 sky130_fd_sc_hd__nor2_1 _06945_ (.A(_05922_),
    .B(_06447_),
    .Y(_06466_));
 sky130_fd_sc_hd__o2bb2a_2 _06946_ (.A1_N(_06464_),
    .A2_N(_06466_),
    .B1(_06465_),
    .B2(_05911_),
    .X(_06467_));
 sky130_fd_sc_hd__a2bb2o_2 _06947_ (.A1_N(_05911_),
    .A2_N(_06465_),
    .B1(_06466_),
    .B2(_06464_),
    .X(_06468_));
 sky130_fd_sc_hd__o22a_1 _06948_ (.A1(net82),
    .A2(net80),
    .B1(net130),
    .B2(net128),
    .X(_06469_));
 sky130_fd_sc_hd__xnor2_1 _06949_ (.A(net158),
    .B(_06469_),
    .Y(_06470_));
 sky130_fd_sc_hd__o21a_1 _06950_ (.A1(net303),
    .A2(_06433_),
    .B1(net274),
    .X(_06471_));
 sky130_fd_sc_hd__o31a_1 _06951_ (.A1(net303),
    .A2(reg1_val[14]),
    .A3(_06433_),
    .B1(net274),
    .X(_06472_));
 sky130_fd_sc_hd__xor2_1 _06952_ (.A(reg1_val[15]),
    .B(_06472_),
    .X(_06473_));
 sky130_fd_sc_hd__xnor2_4 _06953_ (.A(reg1_val[14]),
    .B(_06471_),
    .Y(_06474_));
 sky130_fd_sc_hd__or3_1 _06954_ (.A(net157),
    .B(net155),
    .C(_06474_),
    .X(_06475_));
 sky130_fd_sc_hd__nand2_1 _06955_ (.A(net157),
    .B(_06474_),
    .Y(_06476_));
 sky130_fd_sc_hd__nand3_1 _06956_ (.A(net157),
    .B(net155),
    .C(_06474_),
    .Y(_06477_));
 sky130_fd_sc_hd__and2_1 _06957_ (.A(_06475_),
    .B(_06477_),
    .X(_06478_));
 sky130_fd_sc_hd__o21a_2 _06958_ (.A1(_06181_),
    .A2(_06453_),
    .B1(net193),
    .X(_06479_));
 sky130_fd_sc_hd__o31a_1 _06959_ (.A1(_06127_),
    .A2(_06181_),
    .A3(_06453_),
    .B1(net193),
    .X(_06480_));
 sky130_fd_sc_hd__xnor2_1 _06960_ (.A(_06082_),
    .B(_06480_),
    .Y(_06481_));
 sky130_fd_sc_hd__xnor2_4 _06961_ (.A(net157),
    .B(_06474_),
    .Y(_06482_));
 sky130_fd_sc_hd__xor2_4 _06962_ (.A(_06046_),
    .B(_06454_),
    .X(_06483_));
 sky130_fd_sc_hd__xnor2_4 _06963_ (.A(_06046_),
    .B(_06454_),
    .Y(_06484_));
 sky130_fd_sc_hd__o22a_1 _06964_ (.A1(net79),
    .A2(net127),
    .B1(net124),
    .B2(net121),
    .X(_06485_));
 sky130_fd_sc_hd__xor2_1 _06965_ (.A(net155),
    .B(_06485_),
    .X(_06486_));
 sky130_fd_sc_hd__nor2_1 _06966_ (.A(_06470_),
    .B(_06486_),
    .Y(_06487_));
 sky130_fd_sc_hd__o31a_2 _06967_ (.A1(reg1_val[7]),
    .A2(reg1_val[8]),
    .A3(_06431_),
    .B1(net275),
    .X(_06488_));
 sky130_fd_sc_hd__xnor2_4 _06968_ (.A(reg1_val[9]),
    .B(_06488_),
    .Y(_06489_));
 sky130_fd_sc_hd__inv_6 _06969_ (.A(net191),
    .Y(_06490_));
 sky130_fd_sc_hd__nand2_1 _06970_ (.A(net275),
    .B(_06431_),
    .Y(_06491_));
 sky130_fd_sc_hd__xor2_1 _06971_ (.A(reg1_val[7]),
    .B(_06491_),
    .X(_06492_));
 sky130_fd_sc_hd__o21a_1 _06972_ (.A1(reg1_val[7]),
    .A2(_06431_),
    .B1(net275),
    .X(_06493_));
 sky130_fd_sc_hd__xnor2_1 _06973_ (.A(reg1_val[8]),
    .B(_06493_),
    .Y(_06494_));
 sky130_fd_sc_hd__or2_1 _06974_ (.A(net190),
    .B(_06494_),
    .X(_06495_));
 sky130_fd_sc_hd__nand2_1 _06975_ (.A(net190),
    .B(_06494_),
    .Y(_06496_));
 sky130_fd_sc_hd__mux2_1 _06976_ (.A0(_06495_),
    .A1(_06496_),
    .S(_06490_),
    .X(_06497_));
 sky130_fd_sc_hd__inv_2 _06977_ (.A(net152),
    .Y(_06498_));
 sky130_fd_sc_hd__nor2_1 _06978_ (.A(_05840_),
    .B(_05911_),
    .Y(_06499_));
 sky130_fd_sc_hd__nand3_4 _06979_ (.A(_06450_),
    .B(net178),
    .C(_06499_),
    .Y(_06500_));
 sky130_fd_sc_hd__or2_2 _06980_ (.A(_05696_),
    .B(_05778_),
    .X(_06501_));
 sky130_fd_sc_hd__o21ai_4 _06981_ (.A1(_06500_),
    .A2(_06501_),
    .B1(net194),
    .Y(_06502_));
 sky130_fd_sc_hd__xnor2_4 _06982_ (.A(_05620_),
    .B(_06502_),
    .Y(_06503_));
 sky130_fd_sc_hd__xnor2_4 _06983_ (.A(_05611_),
    .B(_06502_),
    .Y(_00136_));
 sky130_fd_sc_hd__nand2_2 _06984_ (.A(_06495_),
    .B(_06496_),
    .Y(_00137_));
 sky130_fd_sc_hd__inv_2 _06985_ (.A(net150),
    .Y(_00138_));
 sky130_fd_sc_hd__o31a_1 _06986_ (.A1(_05620_),
    .A2(_06500_),
    .A3(_06501_),
    .B1(net194),
    .X(_00139_));
 sky130_fd_sc_hd__xnor2_1 _06987_ (.A(_05544_),
    .B(_00139_),
    .Y(_00140_));
 sky130_fd_sc_hd__o22a_1 _06988_ (.A1(net152),
    .A2(net77),
    .B1(net150),
    .B2(net75),
    .X(_00141_));
 sky130_fd_sc_hd__xnor2_1 _06989_ (.A(net191),
    .B(_00141_),
    .Y(_00142_));
 sky130_fd_sc_hd__a31o_1 _06990_ (.A1(_06450_),
    .A2(net178),
    .A3(_06499_),
    .B1(_06447_),
    .X(_00143_));
 sky130_fd_sc_hd__nor2_1 _06991_ (.A(_05768_),
    .B(_06447_),
    .Y(_00144_));
 sky130_fd_sc_hd__a22o_1 _06992_ (.A1(_05768_),
    .A2(_00143_),
    .B1(_00144_),
    .B2(_06500_),
    .X(_00145_));
 sky130_fd_sc_hd__nand2_1 _06993_ (.A(net275),
    .B(_06432_),
    .Y(_00146_));
 sky130_fd_sc_hd__xor2_1 _06994_ (.A(reg1_val[10]),
    .B(_00146_),
    .X(_00147_));
 sky130_fd_sc_hd__or2_1 _06995_ (.A(net191),
    .B(_00147_),
    .X(_00148_));
 sky130_fd_sc_hd__nand2_1 _06996_ (.A(net191),
    .B(_00147_),
    .Y(_00149_));
 sky130_fd_sc_hd__mux2_1 _06997_ (.A0(_00149_),
    .A1(_00148_),
    .S(net180),
    .X(_00150_));
 sky130_fd_sc_hd__inv_2 _06998_ (.A(net116),
    .Y(_00151_));
 sky130_fd_sc_hd__nand2_2 _06999_ (.A(_00148_),
    .B(_00149_),
    .Y(_00152_));
 sky130_fd_sc_hd__inv_2 _07000_ (.A(net114),
    .Y(_00153_));
 sky130_fd_sc_hd__o21ai_1 _07001_ (.A1(_05778_),
    .A2(_06500_),
    .B1(net194),
    .Y(_00154_));
 sky130_fd_sc_hd__xnor2_1 _07002_ (.A(_05705_),
    .B(_00154_),
    .Y(_00155_));
 sky130_fd_sc_hd__o22a_1 _07003_ (.A1(net120),
    .A2(net116),
    .B1(net114),
    .B2(net72),
    .X(_00156_));
 sky130_fd_sc_hd__xnor2_1 _07004_ (.A(net180),
    .B(_00156_),
    .Y(_00157_));
 sky130_fd_sc_hd__o21a_1 _07005_ (.A1(reg1_val[4]),
    .A2(_06430_),
    .B1(net275),
    .X(_00158_));
 sky130_fd_sc_hd__xnor2_1 _07006_ (.A(reg1_val[5]),
    .B(_00158_),
    .Y(_00159_));
 sky130_fd_sc_hd__o31a_1 _07007_ (.A1(reg1_val[4]),
    .A2(reg1_val[5]),
    .A3(_06430_),
    .B1(net275),
    .X(_00160_));
 sky130_fd_sc_hd__xnor2_1 _07008_ (.A(reg1_val[6]),
    .B(_00160_),
    .Y(_00161_));
 sky130_fd_sc_hd__or2_1 _07009_ (.A(net211),
    .B(_00161_),
    .X(_00162_));
 sky130_fd_sc_hd__nand2_1 _07010_ (.A(net211),
    .B(_00161_),
    .Y(_00163_));
 sky130_fd_sc_hd__mux2_4 _07011_ (.A0(_00163_),
    .A1(_00162_),
    .S(net190),
    .X(_00164_));
 sky130_fd_sc_hd__nand2_1 _07012_ (.A(_05533_),
    .B(_05611_),
    .Y(_00165_));
 sky130_fd_sc_hd__o31a_1 _07013_ (.A1(_06500_),
    .A2(_06501_),
    .A3(_00165_),
    .B1(net193),
    .X(_00166_));
 sky130_fd_sc_hd__xnor2_1 _07014_ (.A(_05458_),
    .B(_00166_),
    .Y(_00167_));
 sky130_fd_sc_hd__nand2_4 _07015_ (.A(_00162_),
    .B(_00163_),
    .Y(_00168_));
 sky130_fd_sc_hd__o41a_1 _07016_ (.A1(_05458_),
    .A2(_06500_),
    .A3(_06501_),
    .A4(_00165_),
    .B1(net194),
    .X(_00169_));
 sky130_fd_sc_hd__xnor2_1 _07017_ (.A(_05382_),
    .B(_00169_),
    .Y(_00170_));
 sky130_fd_sc_hd__o22a_1 _07018_ (.A1(net177),
    .A2(net69),
    .B1(net175),
    .B2(net66),
    .X(_00171_));
 sky130_fd_sc_hd__xnor2_1 _07019_ (.A(net190),
    .B(_00171_),
    .Y(_00172_));
 sky130_fd_sc_hd__nor2_1 _07020_ (.A(_00157_),
    .B(_00172_),
    .Y(_00173_));
 sky130_fd_sc_hd__xor2_1 _07021_ (.A(_00157_),
    .B(_00172_),
    .X(_00174_));
 sky130_fd_sc_hd__and2b_1 _07022_ (.A_N(_00142_),
    .B(_00174_),
    .X(_00175_));
 sky130_fd_sc_hd__xnor2_1 _07023_ (.A(_00142_),
    .B(_00174_),
    .Y(_00176_));
 sky130_fd_sc_hd__nand2_1 _07024_ (.A(_06487_),
    .B(_00176_),
    .Y(_00177_));
 sky130_fd_sc_hd__o31a_2 _07025_ (.A1(reg1_val[0]),
    .A2(reg1_val[1]),
    .A3(reg1_val[2]),
    .B1(net274),
    .X(_00178_));
 sky130_fd_sc_hd__xnor2_4 _07026_ (.A(reg1_val[3]),
    .B(_00178_),
    .Y(_00179_));
 sky130_fd_sc_hd__clkinv_8 _07027_ (.A(net208),
    .Y(_00180_));
 sky130_fd_sc_hd__or4_4 _07028_ (.A(_05382_),
    .B(_05458_),
    .C(_06501_),
    .D(_00165_),
    .X(_00181_));
 sky130_fd_sc_hd__nand2_1 _07029_ (.A(_04980_),
    .B(_05111_),
    .Y(_00182_));
 sky130_fd_sc_hd__o31a_1 _07030_ (.A1(_06500_),
    .A2(_00181_),
    .A3(_00182_),
    .B1(net194),
    .X(_00183_));
 sky130_fd_sc_hd__o31a_1 _07031_ (.A1(_06500_),
    .A2(_00181_),
    .A3(_00182_),
    .B1(_04828_),
    .X(_00184_));
 sky130_fd_sc_hd__a2bb2o_4 _07032_ (.A1_N(_04828_),
    .A2_N(_00183_),
    .B1(_00184_),
    .B2(net194),
    .X(_00185_));
 sky130_fd_sc_hd__and3_4 _07033_ (.A(net304),
    .B(reg1_val[31]),
    .C(net307),
    .X(_00186_));
 sky130_fd_sc_hd__xnor2_4 _07034_ (.A(_04438_),
    .B(_00186_),
    .Y(_00187_));
 sky130_fd_sc_hd__xnor2_4 _07035_ (.A(reg1_val[1]),
    .B(_00186_),
    .Y(_00188_));
 sky130_fd_sc_hd__o21a_1 _07036_ (.A1(net304),
    .A2(reg1_val[1]),
    .B1(net275),
    .X(_00189_));
 sky130_fd_sc_hd__xnor2_2 _07037_ (.A(reg1_val[2]),
    .B(_00189_),
    .Y(_00190_));
 sky130_fd_sc_hd__or2_1 _07038_ (.A(net255),
    .B(_00190_),
    .X(_00191_));
 sky130_fd_sc_hd__nand2_1 _07039_ (.A(net255),
    .B(_00190_),
    .Y(_00192_));
 sky130_fd_sc_hd__mux2_2 _07040_ (.A0(_00191_),
    .A1(_00192_),
    .S(_00180_),
    .X(_00193_));
 sky130_fd_sc_hd__nand2_2 _07041_ (.A(_00191_),
    .B(_00192_),
    .Y(_00194_));
 sky130_fd_sc_hd__o41a_4 _07042_ (.A1(_04828_),
    .A2(_06500_),
    .A3(_00181_),
    .A4(_00182_),
    .B1(net194),
    .X(_00195_));
 sky130_fd_sc_hd__xnor2_2 _07043_ (.A(_04894_),
    .B(_00195_),
    .Y(_00196_));
 sky130_fd_sc_hd__xnor2_4 _07044_ (.A(_04904_),
    .B(_00195_),
    .Y(_00197_));
 sky130_fd_sc_hd__o22a_1 _07045_ (.A1(_00185_),
    .A2(net173),
    .B1(net171),
    .B2(net61),
    .X(_00198_));
 sky130_fd_sc_hd__xnor2_2 _07046_ (.A(net208),
    .B(_00198_),
    .Y(_00199_));
 sky130_fd_sc_hd__o21ai_1 _07047_ (.A1(_06500_),
    .A2(_00181_),
    .B1(net194),
    .Y(_00200_));
 sky130_fd_sc_hd__o211a_1 _07048_ (.A1(_06500_),
    .A2(_00181_),
    .B1(_05122_),
    .C1(net194),
    .X(_00201_));
 sky130_fd_sc_hd__a21o_1 _07049_ (.A1(_05111_),
    .A2(_00200_),
    .B1(_00201_),
    .X(_00202_));
 sky130_fd_sc_hd__nand2_1 _07050_ (.A(net275),
    .B(_06430_),
    .Y(_00203_));
 sky130_fd_sc_hd__xnor2_2 _07051_ (.A(_04449_),
    .B(_00203_),
    .Y(_00204_));
 sky130_fd_sc_hd__or2_1 _07052_ (.A(net208),
    .B(_00204_),
    .X(_00205_));
 sky130_fd_sc_hd__nand2_1 _07053_ (.A(net208),
    .B(_00204_),
    .Y(_00206_));
 sky130_fd_sc_hd__mux2_1 _07054_ (.A0(_00206_),
    .A1(_00205_),
    .S(net211),
    .X(_00207_));
 sky130_fd_sc_hd__inv_2 _07055_ (.A(net169),
    .Y(_00208_));
 sky130_fd_sc_hd__nand2_2 _07056_ (.A(_00205_),
    .B(_00206_),
    .Y(_00209_));
 sky130_fd_sc_hd__inv_2 _07057_ (.A(net167),
    .Y(_00210_));
 sky130_fd_sc_hd__o31a_1 _07058_ (.A1(_05122_),
    .A2(_06500_),
    .A3(_00181_),
    .B1(net194),
    .X(_00211_));
 sky130_fd_sc_hd__xor2_1 _07059_ (.A(_04980_),
    .B(_00211_),
    .X(_00212_));
 sky130_fd_sc_hd__o22a_1 _07060_ (.A1(net59),
    .A2(net169),
    .B1(net167),
    .B2(net56),
    .X(_00213_));
 sky130_fd_sc_hd__xor2_1 _07061_ (.A(net210),
    .B(_00213_),
    .X(_00214_));
 sky130_fd_sc_hd__nor2_2 _07062_ (.A(net304),
    .B(_04438_),
    .Y(_00215_));
 sky130_fd_sc_hd__nand2_1 _07063_ (.A(net301),
    .B(reg1_val[1]),
    .Y(_00216_));
 sky130_fd_sc_hd__or2_1 _07064_ (.A(_04828_),
    .B(_04894_),
    .X(_00217_));
 sky130_fd_sc_hd__or4_4 _07065_ (.A(_06500_),
    .B(_00181_),
    .C(_00182_),
    .D(_00217_),
    .X(_00218_));
 sky130_fd_sc_hd__a21o_4 _07066_ (.A1(net193),
    .A2(_00218_),
    .B1(_05263_),
    .X(_00219_));
 sky130_fd_sc_hd__nor2_2 _07067_ (.A(_05274_),
    .B(_06447_),
    .Y(_00220_));
 sky130_fd_sc_hd__nand2_8 _07068_ (.A(_00218_),
    .B(_00220_),
    .Y(_00221_));
 sky130_fd_sc_hd__and2_2 _07069_ (.A(_00219_),
    .B(_00221_),
    .X(_00222_));
 sky130_fd_sc_hd__nand2_4 _07070_ (.A(_00219_),
    .B(_00221_),
    .Y(_00223_));
 sky130_fd_sc_hd__and3_1 _07071_ (.A(_00215_),
    .B(_00219_),
    .C(_00221_),
    .X(_00224_));
 sky130_fd_sc_hd__o211ai_4 _07072_ (.A1(_05263_),
    .A2(_00218_),
    .B1(net193),
    .C1(_05187_),
    .Y(_00225_));
 sky130_fd_sc_hd__a211o_4 _07073_ (.A1(net193),
    .A2(_00218_),
    .B1(_00220_),
    .C1(_05187_),
    .X(_00226_));
 sky130_fd_sc_hd__and2_1 _07074_ (.A(_00225_),
    .B(_00226_),
    .X(_00227_));
 sky130_fd_sc_hd__nand2_2 _07075_ (.A(_00225_),
    .B(_00226_),
    .Y(_00228_));
 sky130_fd_sc_hd__a21oi_1 _07076_ (.A1(_00225_),
    .A2(_00226_),
    .B1(net302),
    .Y(_00229_));
 sky130_fd_sc_hd__o21ai_1 _07077_ (.A1(_00224_),
    .A2(_00229_),
    .B1(_00187_),
    .Y(_00230_));
 sky130_fd_sc_hd__or3_1 _07078_ (.A(_00187_),
    .B(_00224_),
    .C(_00229_),
    .X(_00231_));
 sky130_fd_sc_hd__and3_1 _07079_ (.A(_00214_),
    .B(_00230_),
    .C(_00231_),
    .X(_00232_));
 sky130_fd_sc_hd__a21oi_1 _07080_ (.A1(_00230_),
    .A2(_00231_),
    .B1(_00214_),
    .Y(_00233_));
 sky130_fd_sc_hd__or2_1 _07081_ (.A(_00232_),
    .B(_00233_),
    .X(_00234_));
 sky130_fd_sc_hd__xnor2_2 _07082_ (.A(_00199_),
    .B(_00234_),
    .Y(_00235_));
 sky130_fd_sc_hd__xnor2_1 _07083_ (.A(_06487_),
    .B(_00176_),
    .Y(_00236_));
 sky130_fd_sc_hd__o21ai_1 _07084_ (.A1(_00235_),
    .A2(_00236_),
    .B1(_00177_),
    .Y(_00237_));
 sky130_fd_sc_hd__or2_2 _07085_ (.A(reg1_val[14]),
    .B(reg1_val[15]),
    .X(_00238_));
 sky130_fd_sc_hd__or2_1 _07086_ (.A(reg1_val[16]),
    .B(reg1_val[17]),
    .X(_00239_));
 sky130_fd_sc_hd__or2_1 _07087_ (.A(reg1_val[18]),
    .B(_00239_),
    .X(_00240_));
 sky130_fd_sc_hd__or2_1 _07088_ (.A(reg1_val[19]),
    .B(_00240_),
    .X(_00241_));
 sky130_fd_sc_hd__or2_1 _07089_ (.A(reg1_val[20]),
    .B(reg1_val[21]),
    .X(_00242_));
 sky130_fd_sc_hd__or4_2 _07090_ (.A(reg1_val[22]),
    .B(reg1_val[23]),
    .C(_00241_),
    .D(_00242_),
    .X(_00243_));
 sky130_fd_sc_hd__or4_4 _07091_ (.A(net303),
    .B(_06433_),
    .C(_00238_),
    .D(_00243_),
    .X(_00244_));
 sky130_fd_sc_hd__or2_2 _07092_ (.A(reg1_val[24]),
    .B(reg1_val[25]),
    .X(_00245_));
 sky130_fd_sc_hd__o21a_4 _07093_ (.A1(_00244_),
    .A2(_00245_),
    .B1(net274),
    .X(_00246_));
 sky130_fd_sc_hd__o31a_2 _07094_ (.A1(reg1_val[26]),
    .A2(_00244_),
    .A3(_00245_),
    .B1(net274),
    .X(_00247_));
 sky130_fd_sc_hd__xor2_4 _07095_ (.A(reg1_val[27]),
    .B(_00247_),
    .X(_00248_));
 sky130_fd_sc_hd__o211a_1 _07096_ (.A1(_06299_),
    .A2(net227),
    .B1(net307),
    .C1(_04752_),
    .X(_00249_));
 sky130_fd_sc_hd__o311a_2 _07097_ (.A1(net233),
    .A2(_06299_),
    .A3(net227),
    .B1(_04752_),
    .C1(net307),
    .X(_00250_));
 sky130_fd_sc_hd__xnor2_2 _07098_ (.A(_06287_),
    .B(_00250_),
    .Y(_00251_));
 sky130_fd_sc_hd__xor2_2 _07099_ (.A(_06287_),
    .B(_00250_),
    .X(_00252_));
 sky130_fd_sc_hd__o41a_2 _07100_ (.A1(net303),
    .A2(_06433_),
    .A3(_00238_),
    .A4(_00243_),
    .B1(net274),
    .X(_00253_));
 sky130_fd_sc_hd__o21ai_2 _07101_ (.A1(reg1_val[24]),
    .A2(_00244_),
    .B1(net274),
    .Y(_00254_));
 sky130_fd_sc_hd__xnor2_4 _07102_ (.A(reg1_val[25]),
    .B(_00254_),
    .Y(_00255_));
 sky130_fd_sc_hd__xnor2_4 _07103_ (.A(_04482_),
    .B(_00246_),
    .Y(_00256_));
 sky130_fd_sc_hd__nand3b_1 _07104_ (.A_N(net113),
    .B(net110),
    .C(_00256_),
    .Y(_00257_));
 sky130_fd_sc_hd__or3b_1 _07105_ (.A(net110),
    .B(_00256_),
    .C_N(net113),
    .X(_00258_));
 sky130_fd_sc_hd__and2_1 _07106_ (.A(_00257_),
    .B(_00258_),
    .X(_00259_));
 sky130_fd_sc_hd__a21oi_2 _07107_ (.A1(net193),
    .A2(_06448_),
    .B1(net240),
    .Y(_00260_));
 sky130_fd_sc_hd__and3_1 _07108_ (.A(net307),
    .B(_04752_),
    .C(net240),
    .X(_00261_));
 sky130_fd_sc_hd__and2_1 _07109_ (.A(_06448_),
    .B(_00261_),
    .X(_00262_));
 sky130_fd_sc_hd__nor2_2 _07110_ (.A(_00260_),
    .B(_00262_),
    .Y(_00263_));
 sky130_fd_sc_hd__or2_1 _07111_ (.A(_00260_),
    .B(_00262_),
    .X(_00264_));
 sky130_fd_sc_hd__xnor2_4 _07112_ (.A(net110),
    .B(_00256_),
    .Y(_00265_));
 sky130_fd_sc_hd__o22a_1 _07113_ (.A1(net165),
    .A2(net15),
    .B1(net149),
    .B2(net53),
    .X(_00266_));
 sky130_fd_sc_hd__xnor2_1 _07114_ (.A(net113),
    .B(_00266_),
    .Y(_00267_));
 sky130_fd_sc_hd__o41a_4 _07115_ (.A1(net303),
    .A2(_06433_),
    .A3(_00238_),
    .A4(_00241_),
    .B1(net274),
    .X(_00268_));
 sky130_fd_sc_hd__o21a_1 _07116_ (.A1(reg1_val[22]),
    .A2(_00242_),
    .B1(net274),
    .X(_00269_));
 sky130_fd_sc_hd__o21ai_2 _07117_ (.A1(_00268_),
    .A2(_00269_),
    .B1(reg1_val[23]),
    .Y(_00270_));
 sky130_fd_sc_hd__or3_2 _07118_ (.A(reg1_val[23]),
    .B(_00268_),
    .C(_00269_),
    .X(_00271_));
 sky130_fd_sc_hd__and2_1 _07119_ (.A(_00270_),
    .B(_00271_),
    .X(_00272_));
 sky130_fd_sc_hd__o31a_2 _07120_ (.A1(_06273_),
    .A2(net240),
    .A3(_06448_),
    .B1(net193),
    .X(_00273_));
 sky130_fd_sc_hd__o41ai_4 _07121_ (.A1(_06265_),
    .A2(_06273_),
    .A3(net240),
    .A4(_06448_),
    .B1(net193),
    .Y(_00274_));
 sky130_fd_sc_hd__xor2_4 _07122_ (.A(_06258_),
    .B(_00274_),
    .X(_00275_));
 sky130_fd_sc_hd__xnor2_2 _07123_ (.A(_06258_),
    .B(_00274_),
    .Y(_00276_));
 sky130_fd_sc_hd__and3_1 _07124_ (.A(reg1_val[20]),
    .B(reg1_val[31]),
    .C(net307),
    .X(_00277_));
 sky130_fd_sc_hd__o21a_1 _07125_ (.A1(_00268_),
    .A2(_00277_),
    .B1(reg1_val[21]),
    .X(_00278_));
 sky130_fd_sc_hd__nor3_1 _07126_ (.A(reg1_val[21]),
    .B(_00268_),
    .C(_00277_),
    .Y(_00279_));
 sky130_fd_sc_hd__nor2_1 _07127_ (.A(_00278_),
    .B(_00279_),
    .Y(_00280_));
 sky130_fd_sc_hd__and2_1 _07128_ (.A(net274),
    .B(_00242_),
    .X(_00281_));
 sky130_fd_sc_hd__o21a_1 _07129_ (.A1(_00268_),
    .A2(_00281_),
    .B1(reg1_val[22]),
    .X(_00282_));
 sky130_fd_sc_hd__nor3_1 _07130_ (.A(reg1_val[22]),
    .B(_00268_),
    .C(_00281_),
    .Y(_00283_));
 sky130_fd_sc_hd__nor2_2 _07131_ (.A(_00282_),
    .B(_00283_),
    .Y(_00284_));
 sky130_fd_sc_hd__or4_2 _07132_ (.A(_00278_),
    .B(_00279_),
    .C(_00282_),
    .D(_00283_),
    .X(_00285_));
 sky130_fd_sc_hd__nor2_1 _07133_ (.A(net106),
    .B(_00285_),
    .Y(_00286_));
 sky130_fd_sc_hd__o22ai_2 _07134_ (.A1(_00278_),
    .A2(_00279_),
    .B1(_00282_),
    .B2(_00283_),
    .Y(_00287_));
 sky130_fd_sc_hd__mux2_1 _07135_ (.A0(_00285_),
    .A1(_00287_),
    .S(net106),
    .X(_00288_));
 sky130_fd_sc_hd__o21a_1 _07136_ (.A1(_06448_),
    .A2(_06449_),
    .B1(net193),
    .X(_00289_));
 sky130_fd_sc_hd__xnor2_4 _07137_ (.A(_06252_),
    .B(_00289_),
    .Y(_00290_));
 sky130_fd_sc_hd__nand2_2 _07138_ (.A(_00285_),
    .B(_00287_),
    .Y(_00291_));
 sky130_fd_sc_hd__o22a_1 _07139_ (.A1(net147),
    .A2(net51),
    .B1(net144),
    .B2(net49),
    .X(_00292_));
 sky130_fd_sc_hd__xnor2_1 _07140_ (.A(net107),
    .B(_00292_),
    .Y(_00293_));
 sky130_fd_sc_hd__and2_1 _07141_ (.A(_00267_),
    .B(_00293_),
    .X(_00294_));
 sky130_fd_sc_hd__nor2_1 _07142_ (.A(_00267_),
    .B(_00293_),
    .Y(_00295_));
 sky130_fd_sc_hd__or2_1 _07143_ (.A(_00294_),
    .B(_00295_),
    .X(_00296_));
 sky130_fd_sc_hd__o211ai_2 _07144_ (.A1(net240),
    .A2(_06448_),
    .B1(net193),
    .C1(_06272_),
    .Y(_00297_));
 sky130_fd_sc_hd__a211o_1 _07145_ (.A1(net193),
    .A2(_06448_),
    .B1(_00261_),
    .C1(_06272_),
    .X(_00298_));
 sky130_fd_sc_hd__and2_1 _07146_ (.A(_00297_),
    .B(_00298_),
    .X(_00299_));
 sky130_fd_sc_hd__nand2_2 _07147_ (.A(_00297_),
    .B(_00298_),
    .Y(_00300_));
 sky130_fd_sc_hd__xor2_4 _07148_ (.A(reg1_val[24]),
    .B(_00253_),
    .X(_00301_));
 sky130_fd_sc_hd__and3_2 _07149_ (.A(_00270_),
    .B(_00271_),
    .C(_00301_),
    .X(_00302_));
 sky130_fd_sc_hd__nand2_1 _07150_ (.A(net107),
    .B(_00301_),
    .Y(_00303_));
 sky130_fd_sc_hd__a21oi_4 _07151_ (.A1(_00270_),
    .A2(_00271_),
    .B1(_00301_),
    .Y(_00304_));
 sky130_fd_sc_hd__or2_1 _07152_ (.A(net107),
    .B(_00301_),
    .X(_00305_));
 sky130_fd_sc_hd__mux2_2 _07153_ (.A0(_00303_),
    .A1(_00305_),
    .S(net109),
    .X(_00306_));
 sky130_fd_sc_hd__mux2_8 _07154_ (.A0(_00302_),
    .A1(_00304_),
    .S(net108),
    .X(_00307_));
 sky130_fd_sc_hd__nor2_8 _07155_ (.A(_00302_),
    .B(_00304_),
    .Y(_00308_));
 sky130_fd_sc_hd__or2_4 _07156_ (.A(_00302_),
    .B(_00304_),
    .X(_00309_));
 sky130_fd_sc_hd__xor2_4 _07157_ (.A(_06265_),
    .B(_00273_),
    .X(_00310_));
 sky130_fd_sc_hd__xnor2_2 _07158_ (.A(_06265_),
    .B(_00273_),
    .Y(_00311_));
 sky130_fd_sc_hd__a22o_1 _07159_ (.A1(_00300_),
    .A2(_00307_),
    .B1(_00308_),
    .B2(_00310_),
    .X(_00312_));
 sky130_fd_sc_hd__xnor2_1 _07160_ (.A(net110),
    .B(_00312_),
    .Y(_00313_));
 sky130_fd_sc_hd__nor2_1 _07161_ (.A(_00296_),
    .B(_00313_),
    .Y(_00314_));
 sky130_fd_sc_hd__and2_1 _07162_ (.A(_00296_),
    .B(_00313_),
    .X(_00315_));
 sky130_fd_sc_hd__nor2_1 _07163_ (.A(_00314_),
    .B(_00315_),
    .Y(_00316_));
 sky130_fd_sc_hd__a31o_1 _07164_ (.A1(_05922_),
    .A2(_06450_),
    .A3(_06463_),
    .B1(_06447_),
    .X(_00317_));
 sky130_fd_sc_hd__xnor2_2 _07165_ (.A(_05850_),
    .B(_00317_),
    .Y(_00318_));
 sky130_fd_sc_hd__o22a_1 _07166_ (.A1(net120),
    .A2(net114),
    .B1(net101),
    .B2(net116),
    .X(_00319_));
 sky130_fd_sc_hd__xnor2_1 _07167_ (.A(net180),
    .B(_00319_),
    .Y(_00320_));
 sky130_fd_sc_hd__o22a_1 _07168_ (.A1(net75),
    .A2(net177),
    .B1(net69),
    .B2(net175),
    .X(_00321_));
 sky130_fd_sc_hd__xnor2_1 _07169_ (.A(net190),
    .B(_00321_),
    .Y(_00322_));
 sky130_fd_sc_hd__nor2_1 _07170_ (.A(_00320_),
    .B(_00322_),
    .Y(_00323_));
 sky130_fd_sc_hd__o22a_1 _07171_ (.A1(net77),
    .A2(net150),
    .B1(net72),
    .B2(net152),
    .X(_00324_));
 sky130_fd_sc_hd__xnor2_2 _07172_ (.A(net191),
    .B(_00324_),
    .Y(_00325_));
 sky130_fd_sc_hd__inv_2 _07173_ (.A(_00325_),
    .Y(_00326_));
 sky130_fd_sc_hd__xor2_1 _07174_ (.A(_00320_),
    .B(_00322_),
    .X(_00327_));
 sky130_fd_sc_hd__a21oi_1 _07175_ (.A1(_00326_),
    .A2(_00327_),
    .B1(_00323_),
    .Y(_00328_));
 sky130_fd_sc_hd__or3_4 _07176_ (.A(reg1_val[26]),
    .B(reg1_val[27]),
    .C(_00245_),
    .X(_00329_));
 sky130_fd_sc_hd__o31a_1 _07177_ (.A1(reg1_val[28]),
    .A2(_00244_),
    .A3(_00329_),
    .B1(net274),
    .X(_00330_));
 sky130_fd_sc_hd__xnor2_2 _07178_ (.A(reg1_val[29]),
    .B(_00330_),
    .Y(_00331_));
 sky130_fd_sc_hd__o21ai_2 _07179_ (.A1(_00244_),
    .A2(_00329_),
    .B1(net274),
    .Y(_00332_));
 sky130_fd_sc_hd__xnor2_4 _07180_ (.A(reg1_val[28]),
    .B(_00332_),
    .Y(_00333_));
 sky130_fd_sc_hd__o21ba_1 _07181_ (.A1(net112),
    .A2(_00333_),
    .B1_N(net97),
    .X(_00334_));
 sky130_fd_sc_hd__a21boi_1 _07182_ (.A1(net112),
    .A2(_00333_),
    .B1_N(net97),
    .Y(_00335_));
 sky130_fd_sc_hd__or2_1 _07183_ (.A(_00334_),
    .B(_00335_),
    .X(_00336_));
 sky130_fd_sc_hd__and3_2 _07184_ (.A(net307),
    .B(_04752_),
    .C(net227),
    .X(_00337_));
 sky130_fd_sc_hd__xnor2_4 _07185_ (.A(net229),
    .B(_00337_),
    .Y(_00338_));
 sky130_fd_sc_hd__xnor2_2 _07186_ (.A(_06299_),
    .B(_00337_),
    .Y(_00339_));
 sky130_fd_sc_hd__xnor2_1 _07187_ (.A(net113),
    .B(_00333_),
    .Y(_00340_));
 sky130_fd_sc_hd__o22a_1 _07188_ (.A1(net226),
    .A2(net12),
    .B1(net163),
    .B2(net46),
    .X(_00341_));
 sky130_fd_sc_hd__xor2_2 _07189_ (.A(net98),
    .B(_00341_),
    .X(_00342_));
 sky130_fd_sc_hd__and2b_1 _07190_ (.A_N(_00328_),
    .B(_00342_),
    .X(_00343_));
 sky130_fd_sc_hd__o22a_1 _07191_ (.A1(net66),
    .A2(net169),
    .B1(net167),
    .B2(net59),
    .X(_00344_));
 sky130_fd_sc_hd__xnor2_1 _07192_ (.A(net210),
    .B(_00344_),
    .Y(_00345_));
 sky130_fd_sc_hd__a22o_1 _07193_ (.A1(_00197_),
    .A2(_00215_),
    .B1(_00222_),
    .B2(net304),
    .X(_00346_));
 sky130_fd_sc_hd__xnor2_2 _07194_ (.A(_00187_),
    .B(_00346_),
    .Y(_00347_));
 sky130_fd_sc_hd__nor2_1 _07195_ (.A(_00345_),
    .B(_00347_),
    .Y(_00348_));
 sky130_fd_sc_hd__o22a_1 _07196_ (.A1(_00185_),
    .A2(net171),
    .B1(net56),
    .B2(net173),
    .X(_00349_));
 sky130_fd_sc_hd__xnor2_1 _07197_ (.A(net208),
    .B(_00349_),
    .Y(_00350_));
 sky130_fd_sc_hd__xor2_1 _07198_ (.A(_00345_),
    .B(_00347_),
    .X(_00351_));
 sky130_fd_sc_hd__and2b_1 _07199_ (.A_N(_00350_),
    .B(_00351_),
    .X(_00352_));
 sky130_fd_sc_hd__xnor2_1 _07200_ (.A(_00328_),
    .B(_00342_),
    .Y(_00353_));
 sky130_fd_sc_hd__o21a_1 _07201_ (.A1(_00348_),
    .A2(_00352_),
    .B1(_00353_),
    .X(_00354_));
 sky130_fd_sc_hd__or2_1 _07202_ (.A(_00343_),
    .B(_00354_),
    .X(_00355_));
 sky130_fd_sc_hd__xnor2_1 _07203_ (.A(_00316_),
    .B(_00355_),
    .Y(_00356_));
 sky130_fd_sc_hd__and2b_1 _07204_ (.A_N(_00356_),
    .B(_00237_),
    .X(_00357_));
 sky130_fd_sc_hd__and2b_1 _07205_ (.A_N(_00237_),
    .B(_00356_),
    .X(_00358_));
 sky130_fd_sc_hd__nor2_1 _07206_ (.A(_00357_),
    .B(_00358_),
    .Y(_00359_));
 sky130_fd_sc_hd__o22a_1 _07207_ (.A1(net82),
    .A2(net128),
    .B1(net101),
    .B2(net130),
    .X(_00360_));
 sky130_fd_sc_hd__xnor2_2 _07208_ (.A(net158),
    .B(_00360_),
    .Y(_00361_));
 sky130_fd_sc_hd__o22a_1 _07209_ (.A1(net80),
    .A2(net124),
    .B1(net121),
    .B2(net79),
    .X(_00362_));
 sky130_fd_sc_hd__xnor2_2 _07210_ (.A(net155),
    .B(_00362_),
    .Y(_00363_));
 sky130_fd_sc_hd__and2b_1 _07211_ (.A_N(_00361_),
    .B(_00363_),
    .X(_00364_));
 sky130_fd_sc_hd__o21ba_1 _07212_ (.A1(_00199_),
    .A2(_00233_),
    .B1_N(_00232_),
    .X(_00365_));
 sky130_fd_sc_hd__and2b_1 _07213_ (.A_N(_00365_),
    .B(_00364_),
    .X(_00366_));
 sky130_fd_sc_hd__xnor2_1 _07214_ (.A(_00364_),
    .B(_00365_),
    .Y(_00367_));
 sky130_fd_sc_hd__o21a_1 _07215_ (.A1(_00173_),
    .A2(_00175_),
    .B1(_00367_),
    .X(_00368_));
 sky130_fd_sc_hd__nor3_1 _07216_ (.A(_00173_),
    .B(_00175_),
    .C(_00367_),
    .Y(_00369_));
 sky130_fd_sc_hd__or2_1 _07217_ (.A(_00368_),
    .B(_00369_),
    .X(_00370_));
 sky130_fd_sc_hd__o22a_1 _07218_ (.A1(net152),
    .A2(net75),
    .B1(net69),
    .B2(net150),
    .X(_00371_));
 sky130_fd_sc_hd__xnor2_2 _07219_ (.A(net191),
    .B(_00371_),
    .Y(_00372_));
 sky130_fd_sc_hd__o22a_1 _07220_ (.A1(net177),
    .A2(net66),
    .B1(net59),
    .B2(net175),
    .X(_00373_));
 sky130_fd_sc_hd__xnor2_2 _07221_ (.A(net190),
    .B(_00373_),
    .Y(_00374_));
 sky130_fd_sc_hd__o22a_1 _07222_ (.A1(net77),
    .A2(net114),
    .B1(net72),
    .B2(net116),
    .X(_00375_));
 sky130_fd_sc_hd__xnor2_2 _07223_ (.A(net180),
    .B(_00375_),
    .Y(_00376_));
 sky130_fd_sc_hd__nor2_1 _07224_ (.A(_00374_),
    .B(_00376_),
    .Y(_00377_));
 sky130_fd_sc_hd__xor2_2 _07225_ (.A(_00374_),
    .B(_00376_),
    .X(_00378_));
 sky130_fd_sc_hd__and2b_1 _07226_ (.A_N(_00372_),
    .B(_00378_),
    .X(_00379_));
 sky130_fd_sc_hd__xnor2_2 _07227_ (.A(_00372_),
    .B(_00378_),
    .Y(_00380_));
 sky130_fd_sc_hd__o22a_1 _07228_ (.A1(net131),
    .A2(net120),
    .B1(net101),
    .B2(net82),
    .X(_00381_));
 sky130_fd_sc_hd__xnor2_1 _07229_ (.A(net158),
    .B(_00381_),
    .Y(_00382_));
 sky130_fd_sc_hd__o31a_2 _07230_ (.A1(net303),
    .A2(_06433_),
    .A3(_00238_),
    .B1(net275),
    .X(_00383_));
 sky130_fd_sc_hd__o41a_1 _07231_ (.A1(reg1_val[13]),
    .A2(reg1_val[16]),
    .A3(_06433_),
    .A4(_00238_),
    .B1(net275),
    .X(_00384_));
 sky130_fd_sc_hd__xor2_1 _07232_ (.A(reg1_val[17]),
    .B(_00384_),
    .X(_00385_));
 sky130_fd_sc_hd__xnor2_4 _07233_ (.A(_04460_),
    .B(_00383_),
    .Y(_00386_));
 sky130_fd_sc_hd__nand3b_1 _07234_ (.A_N(net137),
    .B(_00386_),
    .C(net154),
    .Y(_00387_));
 sky130_fd_sc_hd__or3b_1 _07235_ (.A(net154),
    .B(_00386_),
    .C_N(net137),
    .X(_00388_));
 sky130_fd_sc_hd__and2_1 _07236_ (.A(_00387_),
    .B(_00388_),
    .X(_00389_));
 sky130_fd_sc_hd__nand2_1 _07237_ (.A(_00387_),
    .B(_00388_),
    .Y(_00390_));
 sky130_fd_sc_hd__xnor2_4 _07238_ (.A(net155),
    .B(_00386_),
    .Y(_00391_));
 sky130_fd_sc_hd__inv_2 _07239_ (.A(net94),
    .Y(_00392_));
 sky130_fd_sc_hd__o22a_1 _07240_ (.A1(net127),
    .A2(net42),
    .B1(net94),
    .B2(net121),
    .X(_00393_));
 sky130_fd_sc_hd__xor2_1 _07241_ (.A(net138),
    .B(_00393_),
    .X(_00394_));
 sky130_fd_sc_hd__nor2_1 _07242_ (.A(_00382_),
    .B(_00394_),
    .Y(_00395_));
 sky130_fd_sc_hd__xnor2_1 _07243_ (.A(_00382_),
    .B(_00394_),
    .Y(_00396_));
 sky130_fd_sc_hd__o22a_1 _07244_ (.A1(net80),
    .A2(net78),
    .B1(net124),
    .B2(net128),
    .X(_00397_));
 sky130_fd_sc_hd__xor2_1 _07245_ (.A(net155),
    .B(_00397_),
    .X(_00398_));
 sky130_fd_sc_hd__nor2_1 _07246_ (.A(_00396_),
    .B(_00398_),
    .Y(_00399_));
 sky130_fd_sc_hd__or2_1 _07247_ (.A(_00396_),
    .B(_00398_),
    .X(_00400_));
 sky130_fd_sc_hd__nand2_1 _07248_ (.A(_00396_),
    .B(_00398_),
    .Y(_00401_));
 sky130_fd_sc_hd__nand2_1 _07249_ (.A(_00400_),
    .B(_00401_),
    .Y(_00402_));
 sky130_fd_sc_hd__o22ai_4 _07250_ (.A1(net173),
    .A2(net61),
    .B1(net18),
    .B2(net171),
    .Y(_00403_));
 sky130_fd_sc_hd__xnor2_4 _07251_ (.A(net208),
    .B(_00403_),
    .Y(_00404_));
 sky130_fd_sc_hd__o22a_2 _07252_ (.A1(net62),
    .A2(net167),
    .B1(net54),
    .B2(net169),
    .X(_00405_));
 sky130_fd_sc_hd__xnor2_4 _07253_ (.A(net210),
    .B(_00405_),
    .Y(_00406_));
 sky130_fd_sc_hd__o31a_2 _07254_ (.A1(_05198_),
    .A2(_05263_),
    .A3(_00218_),
    .B1(net193),
    .X(_00407_));
 sky130_fd_sc_hd__xnor2_4 _07255_ (.A(_05046_),
    .B(_00407_),
    .Y(_00408_));
 sky130_fd_sc_hd__o22a_2 _07256_ (.A1(net253),
    .A2(net16),
    .B1(net10),
    .B2(net302),
    .X(_00409_));
 sky130_fd_sc_hd__xnor2_4 _07257_ (.A(net255),
    .B(_00409_),
    .Y(_00410_));
 sky130_fd_sc_hd__nor2_1 _07258_ (.A(_00406_),
    .B(_00410_),
    .Y(_00411_));
 sky130_fd_sc_hd__xor2_4 _07259_ (.A(_00406_),
    .B(_00410_),
    .X(_00412_));
 sky130_fd_sc_hd__xor2_4 _07260_ (.A(_00404_),
    .B(_00412_),
    .X(_00413_));
 sky130_fd_sc_hd__xnor2_2 _07261_ (.A(_00402_),
    .B(_00413_),
    .Y(_00414_));
 sky130_fd_sc_hd__xnor2_1 _07262_ (.A(_00380_),
    .B(_00414_),
    .Y(_00415_));
 sky130_fd_sc_hd__or4_1 _07263_ (.A(reg1_val[28]),
    .B(reg1_val[29]),
    .C(_00244_),
    .D(_00329_),
    .X(_00416_));
 sky130_fd_sc_hd__o41a_2 _07264_ (.A1(reg1_val[28]),
    .A2(reg1_val[29]),
    .A3(_00244_),
    .A4(_00329_),
    .B1(net274),
    .X(_00417_));
 sky130_fd_sc_hd__xnor2_4 _07265_ (.A(reg1_val[30]),
    .B(_00417_),
    .Y(_00418_));
 sky130_fd_sc_hd__or2_1 _07266_ (.A(net98),
    .B(_00418_),
    .X(_00419_));
 sky130_fd_sc_hd__nand2_1 _07267_ (.A(net98),
    .B(_00418_),
    .Y(_00420_));
 sky130_fd_sc_hd__nand2_2 _07268_ (.A(_00419_),
    .B(_00420_),
    .Y(_00421_));
 sky130_fd_sc_hd__or2_1 _07269_ (.A(net226),
    .B(net8),
    .X(_00422_));
 sky130_fd_sc_hd__xnor2_1 _07270_ (.A(net233),
    .B(_00249_),
    .Y(_00423_));
 sky130_fd_sc_hd__xor2_2 _07271_ (.A(net233),
    .B(_00249_),
    .X(_00424_));
 sky130_fd_sc_hd__o22a_1 _07272_ (.A1(net12),
    .A2(net163),
    .B1(net46),
    .B2(net161),
    .X(_00425_));
 sky130_fd_sc_hd__xnor2_1 _07273_ (.A(net98),
    .B(_00425_),
    .Y(_00426_));
 sky130_fd_sc_hd__xnor2_1 _07274_ (.A(_00422_),
    .B(_00426_),
    .Y(_00427_));
 sky130_fd_sc_hd__xnor2_1 _07275_ (.A(_00415_),
    .B(_00427_),
    .Y(_00428_));
 sky130_fd_sc_hd__xor2_1 _07276_ (.A(_00370_),
    .B(_00428_),
    .X(_00429_));
 sky130_fd_sc_hd__xor2_4 _07277_ (.A(_06127_),
    .B(_06479_),
    .X(_00430_));
 sky130_fd_sc_hd__xnor2_1 _07278_ (.A(_06127_),
    .B(_06479_),
    .Y(_00431_));
 sky130_fd_sc_hd__o22a_1 _07279_ (.A1(net127),
    .A2(net95),
    .B1(net92),
    .B2(net42),
    .X(_00432_));
 sky130_fd_sc_hd__xnor2_1 _07280_ (.A(net138),
    .B(_00432_),
    .Y(_00433_));
 sky130_fd_sc_hd__o41a_4 _07281_ (.A1(reg1_val[13]),
    .A2(_06433_),
    .A3(_00238_),
    .A4(_00240_),
    .B1(net274),
    .X(_00434_));
 sky130_fd_sc_hd__xor2_2 _07282_ (.A(reg1_val[19]),
    .B(_00434_),
    .X(_00435_));
 sky130_fd_sc_hd__xnor2_4 _07283_ (.A(reg1_val[19]),
    .B(_00434_),
    .Y(_00436_));
 sky130_fd_sc_hd__xnor2_2 _07284_ (.A(reg1_val[20]),
    .B(_00268_),
    .Y(_00437_));
 sky130_fd_sc_hd__or2_1 _07285_ (.A(_00436_),
    .B(_00437_),
    .X(_00438_));
 sky130_fd_sc_hd__nand2_1 _07286_ (.A(_00436_),
    .B(_00437_),
    .Y(_00439_));
 sky130_fd_sc_hd__mux2_2 _07287_ (.A0(_00438_),
    .A1(_00439_),
    .S(net103),
    .X(_00440_));
 sky130_fd_sc_hd__o31a_1 _07288_ (.A1(_06252_),
    .A2(_06448_),
    .A3(_06449_),
    .B1(net193),
    .X(_00441_));
 sky130_fd_sc_hd__nor2_1 _07289_ (.A(_06246_),
    .B(_06447_),
    .Y(_00442_));
 sky130_fd_sc_hd__a2bb2o_1 _07290_ (.A1_N(_06245_),
    .A2_N(_00441_),
    .B1(_00442_),
    .B2(_06451_),
    .X(_00443_));
 sky130_fd_sc_hd__nand2_2 _07291_ (.A(_00438_),
    .B(_00439_),
    .Y(_00444_));
 sky130_fd_sc_hd__o22a_1 _07292_ (.A1(net144),
    .A2(net40),
    .B1(net134),
    .B2(net38),
    .X(_00445_));
 sky130_fd_sc_hd__xnor2_1 _07293_ (.A(net103),
    .B(_00445_),
    .Y(_00446_));
 sky130_fd_sc_hd__xor2_1 _07294_ (.A(_00433_),
    .B(_00446_),
    .X(_00447_));
 sky130_fd_sc_hd__or2_1 _07295_ (.A(_00441_),
    .B(_00442_),
    .X(_00448_));
 sky130_fd_sc_hd__xnor2_1 _07296_ (.A(_06233_),
    .B(_00448_),
    .Y(_00449_));
 sky130_fd_sc_hd__o41a_2 _07297_ (.A1(reg1_val[13]),
    .A2(_06433_),
    .A3(_00238_),
    .A4(_00239_),
    .B1(net274),
    .X(_00450_));
 sky130_fd_sc_hd__xor2_4 _07298_ (.A(reg1_val[18]),
    .B(_00450_),
    .X(_00451_));
 sky130_fd_sc_hd__and2_1 _07299_ (.A(net137),
    .B(_00451_),
    .X(_00452_));
 sky130_fd_sc_hd__and3_1 _07300_ (.A(net138),
    .B(_00436_),
    .C(_00451_),
    .X(_00453_));
 sky130_fd_sc_hd__nor2_1 _07301_ (.A(net137),
    .B(_00451_),
    .Y(_00454_));
 sky130_fd_sc_hd__a21oi_2 _07302_ (.A1(net135),
    .A2(_00454_),
    .B1(_00453_),
    .Y(_00455_));
 sky130_fd_sc_hd__and2_1 _07303_ (.A(net193),
    .B(_06453_),
    .X(_00456_));
 sky130_fd_sc_hd__xnor2_4 _07304_ (.A(_06181_),
    .B(_00456_),
    .Y(_00457_));
 sky130_fd_sc_hd__or2_4 _07305_ (.A(_00452_),
    .B(_00454_),
    .X(_00458_));
 sky130_fd_sc_hd__o22a_1 _07306_ (.A1(net91),
    .A2(net36),
    .B1(net88),
    .B2(_00458_),
    .X(_00459_));
 sky130_fd_sc_hd__xnor2_1 _07307_ (.A(net135),
    .B(_00459_),
    .Y(_00460_));
 sky130_fd_sc_hd__and2_1 _07308_ (.A(_00447_),
    .B(_00460_),
    .X(_00461_));
 sky130_fd_sc_hd__a21oi_1 _07309_ (.A1(_00433_),
    .A2(_00446_),
    .B1(_00461_),
    .Y(_00462_));
 sky130_fd_sc_hd__o22a_1 _07310_ (.A1(net36),
    .A2(net88),
    .B1(_00458_),
    .B2(net92),
    .X(_00463_));
 sky130_fd_sc_hd__xnor2_1 _07311_ (.A(_00436_),
    .B(_00463_),
    .Y(_00464_));
 sky130_fd_sc_hd__o22a_1 _07312_ (.A1(net40),
    .A2(net134),
    .B1(net38),
    .B2(net91),
    .X(_00465_));
 sky130_fd_sc_hd__xor2_1 _07313_ (.A(net103),
    .B(_00465_),
    .X(_00466_));
 sky130_fd_sc_hd__nor2_1 _07314_ (.A(_00464_),
    .B(_00466_),
    .Y(_00467_));
 sky130_fd_sc_hd__and2_1 _07315_ (.A(_00464_),
    .B(_00466_),
    .X(_00468_));
 sky130_fd_sc_hd__nor2_1 _07316_ (.A(_00467_),
    .B(_00468_),
    .Y(_00469_));
 sky130_fd_sc_hd__o22a_1 _07317_ (.A1(net147),
    .A2(net49),
    .B1(net141),
    .B2(net51),
    .X(_00470_));
 sky130_fd_sc_hd__xnor2_1 _07318_ (.A(net107),
    .B(_00470_),
    .Y(_00471_));
 sky130_fd_sc_hd__o22a_1 _07319_ (.A1(net165),
    .A2(net53),
    .B1(net161),
    .B2(net15),
    .X(_00472_));
 sky130_fd_sc_hd__xnor2_1 _07320_ (.A(net113),
    .B(_00472_),
    .Y(_00473_));
 sky130_fd_sc_hd__and2_1 _07321_ (.A(_00471_),
    .B(_00473_),
    .X(_00474_));
 sky130_fd_sc_hd__xor2_1 _07322_ (.A(_00471_),
    .B(_00473_),
    .X(_00475_));
 sky130_fd_sc_hd__a22o_1 _07323_ (.A1(_00263_),
    .A2(_00307_),
    .B1(_00308_),
    .B2(_00300_),
    .X(_00476_));
 sky130_fd_sc_hd__xor2_1 _07324_ (.A(net110),
    .B(_00476_),
    .X(_00477_));
 sky130_fd_sc_hd__and2_1 _07325_ (.A(_00475_),
    .B(_00477_),
    .X(_00478_));
 sky130_fd_sc_hd__o21a_1 _07326_ (.A1(_00474_),
    .A2(_00478_),
    .B1(_00469_),
    .X(_00479_));
 sky130_fd_sc_hd__or3_1 _07327_ (.A(_00469_),
    .B(_00474_),
    .C(_00478_),
    .X(_00480_));
 sky130_fd_sc_hd__and2b_1 _07328_ (.A_N(_00479_),
    .B(_00480_),
    .X(_00481_));
 sky130_fd_sc_hd__and2b_1 _07329_ (.A_N(_00462_),
    .B(_00481_),
    .X(_00482_));
 sky130_fd_sc_hd__xnor2_1 _07330_ (.A(_00462_),
    .B(_00481_),
    .Y(_00483_));
 sky130_fd_sc_hd__and2_1 _07331_ (.A(_00429_),
    .B(_00483_),
    .X(_00484_));
 sky130_fd_sc_hd__nor2_1 _07332_ (.A(_00429_),
    .B(_00483_),
    .Y(_00485_));
 sky130_fd_sc_hd__nor2_1 _07333_ (.A(_00484_),
    .B(_00485_),
    .Y(_00486_));
 sky130_fd_sc_hd__xor2_1 _07334_ (.A(_00359_),
    .B(_00486_),
    .X(_00487_));
 sky130_fd_sc_hd__nor3_1 _07335_ (.A(_00348_),
    .B(_00352_),
    .C(_00353_),
    .Y(_00488_));
 sky130_fd_sc_hd__or2_1 _07336_ (.A(_00354_),
    .B(_00488_),
    .X(_00489_));
 sky130_fd_sc_hd__xor2_1 _07337_ (.A(_00475_),
    .B(_00477_),
    .X(_00490_));
 sky130_fd_sc_hd__inv_2 _07338_ (.A(_00490_),
    .Y(_00491_));
 sky130_fd_sc_hd__xnor2_1 _07339_ (.A(_00235_),
    .B(_00236_),
    .Y(_00492_));
 sky130_fd_sc_hd__or2_1 _07340_ (.A(_00491_),
    .B(_00492_),
    .X(_00493_));
 sky130_fd_sc_hd__xnor2_1 _07341_ (.A(_00491_),
    .B(_00492_),
    .Y(_00494_));
 sky130_fd_sc_hd__or2_1 _07342_ (.A(_00489_),
    .B(_00494_),
    .X(_00495_));
 sky130_fd_sc_hd__nand2_1 _07343_ (.A(_00489_),
    .B(_00494_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_1 _07344_ (.A(_00495_),
    .B(_00496_),
    .Y(_00497_));
 sky130_fd_sc_hd__o22a_1 _07345_ (.A1(_00391_),
    .A2(net92),
    .B1(net88),
    .B2(net42),
    .X(_00498_));
 sky130_fd_sc_hd__xnor2_1 _07346_ (.A(net138),
    .B(_00498_),
    .Y(_00499_));
 sky130_fd_sc_hd__o22a_1 _07347_ (.A1(net147),
    .A2(net40),
    .B1(net38),
    .B2(net144),
    .X(_00500_));
 sky130_fd_sc_hd__xnor2_1 _07348_ (.A(net103),
    .B(_00500_),
    .Y(_00501_));
 sky130_fd_sc_hd__xnor2_1 _07349_ (.A(_00499_),
    .B(_00501_),
    .Y(_00502_));
 sky130_fd_sc_hd__o22a_1 _07350_ (.A1(net134),
    .A2(net36),
    .B1(net35),
    .B2(net91),
    .X(_00503_));
 sky130_fd_sc_hd__xnor2_1 _07351_ (.A(_00436_),
    .B(_00503_),
    .Y(_00504_));
 sky130_fd_sc_hd__nor2_1 _07352_ (.A(_00502_),
    .B(_00504_),
    .Y(_00505_));
 sky130_fd_sc_hd__a21o_1 _07353_ (.A1(_00499_),
    .A2(_00501_),
    .B1(_00505_),
    .X(_00506_));
 sky130_fd_sc_hd__xor2_2 _07354_ (.A(_00361_),
    .B(_00363_),
    .X(_00507_));
 sky130_fd_sc_hd__o22a_1 _07355_ (.A1(net51),
    .A2(net143),
    .B1(net141),
    .B2(net49),
    .X(_00508_));
 sky130_fd_sc_hd__xor2_1 _07356_ (.A(net107),
    .B(_00508_),
    .X(_00509_));
 sky130_fd_sc_hd__o22a_1 _07357_ (.A1(net15),
    .A2(net163),
    .B1(net161),
    .B2(net53),
    .X(_00510_));
 sky130_fd_sc_hd__nand2_1 _07358_ (.A(net113),
    .B(_00510_),
    .Y(_00511_));
 sky130_fd_sc_hd__or2_1 _07359_ (.A(net113),
    .B(_00510_),
    .X(_00512_));
 sky130_fd_sc_hd__a21o_1 _07360_ (.A1(_00511_),
    .A2(_00512_),
    .B1(_00509_),
    .X(_00513_));
 sky130_fd_sc_hd__nand3_1 _07361_ (.A(_00509_),
    .B(_00511_),
    .C(_00512_),
    .Y(_00514_));
 sky130_fd_sc_hd__a22o_1 _07362_ (.A1(_00252_),
    .A2(_00307_),
    .B1(_00308_),
    .B2(_00263_),
    .X(_00515_));
 sky130_fd_sc_hd__xor2_2 _07363_ (.A(net110),
    .B(_00515_),
    .X(_00516_));
 sky130_fd_sc_hd__and3_1 _07364_ (.A(_00513_),
    .B(_00514_),
    .C(_00516_),
    .X(_00517_));
 sky130_fd_sc_hd__a21boi_2 _07365_ (.A1(_00514_),
    .A2(_00516_),
    .B1_N(_00513_),
    .Y(_00518_));
 sky130_fd_sc_hd__xor2_1 _07366_ (.A(_00507_),
    .B(_00518_),
    .X(_00519_));
 sky130_fd_sc_hd__nand2_1 _07367_ (.A(_00506_),
    .B(_00519_),
    .Y(_00520_));
 sky130_fd_sc_hd__or2_1 _07368_ (.A(_00506_),
    .B(_00519_),
    .X(_00521_));
 sky130_fd_sc_hd__and2_1 _07369_ (.A(_00520_),
    .B(_00521_),
    .X(_00522_));
 sky130_fd_sc_hd__o22a_1 _07370_ (.A1(net77),
    .A2(net177),
    .B1(net175),
    .B2(net75),
    .X(_00523_));
 sky130_fd_sc_hd__xnor2_1 _07371_ (.A(net189),
    .B(_00523_),
    .Y(_00524_));
 sky130_fd_sc_hd__o22a_1 _07372_ (.A1(net152),
    .A2(net120),
    .B1(net72),
    .B2(net150),
    .X(_00525_));
 sky130_fd_sc_hd__xnor2_1 _07373_ (.A(net192),
    .B(_00525_),
    .Y(_00526_));
 sky130_fd_sc_hd__nor2_1 _07374_ (.A(_00524_),
    .B(_00526_),
    .Y(_00527_));
 sky130_fd_sc_hd__xnor2_1 _07375_ (.A(_00325_),
    .B(_00327_),
    .Y(_00528_));
 sky130_fd_sc_hd__nand2_1 _07376_ (.A(_00527_),
    .B(_00528_),
    .Y(_00529_));
 sky130_fd_sc_hd__xor2_1 _07377_ (.A(_00350_),
    .B(_00351_),
    .X(_00530_));
 sky130_fd_sc_hd__xnor2_1 _07378_ (.A(_00527_),
    .B(_00528_),
    .Y(_00531_));
 sky130_fd_sc_hd__o21a_1 _07379_ (.A1(_00530_),
    .A2(_00531_),
    .B1(_00529_),
    .X(_00532_));
 sky130_fd_sc_hd__nor2_1 _07380_ (.A(_00447_),
    .B(_00460_),
    .Y(_00533_));
 sky130_fd_sc_hd__nor2_1 _07381_ (.A(_00461_),
    .B(_00533_),
    .Y(_00534_));
 sky130_fd_sc_hd__o22a_1 _07382_ (.A1(net302),
    .A2(net61),
    .B1(net253),
    .B2(_00185_),
    .X(_00535_));
 sky130_fd_sc_hd__xnor2_2 _07383_ (.A(net255),
    .B(_00535_),
    .Y(_00536_));
 sky130_fd_sc_hd__o22a_1 _07384_ (.A1(net69),
    .A2(net169),
    .B1(net167),
    .B2(net66),
    .X(_00537_));
 sky130_fd_sc_hd__xnor2_1 _07385_ (.A(net210),
    .B(_00537_),
    .Y(_00538_));
 sky130_fd_sc_hd__nor2_1 _07386_ (.A(_00536_),
    .B(_00538_),
    .Y(_00539_));
 sky130_fd_sc_hd__o22a_1 _07387_ (.A1(net173),
    .A2(net59),
    .B1(net56),
    .B2(net171),
    .X(_00540_));
 sky130_fd_sc_hd__xnor2_1 _07388_ (.A(net208),
    .B(_00540_),
    .Y(_00541_));
 sky130_fd_sc_hd__xnor2_1 _07389_ (.A(_00536_),
    .B(_00538_),
    .Y(_00542_));
 sky130_fd_sc_hd__nor2_1 _07390_ (.A(_00541_),
    .B(_00542_),
    .Y(_00543_));
 sky130_fd_sc_hd__or4_1 _07391_ (.A(net226),
    .B(net46),
    .C(_00539_),
    .D(_00543_),
    .X(_00544_));
 sky130_fd_sc_hd__o21ai_1 _07392_ (.A1(net226),
    .A2(net46),
    .B1(net98),
    .Y(_00545_));
 sky130_fd_sc_hd__and3_1 _07393_ (.A(_00534_),
    .B(_00544_),
    .C(_00545_),
    .X(_00546_));
 sky130_fd_sc_hd__a21oi_1 _07394_ (.A1(_00544_),
    .A2(_00545_),
    .B1(_00534_),
    .Y(_00547_));
 sky130_fd_sc_hd__nor2_1 _07395_ (.A(_00546_),
    .B(_00547_),
    .Y(_00548_));
 sky130_fd_sc_hd__xnor2_2 _07396_ (.A(_00532_),
    .B(_00548_),
    .Y(_00549_));
 sky130_fd_sc_hd__xnor2_2 _07397_ (.A(_00497_),
    .B(_00522_),
    .Y(_00550_));
 sky130_fd_sc_hd__a32o_1 _07398_ (.A1(_00495_),
    .A2(_00496_),
    .A3(_00522_),
    .B1(_00549_),
    .B2(_00550_),
    .X(_00551_));
 sky130_fd_sc_hd__o21bai_2 _07399_ (.A1(_00532_),
    .A2(_00547_),
    .B1_N(_00546_),
    .Y(_00552_));
 sky130_fd_sc_hd__o21a_1 _07400_ (.A1(_00489_),
    .A2(_00494_),
    .B1(_00493_),
    .X(_00553_));
 sky130_fd_sc_hd__o21ai_2 _07401_ (.A1(_00507_),
    .A2(_00518_),
    .B1(_00520_),
    .Y(_00554_));
 sky130_fd_sc_hd__nand2b_1 _07402_ (.A_N(_00553_),
    .B(_00554_),
    .Y(_00555_));
 sky130_fd_sc_hd__xnor2_2 _07403_ (.A(_00553_),
    .B(_00554_),
    .Y(_00556_));
 sky130_fd_sc_hd__xnor2_2 _07404_ (.A(_00552_),
    .B(_00556_),
    .Y(_00557_));
 sky130_fd_sc_hd__xnor2_1 _07405_ (.A(_00530_),
    .B(_00531_),
    .Y(_00558_));
 sky130_fd_sc_hd__a21oi_1 _07406_ (.A1(_00513_),
    .A2(_00514_),
    .B1(_00516_),
    .Y(_00559_));
 sky130_fd_sc_hd__nor2_1 _07407_ (.A(_00517_),
    .B(_00559_),
    .Y(_00560_));
 sky130_fd_sc_hd__and2b_1 _07408_ (.A_N(_00558_),
    .B(_00560_),
    .X(_00561_));
 sky130_fd_sc_hd__xnor2_1 _07409_ (.A(_00558_),
    .B(_00560_),
    .Y(_00562_));
 sky130_fd_sc_hd__o22ai_1 _07410_ (.A1(net226),
    .A2(net46),
    .B1(_00539_),
    .B2(_00543_),
    .Y(_00563_));
 sky130_fd_sc_hd__and2_1 _07411_ (.A(_00544_),
    .B(_00563_),
    .X(_00564_));
 sky130_fd_sc_hd__inv_2 _07412_ (.A(_00564_),
    .Y(_00565_));
 sky130_fd_sc_hd__a21oi_1 _07413_ (.A1(_00562_),
    .A2(_00565_),
    .B1(_00561_),
    .Y(_00566_));
 sky130_fd_sc_hd__and2_1 _07414_ (.A(_06470_),
    .B(_06486_),
    .X(_00567_));
 sky130_fd_sc_hd__nor2_1 _07415_ (.A(_06487_),
    .B(_00567_),
    .Y(_00568_));
 sky130_fd_sc_hd__o22a_1 _07416_ (.A1(net42),
    .A2(net91),
    .B1(_00457_),
    .B2(net95),
    .X(_00569_));
 sky130_fd_sc_hd__xnor2_1 _07417_ (.A(net138),
    .B(_00569_),
    .Y(_00570_));
 sky130_fd_sc_hd__o22a_1 _07418_ (.A1(net141),
    .A2(net40),
    .B1(net38),
    .B2(net147),
    .X(_00571_));
 sky130_fd_sc_hd__xnor2_1 _07419_ (.A(net103),
    .B(_00571_),
    .Y(_00572_));
 sky130_fd_sc_hd__xor2_1 _07420_ (.A(_00570_),
    .B(_00572_),
    .X(_00573_));
 sky130_fd_sc_hd__o22a_1 _07421_ (.A1(net144),
    .A2(net36),
    .B1(net34),
    .B2(net134),
    .X(_00574_));
 sky130_fd_sc_hd__xnor2_1 _07422_ (.A(net135),
    .B(_00574_),
    .Y(_00575_));
 sky130_fd_sc_hd__and2_1 _07423_ (.A(_00573_),
    .B(_00575_),
    .X(_00576_));
 sky130_fd_sc_hd__a21o_1 _07424_ (.A1(_00570_),
    .A2(_00572_),
    .B1(_00576_),
    .X(_00577_));
 sky130_fd_sc_hd__o22a_1 _07425_ (.A1(net128),
    .A2(net116),
    .B1(net115),
    .B2(net101),
    .X(_00578_));
 sky130_fd_sc_hd__xnor2_2 _07426_ (.A(net180),
    .B(_00578_),
    .Y(_00579_));
 sky130_fd_sc_hd__o22a_1 _07427_ (.A1(net127),
    .A2(net123),
    .B1(net92),
    .B2(net78),
    .X(_00580_));
 sky130_fd_sc_hd__xor2_2 _07428_ (.A(net155),
    .B(_00580_),
    .X(_00581_));
 sky130_fd_sc_hd__xnor2_1 _07429_ (.A(_00579_),
    .B(_00581_),
    .Y(_00582_));
 sky130_fd_sc_hd__o22a_1 _07430_ (.A1(net80),
    .A2(net130),
    .B1(net121),
    .B2(net82),
    .X(_00583_));
 sky130_fd_sc_hd__xnor2_1 _07431_ (.A(net158),
    .B(_00583_),
    .Y(_00584_));
 sky130_fd_sc_hd__or2_1 _07432_ (.A(_00582_),
    .B(_00584_),
    .X(_00585_));
 sky130_fd_sc_hd__o21ai_2 _07433_ (.A1(_00579_),
    .A2(_00581_),
    .B1(_00585_),
    .Y(_00586_));
 sky130_fd_sc_hd__xnor2_1 _07434_ (.A(_00568_),
    .B(_00577_),
    .Y(_00587_));
 sky130_fd_sc_hd__and2b_1 _07435_ (.A_N(_00587_),
    .B(_00586_),
    .X(_00588_));
 sky130_fd_sc_hd__a21oi_1 _07436_ (.A1(_00568_),
    .A2(_00577_),
    .B1(_00588_),
    .Y(_00589_));
 sky130_fd_sc_hd__nor2_1 _07437_ (.A(_00566_),
    .B(_00589_),
    .Y(_00590_));
 sky130_fd_sc_hd__and2_1 _07438_ (.A(_00502_),
    .B(_00504_),
    .X(_00591_));
 sky130_fd_sc_hd__nor2_1 _07439_ (.A(_00505_),
    .B(_00591_),
    .Y(_00592_));
 sky130_fd_sc_hd__o22a_1 _07440_ (.A1(net226),
    .A2(net15),
    .B1(net53),
    .B2(net163),
    .X(_00593_));
 sky130_fd_sc_hd__xnor2_1 _07441_ (.A(net113),
    .B(_00593_),
    .Y(_00594_));
 sky130_fd_sc_hd__o22a_1 _07442_ (.A1(net149),
    .A2(net51),
    .B1(net49),
    .B2(net143),
    .X(_00595_));
 sky130_fd_sc_hd__xnor2_1 _07443_ (.A(net107),
    .B(_00595_),
    .Y(_00596_));
 sky130_fd_sc_hd__xor2_1 _07444_ (.A(_00594_),
    .B(_00596_),
    .X(_00597_));
 sky130_fd_sc_hd__a22o_1 _07445_ (.A1(_00252_),
    .A2(_00308_),
    .B1(_00424_),
    .B2(_00307_),
    .X(_00598_));
 sky130_fd_sc_hd__xor2_2 _07446_ (.A(net110),
    .B(_00598_),
    .X(_00599_));
 sky130_fd_sc_hd__and2_1 _07447_ (.A(_00597_),
    .B(_00599_),
    .X(_00600_));
 sky130_fd_sc_hd__a21o_1 _07448_ (.A1(_00594_),
    .A2(_00596_),
    .B1(_00600_),
    .X(_00601_));
 sky130_fd_sc_hd__xor2_1 _07449_ (.A(_00541_),
    .B(_00542_),
    .X(_00602_));
 sky130_fd_sc_hd__o22a_1 _07450_ (.A1(net75),
    .A2(net169),
    .B1(net167),
    .B2(net69),
    .X(_00603_));
 sky130_fd_sc_hd__xnor2_2 _07451_ (.A(net210),
    .B(_00603_),
    .Y(_00604_));
 sky130_fd_sc_hd__o22a_1 _07452_ (.A1(net302),
    .A2(_00185_),
    .B1(net56),
    .B2(net253),
    .X(_00605_));
 sky130_fd_sc_hd__xnor2_2 _07453_ (.A(net255),
    .B(_00605_),
    .Y(_00606_));
 sky130_fd_sc_hd__nor2_1 _07454_ (.A(_00604_),
    .B(_00606_),
    .Y(_00607_));
 sky130_fd_sc_hd__o22a_1 _07455_ (.A1(net66),
    .A2(net173),
    .B1(net171),
    .B2(net59),
    .X(_00608_));
 sky130_fd_sc_hd__xnor2_2 _07456_ (.A(net208),
    .B(_00608_),
    .Y(_00609_));
 sky130_fd_sc_hd__inv_2 _07457_ (.A(_00609_),
    .Y(_00610_));
 sky130_fd_sc_hd__xor2_2 _07458_ (.A(_00604_),
    .B(_00606_),
    .X(_00611_));
 sky130_fd_sc_hd__a21o_1 _07459_ (.A1(_00610_),
    .A2(_00611_),
    .B1(_00607_),
    .X(_00612_));
 sky130_fd_sc_hd__and2_1 _07460_ (.A(_00602_),
    .B(_00612_),
    .X(_00613_));
 sky130_fd_sc_hd__o22a_1 _07461_ (.A1(net72),
    .A2(net177),
    .B1(net175),
    .B2(net77),
    .X(_00614_));
 sky130_fd_sc_hd__xnor2_1 _07462_ (.A(net189),
    .B(_00614_),
    .Y(_00615_));
 sky130_fd_sc_hd__o22a_1 _07463_ (.A1(net150),
    .A2(net120),
    .B1(net101),
    .B2(net152),
    .X(_00616_));
 sky130_fd_sc_hd__xnor2_1 _07464_ (.A(_06489_),
    .B(_00616_),
    .Y(_00617_));
 sky130_fd_sc_hd__nor2_1 _07465_ (.A(_00615_),
    .B(_00617_),
    .Y(_00618_));
 sky130_fd_sc_hd__xor2_1 _07466_ (.A(_00602_),
    .B(_00612_),
    .X(_00619_));
 sky130_fd_sc_hd__a21o_1 _07467_ (.A1(_00618_),
    .A2(_00619_),
    .B1(_00613_),
    .X(_00620_));
 sky130_fd_sc_hd__xnor2_1 _07468_ (.A(_00592_),
    .B(_00601_),
    .Y(_00621_));
 sky130_fd_sc_hd__nand2b_1 _07469_ (.A_N(_00621_),
    .B(_00620_),
    .Y(_00622_));
 sky130_fd_sc_hd__a21bo_1 _07470_ (.A1(_00592_),
    .A2(_00601_),
    .B1_N(_00622_),
    .X(_00623_));
 sky130_fd_sc_hd__xor2_1 _07471_ (.A(_00566_),
    .B(_00589_),
    .X(_00624_));
 sky130_fd_sc_hd__a21oi_2 _07472_ (.A1(_00623_),
    .A2(_00624_),
    .B1(_00590_),
    .Y(_00625_));
 sky130_fd_sc_hd__xnor2_1 _07473_ (.A(_00557_),
    .B(_00625_),
    .Y(_00626_));
 sky130_fd_sc_hd__nand2b_1 _07474_ (.A_N(_00626_),
    .B(_00551_),
    .Y(_00627_));
 sky130_fd_sc_hd__xnor2_1 _07475_ (.A(_00551_),
    .B(_00626_),
    .Y(_00628_));
 sky130_fd_sc_hd__nand2_1 _07476_ (.A(_00487_),
    .B(_00628_),
    .Y(_00629_));
 sky130_fd_sc_hd__and2_1 _07477_ (.A(_00524_),
    .B(_00526_),
    .X(_00630_));
 sky130_fd_sc_hd__nor2_1 _07478_ (.A(_00527_),
    .B(_00630_),
    .Y(_00631_));
 sky130_fd_sc_hd__o22a_1 _07479_ (.A1(net43),
    .A2(net134),
    .B1(net91),
    .B2(net95),
    .X(_00632_));
 sky130_fd_sc_hd__xnor2_1 _07480_ (.A(net138),
    .B(_00632_),
    .Y(_00633_));
 sky130_fd_sc_hd__o22a_1 _07481_ (.A1(net143),
    .A2(_00440_),
    .B1(_00444_),
    .B2(net141),
    .X(_00634_));
 sky130_fd_sc_hd__xnor2_1 _07482_ (.A(net103),
    .B(_00634_),
    .Y(_00635_));
 sky130_fd_sc_hd__and2_1 _07483_ (.A(_00633_),
    .B(_00635_),
    .X(_00636_));
 sky130_fd_sc_hd__xor2_1 _07484_ (.A(_00633_),
    .B(_00635_),
    .X(_00637_));
 sky130_fd_sc_hd__o22a_1 _07485_ (.A1(net147),
    .A2(net36),
    .B1(net34),
    .B2(_00290_),
    .X(_00638_));
 sky130_fd_sc_hd__xnor2_1 _07486_ (.A(net136),
    .B(_00638_),
    .Y(_00639_));
 sky130_fd_sc_hd__and2_1 _07487_ (.A(_00637_),
    .B(_00639_),
    .X(_00640_));
 sky130_fd_sc_hd__o21ai_1 _07488_ (.A1(_00636_),
    .A2(_00640_),
    .B1(_00631_),
    .Y(_00641_));
 sky130_fd_sc_hd__or3_1 _07489_ (.A(_00631_),
    .B(_00636_),
    .C(_00640_),
    .X(_00642_));
 sky130_fd_sc_hd__nand2_1 _07490_ (.A(_00641_),
    .B(_00642_),
    .Y(_00643_));
 sky130_fd_sc_hd__o22a_1 _07491_ (.A1(net80),
    .A2(net117),
    .B1(net115),
    .B2(net128),
    .X(_00644_));
 sky130_fd_sc_hd__xnor2_2 _07492_ (.A(net180),
    .B(_00644_),
    .Y(_00645_));
 sky130_fd_sc_hd__o22a_1 _07493_ (.A1(net123),
    .A2(net92),
    .B1(_00457_),
    .B2(net78),
    .X(_00646_));
 sky130_fd_sc_hd__xor2_1 _07494_ (.A(net155),
    .B(_00646_),
    .X(_00647_));
 sky130_fd_sc_hd__xnor2_1 _07495_ (.A(_00645_),
    .B(_00647_),
    .Y(_00648_));
 sky130_fd_sc_hd__o22a_1 _07496_ (.A1(net82),
    .A2(net127),
    .B1(net121),
    .B2(net130),
    .X(_00649_));
 sky130_fd_sc_hd__xnor2_1 _07497_ (.A(net158),
    .B(_00649_),
    .Y(_00650_));
 sky130_fd_sc_hd__or2_1 _07498_ (.A(_00648_),
    .B(_00650_),
    .X(_00651_));
 sky130_fd_sc_hd__o21ai_2 _07499_ (.A1(_00645_),
    .A2(_00647_),
    .B1(_00651_),
    .Y(_00652_));
 sky130_fd_sc_hd__nand2b_1 _07500_ (.A_N(_00643_),
    .B(_00652_),
    .Y(_00653_));
 sky130_fd_sc_hd__nand2_1 _07501_ (.A(_00641_),
    .B(_00653_),
    .Y(_00654_));
 sky130_fd_sc_hd__xnor2_1 _07502_ (.A(_00618_),
    .B(_00619_),
    .Y(_00655_));
 sky130_fd_sc_hd__nor2_1 _07503_ (.A(_00573_),
    .B(_00575_),
    .Y(_00656_));
 sky130_fd_sc_hd__nor2_1 _07504_ (.A(_00576_),
    .B(_00656_),
    .Y(_00657_));
 sky130_fd_sc_hd__and2b_1 _07505_ (.A_N(_00655_),
    .B(_00657_),
    .X(_00658_));
 sky130_fd_sc_hd__nor2_1 _07506_ (.A(_00597_),
    .B(_00599_),
    .Y(_00659_));
 sky130_fd_sc_hd__nor2_1 _07507_ (.A(_00600_),
    .B(_00659_),
    .Y(_00660_));
 sky130_fd_sc_hd__xnor2_1 _07508_ (.A(_00655_),
    .B(_00657_),
    .Y(_00661_));
 sky130_fd_sc_hd__a21oi_1 _07509_ (.A1(_00660_),
    .A2(_00661_),
    .B1(_00658_),
    .Y(_00662_));
 sky130_fd_sc_hd__a21o_1 _07510_ (.A1(_00641_),
    .A2(_00653_),
    .B1(_00662_),
    .X(_00663_));
 sky130_fd_sc_hd__o22a_1 _07511_ (.A1(net165),
    .A2(net51),
    .B1(net49),
    .B2(net149),
    .X(_00664_));
 sky130_fd_sc_hd__xnor2_1 _07512_ (.A(net107),
    .B(_00664_),
    .Y(_00665_));
 sky130_fd_sc_hd__or2_1 _07513_ (.A(net226),
    .B(net53),
    .X(_00666_));
 sky130_fd_sc_hd__xnor2_1 _07514_ (.A(net113),
    .B(_00666_),
    .Y(_00667_));
 sky130_fd_sc_hd__nand2_1 _07515_ (.A(_00665_),
    .B(_00667_),
    .Y(_00668_));
 sky130_fd_sc_hd__or2_1 _07516_ (.A(_00665_),
    .B(_00667_),
    .X(_00669_));
 sky130_fd_sc_hd__nand2_1 _07517_ (.A(_00668_),
    .B(_00669_),
    .Y(_00670_));
 sky130_fd_sc_hd__a22o_1 _07518_ (.A1(_00307_),
    .A2(_00338_),
    .B1(_00424_),
    .B2(_00308_),
    .X(_00671_));
 sky130_fd_sc_hd__xnor2_1 _07519_ (.A(net110),
    .B(_00671_),
    .Y(_00672_));
 sky130_fd_sc_hd__or2_1 _07520_ (.A(_00670_),
    .B(_00672_),
    .X(_00673_));
 sky130_fd_sc_hd__nand2_1 _07521_ (.A(_00582_),
    .B(_00584_),
    .Y(_00674_));
 sky130_fd_sc_hd__nand2_1 _07522_ (.A(_00585_),
    .B(_00674_),
    .Y(_00675_));
 sky130_fd_sc_hd__a21oi_1 _07523_ (.A1(_00668_),
    .A2(_00673_),
    .B1(_00675_),
    .Y(_00676_));
 sky130_fd_sc_hd__xnor2_2 _07524_ (.A(_00609_),
    .B(_00611_),
    .Y(_00677_));
 sky130_fd_sc_hd__xnor2_2 _07525_ (.A(net113),
    .B(_00677_),
    .Y(_00678_));
 sky130_fd_sc_hd__o22a_1 _07526_ (.A1(net69),
    .A2(net173),
    .B1(net171),
    .B2(net66),
    .X(_00679_));
 sky130_fd_sc_hd__xnor2_1 _07527_ (.A(net208),
    .B(_00679_),
    .Y(_00680_));
 sky130_fd_sc_hd__o22a_1 _07528_ (.A1(net302),
    .A2(net56),
    .B1(net253),
    .B2(net59),
    .X(_00681_));
 sky130_fd_sc_hd__xnor2_1 _07529_ (.A(net255),
    .B(_00681_),
    .Y(_00682_));
 sky130_fd_sc_hd__nor2_1 _07530_ (.A(_00680_),
    .B(_00682_),
    .Y(_00683_));
 sky130_fd_sc_hd__or3_1 _07531_ (.A(_00678_),
    .B(_00680_),
    .C(_00682_),
    .X(_00684_));
 sky130_fd_sc_hd__a21bo_1 _07532_ (.A1(net113),
    .A2(_00677_),
    .B1_N(_00684_),
    .X(_00685_));
 sky130_fd_sc_hd__and3_1 _07533_ (.A(_00668_),
    .B(_00673_),
    .C(_00675_),
    .X(_00686_));
 sky130_fd_sc_hd__nor2_1 _07534_ (.A(_00676_),
    .B(_00686_),
    .Y(_00687_));
 sky130_fd_sc_hd__a21o_1 _07535_ (.A1(_00685_),
    .A2(_00687_),
    .B1(_00676_),
    .X(_00688_));
 sky130_fd_sc_hd__xnor2_1 _07536_ (.A(_00654_),
    .B(_00662_),
    .Y(_00689_));
 sky130_fd_sc_hd__nand2_1 _07537_ (.A(_00688_),
    .B(_00689_),
    .Y(_00690_));
 sky130_fd_sc_hd__xnor2_1 _07538_ (.A(_00623_),
    .B(_00624_),
    .Y(_00691_));
 sky130_fd_sc_hd__a21o_1 _07539_ (.A1(_00663_),
    .A2(_00690_),
    .B1(_00691_),
    .X(_00692_));
 sky130_fd_sc_hd__xnor2_1 _07540_ (.A(_00562_),
    .B(_00564_),
    .Y(_00693_));
 sky130_fd_sc_hd__xnor2_1 _07541_ (.A(_00586_),
    .B(_00587_),
    .Y(_00694_));
 sky130_fd_sc_hd__xor2_1 _07542_ (.A(_00620_),
    .B(_00621_),
    .X(_00695_));
 sky130_fd_sc_hd__xnor2_1 _07543_ (.A(_00693_),
    .B(_00694_),
    .Y(_00696_));
 sky130_fd_sc_hd__or2_1 _07544_ (.A(_00695_),
    .B(_00696_),
    .X(_00697_));
 sky130_fd_sc_hd__a21bo_1 _07545_ (.A1(_00693_),
    .A2(_00694_),
    .B1_N(_00697_),
    .X(_00698_));
 sky130_fd_sc_hd__nand3_1 _07546_ (.A(_00663_),
    .B(_00690_),
    .C(_00691_),
    .Y(_00699_));
 sky130_fd_sc_hd__nand2_1 _07547_ (.A(_00692_),
    .B(_00699_),
    .Y(_00700_));
 sky130_fd_sc_hd__nand2b_1 _07548_ (.A_N(_00700_),
    .B(_00698_),
    .Y(_00701_));
 sky130_fd_sc_hd__or2_1 _07549_ (.A(_00487_),
    .B(_00628_),
    .X(_00702_));
 sky130_fd_sc_hd__nand2_1 _07550_ (.A(_00629_),
    .B(_00702_),
    .Y(_00703_));
 sky130_fd_sc_hd__a21o_1 _07551_ (.A1(_00692_),
    .A2(_00701_),
    .B1(_00703_),
    .X(_00704_));
 sky130_fd_sc_hd__o21ai_2 _07552_ (.A1(_00557_),
    .A2(_00625_),
    .B1(_00627_),
    .Y(_00705_));
 sky130_fd_sc_hd__a32oi_4 _07553_ (.A1(_00400_),
    .A2(_00401_),
    .A3(_00413_),
    .B1(_00414_),
    .B2(_00380_),
    .Y(_00706_));
 sky130_fd_sc_hd__o22a_1 _07554_ (.A1(net15),
    .A2(net149),
    .B1(net53),
    .B2(net143),
    .X(_00707_));
 sky130_fd_sc_hd__xnor2_1 _07555_ (.A(net113),
    .B(_00707_),
    .Y(_00708_));
 sky130_fd_sc_hd__o22a_1 _07556_ (.A1(net51),
    .A2(_00290_),
    .B1(net49),
    .B2(net134),
    .X(_00709_));
 sky130_fd_sc_hd__xnor2_1 _07557_ (.A(net107),
    .B(_00709_),
    .Y(_00710_));
 sky130_fd_sc_hd__and2_1 _07558_ (.A(_00708_),
    .B(_00710_),
    .X(_00711_));
 sky130_fd_sc_hd__nor2_1 _07559_ (.A(_00708_),
    .B(_00710_),
    .Y(_00712_));
 sky130_fd_sc_hd__nor2_1 _07560_ (.A(_00711_),
    .B(_00712_),
    .Y(_00713_));
 sky130_fd_sc_hd__a22o_1 _07561_ (.A1(_00276_),
    .A2(_00308_),
    .B1(_00310_),
    .B2(_00307_),
    .X(_00714_));
 sky130_fd_sc_hd__xnor2_2 _07562_ (.A(net110),
    .B(_00714_),
    .Y(_00715_));
 sky130_fd_sc_hd__xnor2_1 _07563_ (.A(_00713_),
    .B(_00715_),
    .Y(_00716_));
 sky130_fd_sc_hd__o21ai_2 _07564_ (.A1(_00366_),
    .A2(_00368_),
    .B1(_00716_),
    .Y(_00717_));
 sky130_fd_sc_hd__or3_1 _07565_ (.A(_00366_),
    .B(_00368_),
    .C(_00716_),
    .X(_00718_));
 sky130_fd_sc_hd__nand2_1 _07566_ (.A(_00717_),
    .B(_00718_),
    .Y(_00719_));
 sky130_fd_sc_hd__xor2_1 _07567_ (.A(_00706_),
    .B(_00719_),
    .X(_00720_));
 sky130_fd_sc_hd__o21ai_1 _07568_ (.A1(_00377_),
    .A2(_00379_),
    .B1(_00467_),
    .Y(_00721_));
 sky130_fd_sc_hd__or3_1 _07569_ (.A(_00377_),
    .B(_00379_),
    .C(_00467_),
    .X(_00722_));
 sky130_fd_sc_hd__and2_1 _07570_ (.A(_00721_),
    .B(_00722_),
    .X(_00723_));
 sky130_fd_sc_hd__o21ai_1 _07571_ (.A1(_00395_),
    .A2(_00399_),
    .B1(_00723_),
    .Y(_00724_));
 sky130_fd_sc_hd__or3_1 _07572_ (.A(_00395_),
    .B(_00399_),
    .C(_00723_),
    .X(_00725_));
 sky130_fd_sc_hd__nand2_1 _07573_ (.A(_00724_),
    .B(_00725_),
    .Y(_00726_));
 sky130_fd_sc_hd__nor2_1 _07574_ (.A(reg1_val[30]),
    .B(_00416_),
    .Y(_00727_));
 sky130_fd_sc_hd__o21a_2 _07575_ (.A1(_04504_),
    .A2(_00727_),
    .B1(reg1_val[31]),
    .X(_00728_));
 sky130_fd_sc_hd__o21ai_1 _07576_ (.A1(_04504_),
    .A2(_00727_),
    .B1(reg1_val[31]),
    .Y(_00729_));
 sky130_fd_sc_hd__mux2_1 _07577_ (.A0(_00419_),
    .A1(_00420_),
    .S(net33),
    .X(_00730_));
 sky130_fd_sc_hd__o22a_1 _07578_ (.A1(net163),
    .A2(net8),
    .B1(net6),
    .B2(_06309_),
    .X(_00731_));
 sky130_fd_sc_hd__xnor2_2 _07579_ (.A(net32),
    .B(_00731_),
    .Y(_00732_));
 sky130_fd_sc_hd__a21oi_2 _07580_ (.A1(_00404_),
    .A2(_00412_),
    .B1(_00411_),
    .Y(_00733_));
 sky130_fd_sc_hd__o22a_1 _07581_ (.A1(net165),
    .A2(net46),
    .B1(net161),
    .B2(net12),
    .X(_00734_));
 sky130_fd_sc_hd__xnor2_2 _07582_ (.A(net98),
    .B(_00734_),
    .Y(_00735_));
 sky130_fd_sc_hd__or2_1 _07583_ (.A(_00733_),
    .B(_00735_),
    .X(_00736_));
 sky130_fd_sc_hd__xnor2_2 _07584_ (.A(_00733_),
    .B(_00735_),
    .Y(_00737_));
 sky130_fd_sc_hd__xnor2_2 _07585_ (.A(_00732_),
    .B(_00737_),
    .Y(_00738_));
 sky130_fd_sc_hd__o22a_1 _07586_ (.A1(net152),
    .A2(net68),
    .B1(net65),
    .B2(net150),
    .X(_00739_));
 sky130_fd_sc_hd__xnor2_1 _07587_ (.A(_06489_),
    .B(_00739_),
    .Y(_00740_));
 sky130_fd_sc_hd__inv_2 _07588_ (.A(_00740_),
    .Y(_00741_));
 sky130_fd_sc_hd__o22a_1 _07589_ (.A1(net177),
    .A2(net57),
    .B1(net54),
    .B2(net175),
    .X(_00742_));
 sky130_fd_sc_hd__xnor2_1 _07590_ (.A(net189),
    .B(_00742_),
    .Y(_00743_));
 sky130_fd_sc_hd__o22a_1 _07591_ (.A1(net77),
    .A2(net116),
    .B1(net114),
    .B2(net74),
    .X(_00744_));
 sky130_fd_sc_hd__xnor2_1 _07592_ (.A(net180),
    .B(_00744_),
    .Y(_00745_));
 sky130_fd_sc_hd__nor2_1 _07593_ (.A(_00743_),
    .B(_00745_),
    .Y(_00746_));
 sky130_fd_sc_hd__xor2_1 _07594_ (.A(_00743_),
    .B(_00745_),
    .X(_00747_));
 sky130_fd_sc_hd__xnor2_1 _07595_ (.A(_00740_),
    .B(_00747_),
    .Y(_00748_));
 sky130_fd_sc_hd__inv_2 _07596_ (.A(_00748_),
    .Y(_00749_));
 sky130_fd_sc_hd__o22a_2 _07597_ (.A1(net173),
    .A2(_00223_),
    .B1(net16),
    .B2(net171),
    .X(_00750_));
 sky130_fd_sc_hd__xnor2_4 _07598_ (.A(net208),
    .B(_00750_),
    .Y(_00751_));
 sky130_fd_sc_hd__inv_2 _07599_ (.A(_00751_),
    .Y(_00752_));
 sky130_fd_sc_hd__o22a_2 _07600_ (.A1(net63),
    .A2(net169),
    .B1(net167),
    .B2(net61),
    .X(_00753_));
 sky130_fd_sc_hd__xnor2_4 _07601_ (.A(net210),
    .B(_00753_),
    .Y(_00754_));
 sky130_fd_sc_hd__o41a_1 _07602_ (.A1(_05046_),
    .A2(_05198_),
    .A3(_05263_),
    .A4(_00218_),
    .B1(net307),
    .X(_00755_));
 sky130_fd_sc_hd__nor2_4 _07603_ (.A(_04741_),
    .B(_00755_),
    .Y(_00756_));
 sky130_fd_sc_hd__or2_2 _07604_ (.A(_04741_),
    .B(_00755_),
    .X(_00757_));
 sky130_fd_sc_hd__o22a_1 _07605_ (.A1(net253),
    .A2(net10),
    .B1(net4),
    .B2(net302),
    .X(_00758_));
 sky130_fd_sc_hd__xnor2_2 _07606_ (.A(net255),
    .B(_00758_),
    .Y(_00759_));
 sky130_fd_sc_hd__nor2_1 _07607_ (.A(_00754_),
    .B(_00759_),
    .Y(_00760_));
 sky130_fd_sc_hd__xor2_4 _07608_ (.A(_00754_),
    .B(_00759_),
    .X(_00761_));
 sky130_fd_sc_hd__xnor2_4 _07609_ (.A(_00751_),
    .B(_00761_),
    .Y(_00762_));
 sky130_fd_sc_hd__o22a_1 _07610_ (.A1(_06484_),
    .A2(net43),
    .B1(net94),
    .B2(net80),
    .X(_00763_));
 sky130_fd_sc_hd__xnor2_2 _07611_ (.A(net137),
    .B(_00763_),
    .Y(_00764_));
 sky130_fd_sc_hd__inv_2 _07612_ (.A(_00764_),
    .Y(_00765_));
 sky130_fd_sc_hd__o22a_1 _07613_ (.A1(net82),
    .A2(net119),
    .B1(net70),
    .B2(net130),
    .X(_00766_));
 sky130_fd_sc_hd__xnor2_1 _07614_ (.A(net157),
    .B(_00766_),
    .Y(_00767_));
 sky130_fd_sc_hd__nor2_1 _07615_ (.A(_00765_),
    .B(_00767_),
    .Y(_00768_));
 sky130_fd_sc_hd__xnor2_1 _07616_ (.A(_00764_),
    .B(_00767_),
    .Y(_00769_));
 sky130_fd_sc_hd__o22a_1 _07617_ (.A1(net128),
    .A2(net79),
    .B1(net124),
    .B2(net100),
    .X(_00770_));
 sky130_fd_sc_hd__xnor2_1 _07618_ (.A(net154),
    .B(_00770_),
    .Y(_00771_));
 sky130_fd_sc_hd__and2_1 _07619_ (.A(_00769_),
    .B(_00771_),
    .X(_00772_));
 sky130_fd_sc_hd__nor2_1 _07620_ (.A(_00769_),
    .B(_00771_),
    .Y(_00773_));
 sky130_fd_sc_hd__nor2_2 _07621_ (.A(_00772_),
    .B(_00773_),
    .Y(_00774_));
 sky130_fd_sc_hd__nand2_1 _07622_ (.A(_00762_),
    .B(_00774_),
    .Y(_00775_));
 sky130_fd_sc_hd__xnor2_4 _07623_ (.A(_00762_),
    .B(_00774_),
    .Y(_00776_));
 sky130_fd_sc_hd__xnor2_2 _07624_ (.A(_00749_),
    .B(_00776_),
    .Y(_00777_));
 sky130_fd_sc_hd__or2_1 _07625_ (.A(_00738_),
    .B(_00777_),
    .X(_00778_));
 sky130_fd_sc_hd__xnor2_2 _07626_ (.A(_00738_),
    .B(_00777_),
    .Y(_00779_));
 sky130_fd_sc_hd__xnor2_2 _07627_ (.A(_00726_),
    .B(_00779_),
    .Y(_00780_));
 sky130_fd_sc_hd__o22a_1 _07628_ (.A1(net92),
    .A2(net37),
    .B1(net34),
    .B2(net127),
    .X(_00781_));
 sky130_fd_sc_hd__xnor2_1 _07629_ (.A(net136),
    .B(_00781_),
    .Y(_00782_));
 sky130_fd_sc_hd__o22a_1 _07630_ (.A1(net41),
    .A2(net91),
    .B1(net88),
    .B2(net39),
    .X(_00783_));
 sky130_fd_sc_hd__xnor2_1 _07631_ (.A(net103),
    .B(_00783_),
    .Y(_00784_));
 sky130_fd_sc_hd__and2_1 _07632_ (.A(_00782_),
    .B(_00784_),
    .X(_00785_));
 sky130_fd_sc_hd__nor2_1 _07633_ (.A(_00782_),
    .B(_00784_),
    .Y(_00786_));
 sky130_fd_sc_hd__nor2_1 _07634_ (.A(_00785_),
    .B(_00786_),
    .Y(_00787_));
 sky130_fd_sc_hd__mux2_1 _07635_ (.A0(_00426_),
    .A1(net32),
    .S(_00422_),
    .X(_00788_));
 sky130_fd_sc_hd__inv_2 _07636_ (.A(_00788_),
    .Y(_00789_));
 sky130_fd_sc_hd__xnor2_1 _07637_ (.A(_00787_),
    .B(_00788_),
    .Y(_00790_));
 sky130_fd_sc_hd__o21a_1 _07638_ (.A1(_00294_),
    .A2(_00314_),
    .B1(_00790_),
    .X(_00791_));
 sky130_fd_sc_hd__nor3_1 _07639_ (.A(_00294_),
    .B(_00314_),
    .C(_00790_),
    .Y(_00792_));
 sky130_fd_sc_hd__nor2_1 _07640_ (.A(_00791_),
    .B(_00792_),
    .Y(_00793_));
 sky130_fd_sc_hd__xnor2_1 _07641_ (.A(_00780_),
    .B(_00793_),
    .Y(_00794_));
 sky130_fd_sc_hd__nand2_1 _07642_ (.A(_00720_),
    .B(_00794_),
    .Y(_00795_));
 sky130_fd_sc_hd__or2_1 _07643_ (.A(_00720_),
    .B(_00794_),
    .X(_00796_));
 sky130_fd_sc_hd__and2_1 _07644_ (.A(_00795_),
    .B(_00796_),
    .X(_00797_));
 sky130_fd_sc_hd__a21o_1 _07645_ (.A1(_00359_),
    .A2(_00486_),
    .B1(_00484_),
    .X(_00798_));
 sky130_fd_sc_hd__a21bo_1 _07646_ (.A1(_00552_),
    .A2(_00556_),
    .B1_N(_00555_),
    .X(_00799_));
 sky130_fd_sc_hd__a21o_1 _07647_ (.A1(_00316_),
    .A2(_00355_),
    .B1(_00357_),
    .X(_00800_));
 sky130_fd_sc_hd__o32a_1 _07648_ (.A1(_00368_),
    .A2(_00369_),
    .A3(_00428_),
    .B1(_00427_),
    .B2(_00415_),
    .X(_00801_));
 sky130_fd_sc_hd__nor2_1 _07649_ (.A(_00479_),
    .B(_00482_),
    .Y(_00802_));
 sky130_fd_sc_hd__nor2_1 _07650_ (.A(_00801_),
    .B(_00802_),
    .Y(_00803_));
 sky130_fd_sc_hd__xor2_2 _07651_ (.A(_00801_),
    .B(_00802_),
    .X(_00804_));
 sky130_fd_sc_hd__xor2_2 _07652_ (.A(_00800_),
    .B(_00804_),
    .X(_00805_));
 sky130_fd_sc_hd__xnor2_2 _07653_ (.A(_00799_),
    .B(_00805_),
    .Y(_00806_));
 sky130_fd_sc_hd__nand2b_1 _07654_ (.A_N(_00806_),
    .B(_00798_),
    .Y(_00807_));
 sky130_fd_sc_hd__xnor2_2 _07655_ (.A(_00798_),
    .B(_00806_),
    .Y(_00808_));
 sky130_fd_sc_hd__and2_1 _07656_ (.A(_00797_),
    .B(_00808_),
    .X(_00809_));
 sky130_fd_sc_hd__xor2_2 _07657_ (.A(_00797_),
    .B(_00808_),
    .X(_00810_));
 sky130_fd_sc_hd__xnor2_1 _07658_ (.A(_00705_),
    .B(_00810_),
    .Y(_00811_));
 sky130_fd_sc_hd__a21oi_1 _07659_ (.A1(_00629_),
    .A2(_00704_),
    .B1(_00811_),
    .Y(_00812_));
 sky130_fd_sc_hd__and3_1 _07660_ (.A(_00629_),
    .B(_00704_),
    .C(_00811_),
    .X(_00813_));
 sky130_fd_sc_hd__nand3_1 _07661_ (.A(_00692_),
    .B(_00701_),
    .C(_00703_),
    .Y(_00814_));
 sky130_fd_sc_hd__nand2_1 _07662_ (.A(_00704_),
    .B(_00814_),
    .Y(_00815_));
 sky130_fd_sc_hd__xor2_2 _07663_ (.A(_00549_),
    .B(_00550_),
    .X(_00816_));
 sky130_fd_sc_hd__xnor2_2 _07664_ (.A(_00698_),
    .B(_00700_),
    .Y(_00817_));
 sky130_fd_sc_hd__xnor2_1 _07665_ (.A(_00688_),
    .B(_00689_),
    .Y(_00818_));
 sky130_fd_sc_hd__xnor2_2 _07666_ (.A(_00678_),
    .B(_00683_),
    .Y(_00819_));
 sky130_fd_sc_hd__nor2_1 _07667_ (.A(_00637_),
    .B(_00639_),
    .Y(_00820_));
 sky130_fd_sc_hd__nor2_1 _07668_ (.A(_00640_),
    .B(_00820_),
    .Y(_00821_));
 sky130_fd_sc_hd__nand2_1 _07669_ (.A(_00819_),
    .B(_00821_),
    .Y(_00822_));
 sky130_fd_sc_hd__nand2_1 _07670_ (.A(_00670_),
    .B(_00672_),
    .Y(_00823_));
 sky130_fd_sc_hd__nand2_1 _07671_ (.A(_00673_),
    .B(_00823_),
    .Y(_00824_));
 sky130_fd_sc_hd__xnor2_2 _07672_ (.A(_00819_),
    .B(_00821_),
    .Y(_00825_));
 sky130_fd_sc_hd__o21a_1 _07673_ (.A1(_00824_),
    .A2(_00825_),
    .B1(_00822_),
    .X(_00826_));
 sky130_fd_sc_hd__and2_1 _07674_ (.A(_00615_),
    .B(_00617_),
    .X(_00827_));
 sky130_fd_sc_hd__nor2_1 _07675_ (.A(_00618_),
    .B(_00827_),
    .Y(_00828_));
 sky130_fd_sc_hd__o22a_1 _07676_ (.A1(net122),
    .A2(net117),
    .B1(net114),
    .B2(net80),
    .X(_00829_));
 sky130_fd_sc_hd__xnor2_1 _07677_ (.A(net180),
    .B(_00829_),
    .Y(_00830_));
 sky130_fd_sc_hd__o22a_1 _07678_ (.A1(net79),
    .A2(net91),
    .B1(_00457_),
    .B2(net124),
    .X(_00831_));
 sky130_fd_sc_hd__xor2_1 _07679_ (.A(net155),
    .B(_00831_),
    .X(_00832_));
 sky130_fd_sc_hd__nor2_1 _07680_ (.A(_00830_),
    .B(_00832_),
    .Y(_00833_));
 sky130_fd_sc_hd__xnor2_1 _07681_ (.A(_00830_),
    .B(_00832_),
    .Y(_00834_));
 sky130_fd_sc_hd__o22a_1 _07682_ (.A1(net130),
    .A2(net127),
    .B1(net92),
    .B2(net82),
    .X(_00835_));
 sky130_fd_sc_hd__xnor2_1 _07683_ (.A(net158),
    .B(_00835_),
    .Y(_00836_));
 sky130_fd_sc_hd__nor2_1 _07684_ (.A(_00834_),
    .B(_00836_),
    .Y(_00837_));
 sky130_fd_sc_hd__o21a_1 _07685_ (.A1(_00833_),
    .A2(_00837_),
    .B1(_00828_),
    .X(_00838_));
 sky130_fd_sc_hd__o22a_1 _07686_ (.A1(_00136_),
    .A2(net169),
    .B1(net167),
    .B2(net75),
    .X(_00839_));
 sky130_fd_sc_hd__xnor2_1 _07687_ (.A(net210),
    .B(_00839_),
    .Y(_00840_));
 sky130_fd_sc_hd__o22a_1 _07688_ (.A1(net128),
    .A2(net153),
    .B1(_00137_),
    .B2(net101),
    .X(_00841_));
 sky130_fd_sc_hd__xnor2_1 _07689_ (.A(_06489_),
    .B(_00841_),
    .Y(_00842_));
 sky130_fd_sc_hd__o22a_1 _07690_ (.A1(net120),
    .A2(net177),
    .B1(net175),
    .B2(net72),
    .X(_00843_));
 sky130_fd_sc_hd__xnor2_1 _07691_ (.A(net189),
    .B(_00843_),
    .Y(_00844_));
 sky130_fd_sc_hd__xnor2_1 _07692_ (.A(_00840_),
    .B(_00842_),
    .Y(_00845_));
 sky130_fd_sc_hd__nor2_1 _07693_ (.A(_00844_),
    .B(_00845_),
    .Y(_00846_));
 sky130_fd_sc_hd__o21bai_2 _07694_ (.A1(_00840_),
    .A2(_00842_),
    .B1_N(_00846_),
    .Y(_00847_));
 sky130_fd_sc_hd__nor3_1 _07695_ (.A(_00828_),
    .B(_00833_),
    .C(_00837_),
    .Y(_00848_));
 sky130_fd_sc_hd__nor2_1 _07696_ (.A(_00838_),
    .B(_00848_),
    .Y(_00849_));
 sky130_fd_sc_hd__a21o_1 _07697_ (.A1(_00847_),
    .A2(_00849_),
    .B1(_00838_),
    .X(_00850_));
 sky130_fd_sc_hd__nand2b_1 _07698_ (.A_N(_00826_),
    .B(_00850_),
    .Y(_00851_));
 sky130_fd_sc_hd__nand2_1 _07699_ (.A(_00648_),
    .B(_00650_),
    .Y(_00852_));
 sky130_fd_sc_hd__nand2_1 _07700_ (.A(_00651_),
    .B(_00852_),
    .Y(_00853_));
 sky130_fd_sc_hd__o22a_1 _07701_ (.A1(_00290_),
    .A2(net43),
    .B1(net95),
    .B2(net134),
    .X(_00854_));
 sky130_fd_sc_hd__xnor2_1 _07702_ (.A(net138),
    .B(_00854_),
    .Y(_00855_));
 sky130_fd_sc_hd__o22a_1 _07703_ (.A1(net149),
    .A2(net41),
    .B1(net39),
    .B2(net143),
    .X(_00856_));
 sky130_fd_sc_hd__xnor2_1 _07704_ (.A(net103),
    .B(_00856_),
    .Y(_00857_));
 sky130_fd_sc_hd__xor2_1 _07705_ (.A(_00855_),
    .B(_00857_),
    .X(_00858_));
 sky130_fd_sc_hd__o22a_1 _07706_ (.A1(net141),
    .A2(net37),
    .B1(net34),
    .B2(net147),
    .X(_00859_));
 sky130_fd_sc_hd__xnor2_1 _07707_ (.A(net135),
    .B(_00859_),
    .Y(_00860_));
 sky130_fd_sc_hd__and2_1 _07708_ (.A(_00858_),
    .B(_00860_),
    .X(_00861_));
 sky130_fd_sc_hd__a21oi_1 _07709_ (.A1(_00855_),
    .A2(_00857_),
    .B1(_00861_),
    .Y(_00862_));
 sky130_fd_sc_hd__o22a_1 _07710_ (.A1(net75),
    .A2(net173),
    .B1(net171),
    .B2(net69),
    .X(_00863_));
 sky130_fd_sc_hd__xnor2_2 _07711_ (.A(_00180_),
    .B(_00863_),
    .Y(_00864_));
 sky130_fd_sc_hd__o22a_1 _07712_ (.A1(net302),
    .A2(net59),
    .B1(net253),
    .B2(net66),
    .X(_00865_));
 sky130_fd_sc_hd__xnor2_2 _07713_ (.A(net256),
    .B(_00865_),
    .Y(_00866_));
 sky130_fd_sc_hd__and2_1 _07714_ (.A(_00864_),
    .B(_00866_),
    .X(_00867_));
 sky130_fd_sc_hd__o22a_1 _07715_ (.A1(net165),
    .A2(net49),
    .B1(net161),
    .B2(net51),
    .X(_00868_));
 sky130_fd_sc_hd__xnor2_1 _07716_ (.A(net107),
    .B(_00868_),
    .Y(_00869_));
 sky130_fd_sc_hd__and3_1 _07717_ (.A(_00864_),
    .B(_00866_),
    .C(_00869_),
    .X(_00870_));
 sky130_fd_sc_hd__nand3_1 _07718_ (.A(_00864_),
    .B(_00866_),
    .C(_00869_),
    .Y(_00871_));
 sky130_fd_sc_hd__a21o_1 _07719_ (.A1(_00864_),
    .A2(_00866_),
    .B1(_00869_),
    .X(_00872_));
 sky130_fd_sc_hd__a22o_1 _07720_ (.A1(net227),
    .A2(_00307_),
    .B1(_00308_),
    .B2(_00338_),
    .X(_00873_));
 sky130_fd_sc_hd__xor2_1 _07721_ (.A(net110),
    .B(_00873_),
    .X(_00874_));
 sky130_fd_sc_hd__and3_1 _07722_ (.A(_00871_),
    .B(_00872_),
    .C(_00874_),
    .X(_00875_));
 sky130_fd_sc_hd__xor2_1 _07723_ (.A(_00853_),
    .B(_00862_),
    .X(_00876_));
 sky130_fd_sc_hd__o21ai_1 _07724_ (.A1(_00870_),
    .A2(_00875_),
    .B1(_00876_),
    .Y(_00877_));
 sky130_fd_sc_hd__o21ai_2 _07725_ (.A1(_00853_),
    .A2(_00862_),
    .B1(_00877_),
    .Y(_00878_));
 sky130_fd_sc_hd__xnor2_2 _07726_ (.A(_00826_),
    .B(_00850_),
    .Y(_00879_));
 sky130_fd_sc_hd__nand2_1 _07727_ (.A(_00878_),
    .B(_00879_),
    .Y(_00880_));
 sky130_fd_sc_hd__a21o_1 _07728_ (.A1(_00851_),
    .A2(_00880_),
    .B1(_00818_),
    .X(_00881_));
 sky130_fd_sc_hd__xor2_1 _07729_ (.A(_00643_),
    .B(_00652_),
    .X(_00882_));
 sky130_fd_sc_hd__xnor2_1 _07730_ (.A(_00660_),
    .B(_00661_),
    .Y(_00883_));
 sky130_fd_sc_hd__xnor2_1 _07731_ (.A(_00685_),
    .B(_00687_),
    .Y(_00884_));
 sky130_fd_sc_hd__xnor2_1 _07732_ (.A(_00882_),
    .B(_00883_),
    .Y(_00885_));
 sky130_fd_sc_hd__nor2_1 _07733_ (.A(_00884_),
    .B(_00885_),
    .Y(_00886_));
 sky130_fd_sc_hd__o21ba_1 _07734_ (.A1(_00882_),
    .A2(_00883_),
    .B1_N(_00886_),
    .X(_00887_));
 sky130_fd_sc_hd__nand3_1 _07735_ (.A(_00818_),
    .B(_00851_),
    .C(_00880_),
    .Y(_00888_));
 sky130_fd_sc_hd__and2_1 _07736_ (.A(_00881_),
    .B(_00888_),
    .X(_00889_));
 sky130_fd_sc_hd__nand2b_1 _07737_ (.A_N(_00887_),
    .B(_00889_),
    .Y(_00890_));
 sky130_fd_sc_hd__nand2_2 _07738_ (.A(_00881_),
    .B(_00890_),
    .Y(_00891_));
 sky130_fd_sc_hd__xnor2_2 _07739_ (.A(_00816_),
    .B(_00817_),
    .Y(_00892_));
 sky130_fd_sc_hd__and2b_1 _07740_ (.A_N(_00892_),
    .B(_00891_),
    .X(_00893_));
 sky130_fd_sc_hd__a21oi_1 _07741_ (.A1(_00816_),
    .A2(_00817_),
    .B1(_00893_),
    .Y(_00894_));
 sky130_fd_sc_hd__or2_1 _07742_ (.A(_00815_),
    .B(_00894_),
    .X(_00895_));
 sky130_fd_sc_hd__nand2_1 _07743_ (.A(_00815_),
    .B(_00894_),
    .Y(_00896_));
 sky130_fd_sc_hd__and2_2 _07744_ (.A(_00895_),
    .B(_00896_),
    .X(_00897_));
 sky130_fd_sc_hd__nand2_1 _07745_ (.A(_00695_),
    .B(_00696_),
    .Y(_00898_));
 sky130_fd_sc_hd__and2_2 _07746_ (.A(_00697_),
    .B(_00898_),
    .X(_00899_));
 sky130_fd_sc_hd__xnor2_2 _07747_ (.A(_00887_),
    .B(_00889_),
    .Y(_00900_));
 sky130_fd_sc_hd__nand2_1 _07748_ (.A(_00899_),
    .B(_00900_),
    .Y(_00901_));
 sky130_fd_sc_hd__xnor2_2 _07749_ (.A(_00878_),
    .B(_00879_),
    .Y(_00902_));
 sky130_fd_sc_hd__xor2_1 _07750_ (.A(_00834_),
    .B(_00836_),
    .X(_00903_));
 sky130_fd_sc_hd__a21oi_1 _07751_ (.A1(_00871_),
    .A2(_00872_),
    .B1(_00874_),
    .Y(_00904_));
 sky130_fd_sc_hd__or3b_1 _07752_ (.A(_00875_),
    .B(_00904_),
    .C_N(_00903_),
    .X(_00905_));
 sky130_fd_sc_hd__nor2_1 _07753_ (.A(_00858_),
    .B(_00860_),
    .Y(_00906_));
 sky130_fd_sc_hd__nor2_1 _07754_ (.A(_00861_),
    .B(_00906_),
    .Y(_00907_));
 sky130_fd_sc_hd__o21bai_2 _07755_ (.A1(_00875_),
    .A2(_00904_),
    .B1_N(_00903_),
    .Y(_00908_));
 sky130_fd_sc_hd__and3_1 _07756_ (.A(_00905_),
    .B(_00907_),
    .C(_00908_),
    .X(_00909_));
 sky130_fd_sc_hd__a21boi_2 _07757_ (.A1(_00907_),
    .A2(_00908_),
    .B1_N(_00905_),
    .Y(_00910_));
 sky130_fd_sc_hd__and2_1 _07758_ (.A(_00680_),
    .B(_00682_),
    .X(_00911_));
 sky130_fd_sc_hd__nor2_1 _07759_ (.A(_00683_),
    .B(_00911_),
    .Y(_00912_));
 sky130_fd_sc_hd__o22a_1 _07760_ (.A1(net126),
    .A2(net117),
    .B1(_00152_),
    .B2(net121),
    .X(_00913_));
 sky130_fd_sc_hd__xnor2_1 _07761_ (.A(net180),
    .B(_00913_),
    .Y(_00914_));
 sky130_fd_sc_hd__a21o_1 _07762_ (.A1(_06475_),
    .A2(_06477_),
    .B1(net132),
    .X(_00915_));
 sky130_fd_sc_hd__or2_1 _07763_ (.A(net124),
    .B(net90),
    .X(_00916_));
 sky130_fd_sc_hd__nand3_1 _07764_ (.A(net156),
    .B(_00915_),
    .C(_00916_),
    .Y(_00917_));
 sky130_fd_sc_hd__a21o_1 _07765_ (.A1(_00915_),
    .A2(_00916_),
    .B1(net156),
    .X(_00918_));
 sky130_fd_sc_hd__a21oi_1 _07766_ (.A1(_00917_),
    .A2(_00918_),
    .B1(_00914_),
    .Y(_00919_));
 sky130_fd_sc_hd__a21o_1 _07767_ (.A1(_00917_),
    .A2(_00918_),
    .B1(_00914_),
    .X(_00920_));
 sky130_fd_sc_hd__nand3_1 _07768_ (.A(_00914_),
    .B(_00917_),
    .C(_00918_),
    .Y(_00921_));
 sky130_fd_sc_hd__o22a_1 _07769_ (.A1(net130),
    .A2(net92),
    .B1(net87),
    .B2(net82),
    .X(_00922_));
 sky130_fd_sc_hd__xnor2_1 _07770_ (.A(_06435_),
    .B(_00922_),
    .Y(_00923_));
 sky130_fd_sc_hd__and3_1 _07771_ (.A(_00920_),
    .B(_00921_),
    .C(_00923_),
    .X(_00924_));
 sky130_fd_sc_hd__o21a_1 _07772_ (.A1(_00919_),
    .A2(_00924_),
    .B1(_00912_),
    .X(_00925_));
 sky130_fd_sc_hd__o22a_1 _07773_ (.A1(net81),
    .A2(net152),
    .B1(net150),
    .B2(_06468_),
    .X(_00926_));
 sky130_fd_sc_hd__xnor2_2 _07774_ (.A(net191),
    .B(_00926_),
    .Y(_00927_));
 sky130_fd_sc_hd__o22a_1 _07775_ (.A1(net72),
    .A2(net169),
    .B1(net167),
    .B2(net77),
    .X(_00928_));
 sky130_fd_sc_hd__xnor2_2 _07776_ (.A(net211),
    .B(_00928_),
    .Y(_00929_));
 sky130_fd_sc_hd__o22a_1 _07777_ (.A1(net120),
    .A2(net175),
    .B1(net101),
    .B2(net177),
    .X(_00930_));
 sky130_fd_sc_hd__xnor2_1 _07778_ (.A(net189),
    .B(_00930_),
    .Y(_00931_));
 sky130_fd_sc_hd__xnor2_1 _07779_ (.A(_00927_),
    .B(_00929_),
    .Y(_00932_));
 sky130_fd_sc_hd__nor2_1 _07780_ (.A(_00931_),
    .B(_00932_),
    .Y(_00933_));
 sky130_fd_sc_hd__o21bai_2 _07781_ (.A1(_00927_),
    .A2(_00929_),
    .B1_N(_00933_),
    .Y(_00934_));
 sky130_fd_sc_hd__nor3_1 _07782_ (.A(_00912_),
    .B(_00919_),
    .C(_00924_),
    .Y(_00935_));
 sky130_fd_sc_hd__nor2_1 _07783_ (.A(_00925_),
    .B(_00935_),
    .Y(_00936_));
 sky130_fd_sc_hd__a21oi_2 _07784_ (.A1(_00934_),
    .A2(_00936_),
    .B1(_00925_),
    .Y(_00937_));
 sky130_fd_sc_hd__and2_1 _07785_ (.A(_00844_),
    .B(_00845_),
    .X(_00938_));
 sky130_fd_sc_hd__nor2_1 _07786_ (.A(_00846_),
    .B(_00938_),
    .Y(_00939_));
 sky130_fd_sc_hd__o22a_1 _07787_ (.A1(net147),
    .A2(net42),
    .B1(net95),
    .B2(net144),
    .X(_00940_));
 sky130_fd_sc_hd__xnor2_1 _07788_ (.A(net138),
    .B(_00940_),
    .Y(_00941_));
 sky130_fd_sc_hd__o22a_1 _07789_ (.A1(net165),
    .A2(net40),
    .B1(net38),
    .B2(net149),
    .X(_00942_));
 sky130_fd_sc_hd__xnor2_1 _07790_ (.A(net103),
    .B(_00942_),
    .Y(_00943_));
 sky130_fd_sc_hd__and2_1 _07791_ (.A(_00941_),
    .B(_00943_),
    .X(_00944_));
 sky130_fd_sc_hd__xnor2_1 _07792_ (.A(_00941_),
    .B(_00943_),
    .Y(_00945_));
 sky130_fd_sc_hd__o22a_1 _07793_ (.A1(net143),
    .A2(net37),
    .B1(net34),
    .B2(net141),
    .X(_00946_));
 sky130_fd_sc_hd__xnor2_1 _07794_ (.A(_00436_),
    .B(_00946_),
    .Y(_00947_));
 sky130_fd_sc_hd__nor2_1 _07795_ (.A(_00945_),
    .B(_00947_),
    .Y(_00948_));
 sky130_fd_sc_hd__o21a_1 _07796_ (.A1(_00944_),
    .A2(_00948_),
    .B1(_00939_),
    .X(_00949_));
 sky130_fd_sc_hd__nor3_1 _07797_ (.A(_00939_),
    .B(_00944_),
    .C(_00948_),
    .Y(_00950_));
 sky130_fd_sc_hd__nor2_1 _07798_ (.A(_00949_),
    .B(_00950_),
    .Y(_00951_));
 sky130_fd_sc_hd__nand2_1 _07799_ (.A(net227),
    .B(_00308_),
    .Y(_00952_));
 sky130_fd_sc_hd__o22a_1 _07800_ (.A1(net51),
    .A2(net163),
    .B1(net161),
    .B2(net49),
    .X(_00953_));
 sky130_fd_sc_hd__xnor2_1 _07801_ (.A(net107),
    .B(_00953_),
    .Y(_00954_));
 sky130_fd_sc_hd__mux2_1 _07802_ (.A0(_00954_),
    .A1(net110),
    .S(_00952_),
    .X(_00955_));
 sky130_fd_sc_hd__a21o_1 _07803_ (.A1(_00951_),
    .A2(_00955_),
    .B1(_00949_),
    .X(_00956_));
 sky130_fd_sc_hd__xnor2_2 _07804_ (.A(_00910_),
    .B(_00937_),
    .Y(_00957_));
 sky130_fd_sc_hd__nand2b_1 _07805_ (.A_N(_00957_),
    .B(_00956_),
    .Y(_00958_));
 sky130_fd_sc_hd__o21ai_2 _07806_ (.A1(_00910_),
    .A2(_00937_),
    .B1(_00958_),
    .Y(_00959_));
 sky130_fd_sc_hd__nand2b_1 _07807_ (.A_N(_00902_),
    .B(_00959_),
    .Y(_00960_));
 sky130_fd_sc_hd__xor2_2 _07808_ (.A(_00824_),
    .B(_00825_),
    .X(_00961_));
 sky130_fd_sc_hd__inv_2 _07809_ (.A(_00961_),
    .Y(_00962_));
 sky130_fd_sc_hd__xnor2_1 _07810_ (.A(_00847_),
    .B(_00849_),
    .Y(_00963_));
 sky130_fd_sc_hd__or3_1 _07811_ (.A(_00870_),
    .B(_00875_),
    .C(_00876_),
    .X(_00964_));
 sky130_fd_sc_hd__nand2_1 _07812_ (.A(_00877_),
    .B(_00964_),
    .Y(_00965_));
 sky130_fd_sc_hd__xor2_1 _07813_ (.A(_00961_),
    .B(_00963_),
    .X(_00966_));
 sky130_fd_sc_hd__nor2_1 _07814_ (.A(_00965_),
    .B(_00966_),
    .Y(_00967_));
 sky130_fd_sc_hd__o21ba_1 _07815_ (.A1(_00962_),
    .A2(_00963_),
    .B1_N(_00967_),
    .X(_00968_));
 sky130_fd_sc_hd__xnor2_2 _07816_ (.A(_00902_),
    .B(_00959_),
    .Y(_00969_));
 sky130_fd_sc_hd__nand2b_1 _07817_ (.A_N(_00968_),
    .B(_00969_),
    .Y(_00970_));
 sky130_fd_sc_hd__nand2_1 _07818_ (.A(_00960_),
    .B(_00970_),
    .Y(_00971_));
 sky130_fd_sc_hd__xnor2_2 _07819_ (.A(_00899_),
    .B(_00900_),
    .Y(_00972_));
 sky130_fd_sc_hd__nand2b_1 _07820_ (.A_N(_00972_),
    .B(_00971_),
    .Y(_00973_));
 sky130_fd_sc_hd__xor2_2 _07821_ (.A(_00891_),
    .B(_00892_),
    .X(_00974_));
 sky130_fd_sc_hd__a21oi_1 _07822_ (.A1(_00901_),
    .A2(_00973_),
    .B1(_00974_),
    .Y(_00975_));
 sky130_fd_sc_hd__and3_1 _07823_ (.A(_00901_),
    .B(_00973_),
    .C(_00974_),
    .X(_00976_));
 sky130_fd_sc_hd__xor2_2 _07824_ (.A(_00971_),
    .B(_00972_),
    .X(_00977_));
 sky130_fd_sc_hd__and2_1 _07825_ (.A(_00884_),
    .B(_00885_),
    .X(_00978_));
 sky130_fd_sc_hd__nor2_2 _07826_ (.A(_00886_),
    .B(_00978_),
    .Y(_00979_));
 sky130_fd_sc_hd__xnor2_2 _07827_ (.A(_00968_),
    .B(_00969_),
    .Y(_00980_));
 sky130_fd_sc_hd__xor2_2 _07828_ (.A(_00956_),
    .B(_00957_),
    .X(_00981_));
 sky130_fd_sc_hd__nor2_1 _07829_ (.A(_00864_),
    .B(_00866_),
    .Y(_00982_));
 sky130_fd_sc_hd__xor2_1 _07830_ (.A(_00864_),
    .B(_00866_),
    .X(_00983_));
 sky130_fd_sc_hd__o22a_1 _07831_ (.A1(net127),
    .A2(net114),
    .B1(net93),
    .B2(net116),
    .X(_00984_));
 sky130_fd_sc_hd__xnor2_1 _07832_ (.A(net180),
    .B(_00984_),
    .Y(_00985_));
 sky130_fd_sc_hd__o22a_1 _07833_ (.A1(net128),
    .A2(net177),
    .B1(net175),
    .B2(net101),
    .X(_00986_));
 sky130_fd_sc_hd__xnor2_1 _07834_ (.A(net189),
    .B(_00986_),
    .Y(_00987_));
 sky130_fd_sc_hd__or2_1 _07835_ (.A(_00985_),
    .B(_00987_),
    .X(_00988_));
 sky130_fd_sc_hd__o22a_1 _07836_ (.A1(net122),
    .A2(net152),
    .B1(net150),
    .B2(net80),
    .X(_00989_));
 sky130_fd_sc_hd__xnor2_1 _07837_ (.A(net191),
    .B(_00989_),
    .Y(_00990_));
 sky130_fd_sc_hd__and2_1 _07838_ (.A(_00985_),
    .B(_00987_),
    .X(_00991_));
 sky130_fd_sc_hd__xor2_1 _07839_ (.A(_00985_),
    .B(_00987_),
    .X(_00992_));
 sky130_fd_sc_hd__o21a_1 _07840_ (.A1(_00990_),
    .A2(_00991_),
    .B1(_00988_),
    .X(_00993_));
 sky130_fd_sc_hd__o22a_1 _07841_ (.A1(net302),
    .A2(net66),
    .B1(net253),
    .B2(net69),
    .X(_00994_));
 sky130_fd_sc_hd__xnor2_1 _07842_ (.A(_00188_),
    .B(_00994_),
    .Y(_00995_));
 sky130_fd_sc_hd__o22a_1 _07843_ (.A1(net120),
    .A2(net169),
    .B1(net167),
    .B2(net72),
    .X(_00996_));
 sky130_fd_sc_hd__xnor2_1 _07844_ (.A(net210),
    .B(_00996_),
    .Y(_00997_));
 sky130_fd_sc_hd__nor2_1 _07845_ (.A(_00995_),
    .B(_00997_),
    .Y(_00998_));
 sky130_fd_sc_hd__o22a_1 _07846_ (.A1(net77),
    .A2(_00193_),
    .B1(_00194_),
    .B2(net75),
    .X(_00999_));
 sky130_fd_sc_hd__xnor2_1 _07847_ (.A(_00179_),
    .B(_00999_),
    .Y(_01000_));
 sky130_fd_sc_hd__xnor2_1 _07848_ (.A(_00995_),
    .B(_00997_),
    .Y(_01001_));
 sky130_fd_sc_hd__nor2_1 _07849_ (.A(_01000_),
    .B(_01001_),
    .Y(_01002_));
 sky130_fd_sc_hd__xnor2_1 _07850_ (.A(_00983_),
    .B(_00993_),
    .Y(_01003_));
 sky130_fd_sc_hd__o21ai_1 _07851_ (.A1(_00998_),
    .A2(_01002_),
    .B1(_01003_),
    .Y(_01004_));
 sky130_fd_sc_hd__o31a_1 _07852_ (.A1(_00867_),
    .A2(_00982_),
    .A3(_00993_),
    .B1(_01004_),
    .X(_01005_));
 sky130_fd_sc_hd__a21oi_1 _07853_ (.A1(_00920_),
    .A2(_00921_),
    .B1(_00923_),
    .Y(_01006_));
 sky130_fd_sc_hd__or2_1 _07854_ (.A(_00924_),
    .B(_01006_),
    .X(_01007_));
 sky130_fd_sc_hd__xor2_1 _07855_ (.A(_00952_),
    .B(_00954_),
    .X(_01008_));
 sky130_fd_sc_hd__nor2_1 _07856_ (.A(_01007_),
    .B(_01008_),
    .Y(_01009_));
 sky130_fd_sc_hd__and2_1 _07857_ (.A(_00945_),
    .B(_00947_),
    .X(_01010_));
 sky130_fd_sc_hd__nor2_1 _07858_ (.A(_00948_),
    .B(_01010_),
    .Y(_01011_));
 sky130_fd_sc_hd__xor2_1 _07859_ (.A(_01007_),
    .B(_01008_),
    .X(_01012_));
 sky130_fd_sc_hd__a21oi_1 _07860_ (.A1(_01011_),
    .A2(_01012_),
    .B1(_01009_),
    .Y(_01013_));
 sky130_fd_sc_hd__and2_1 _07861_ (.A(_00931_),
    .B(_00932_),
    .X(_01014_));
 sky130_fd_sc_hd__nor2_1 _07862_ (.A(_00933_),
    .B(_01014_),
    .Y(_01015_));
 sky130_fd_sc_hd__o22a_1 _07863_ (.A1(net82),
    .A2(net91),
    .B1(net88),
    .B2(_06460_),
    .X(_01016_));
 sky130_fd_sc_hd__xnor2_1 _07864_ (.A(net158),
    .B(_01016_),
    .Y(_01017_));
 sky130_fd_sc_hd__o22a_1 _07865_ (.A1(net141),
    .A2(net43),
    .B1(net94),
    .B2(net147),
    .X(_01018_));
 sky130_fd_sc_hd__xor2_1 _07866_ (.A(net139),
    .B(_01018_),
    .X(_01019_));
 sky130_fd_sc_hd__or2_1 _07867_ (.A(_01017_),
    .B(_01019_),
    .X(_01020_));
 sky130_fd_sc_hd__xnor2_1 _07868_ (.A(_01017_),
    .B(_01019_),
    .Y(_01021_));
 sky130_fd_sc_hd__o22a_1 _07869_ (.A1(net79),
    .A2(net144),
    .B1(net134),
    .B2(_06482_),
    .X(_01022_));
 sky130_fd_sc_hd__xor2_1 _07870_ (.A(net155),
    .B(_01022_),
    .X(_01023_));
 sky130_fd_sc_hd__o21ai_2 _07871_ (.A1(_01021_),
    .A2(_01023_),
    .B1(_01020_),
    .Y(_01024_));
 sky130_fd_sc_hd__o22a_1 _07872_ (.A1(net149),
    .A2(net37),
    .B1(net35),
    .B2(net143),
    .X(_01025_));
 sky130_fd_sc_hd__xnor2_2 _07873_ (.A(net135),
    .B(_01025_),
    .Y(_01026_));
 sky130_fd_sc_hd__o22a_1 _07874_ (.A1(net161),
    .A2(net41),
    .B1(net39),
    .B2(net165),
    .X(_01027_));
 sky130_fd_sc_hd__xnor2_2 _07875_ (.A(net103),
    .B(_01027_),
    .Y(_01028_));
 sky130_fd_sc_hd__nand2_1 _07876_ (.A(_01026_),
    .B(_01028_),
    .Y(_01029_));
 sky130_fd_sc_hd__xor2_1 _07877_ (.A(_01015_),
    .B(_01024_),
    .X(_01030_));
 sky130_fd_sc_hd__a32o_1 _07878_ (.A1(_01026_),
    .A2(_01028_),
    .A3(_01030_),
    .B1(_01024_),
    .B2(_01015_),
    .X(_01031_));
 sky130_fd_sc_hd__xnor2_1 _07879_ (.A(_01005_),
    .B(_01013_),
    .Y(_01032_));
 sky130_fd_sc_hd__nand2b_1 _07880_ (.A_N(_01032_),
    .B(_01031_),
    .Y(_01033_));
 sky130_fd_sc_hd__o21a_1 _07881_ (.A1(_01005_),
    .A2(_01013_),
    .B1(_01033_),
    .X(_01034_));
 sky130_fd_sc_hd__a21oi_1 _07882_ (.A1(_00905_),
    .A2(_00908_),
    .B1(_00907_),
    .Y(_01035_));
 sky130_fd_sc_hd__or2_1 _07883_ (.A(_00909_),
    .B(_01035_),
    .X(_01036_));
 sky130_fd_sc_hd__xnor2_2 _07884_ (.A(_00934_),
    .B(_00936_),
    .Y(_01037_));
 sky130_fd_sc_hd__xnor2_1 _07885_ (.A(_00951_),
    .B(_00955_),
    .Y(_01038_));
 sky130_fd_sc_hd__xnor2_1 _07886_ (.A(_01036_),
    .B(_01037_),
    .Y(_01039_));
 sky130_fd_sc_hd__or2_1 _07887_ (.A(_01038_),
    .B(_01039_),
    .X(_01040_));
 sky130_fd_sc_hd__o21ai_2 _07888_ (.A1(_01036_),
    .A2(_01037_),
    .B1(_01040_),
    .Y(_01041_));
 sky130_fd_sc_hd__xnor2_2 _07889_ (.A(_00981_),
    .B(_01034_),
    .Y(_01042_));
 sky130_fd_sc_hd__nand2b_1 _07890_ (.A_N(_01042_),
    .B(_01041_),
    .Y(_01043_));
 sky130_fd_sc_hd__o21ai_2 _07891_ (.A1(_00981_),
    .A2(_01034_),
    .B1(_01043_),
    .Y(_01044_));
 sky130_fd_sc_hd__xnor2_2 _07892_ (.A(_00979_),
    .B(_00980_),
    .Y(_01045_));
 sky130_fd_sc_hd__and2b_1 _07893_ (.A_N(_01045_),
    .B(_01044_),
    .X(_01046_));
 sky130_fd_sc_hd__a21oi_1 _07894_ (.A1(_00979_),
    .A2(_00980_),
    .B1(_01046_),
    .Y(_01047_));
 sky130_fd_sc_hd__or2_1 _07895_ (.A(_00977_),
    .B(_01047_),
    .X(_01048_));
 sky130_fd_sc_hd__xnor2_2 _07896_ (.A(_00977_),
    .B(_01047_),
    .Y(_01049_));
 sky130_fd_sc_hd__inv_2 _07897_ (.A(_01049_),
    .Y(_01050_));
 sky130_fd_sc_hd__and2_1 _07898_ (.A(_00965_),
    .B(_00966_),
    .X(_01051_));
 sky130_fd_sc_hd__nor2_1 _07899_ (.A(_00967_),
    .B(_01051_),
    .Y(_01052_));
 sky130_fd_sc_hd__xnor2_2 _07900_ (.A(_01041_),
    .B(_01042_),
    .Y(_01053_));
 sky130_fd_sc_hd__nand2_1 _07901_ (.A(_01052_),
    .B(_01053_),
    .Y(_01054_));
 sky130_fd_sc_hd__xor2_2 _07902_ (.A(_01031_),
    .B(_01032_),
    .X(_01055_));
 sky130_fd_sc_hd__o22a_1 _07903_ (.A1(net115),
    .A2(net93),
    .B1(net88),
    .B2(net117),
    .X(_01056_));
 sky130_fd_sc_hd__xor2_1 _07904_ (.A(net181),
    .B(_01056_),
    .X(_01057_));
 sky130_fd_sc_hd__a21o_1 _07905_ (.A1(_06456_),
    .A2(_06457_),
    .B1(net176),
    .X(_01058_));
 sky130_fd_sc_hd__or2_1 _07906_ (.A(net129),
    .B(net174),
    .X(_01059_));
 sky130_fd_sc_hd__a21o_1 _07907_ (.A1(_01058_),
    .A2(_01059_),
    .B1(net188),
    .X(_01060_));
 sky130_fd_sc_hd__nand3_1 _07908_ (.A(net188),
    .B(_01058_),
    .C(_01059_),
    .Y(_01061_));
 sky130_fd_sc_hd__nand3_2 _07909_ (.A(_01057_),
    .B(_01060_),
    .C(_01061_),
    .Y(_01062_));
 sky130_fd_sc_hd__o22a_1 _07910_ (.A1(net125),
    .A2(net153),
    .B1(net151),
    .B2(net122),
    .X(_01063_));
 sky130_fd_sc_hd__xnor2_2 _07911_ (.A(_06490_),
    .B(_01063_),
    .Y(_01064_));
 sky130_fd_sc_hd__a21o_1 _07912_ (.A1(_01060_),
    .A2(_01061_),
    .B1(_01057_),
    .X(_01065_));
 sky130_fd_sc_hd__nand3_2 _07913_ (.A(_01062_),
    .B(_01064_),
    .C(_01065_),
    .Y(_01066_));
 sky130_fd_sc_hd__a21bo_1 _07914_ (.A1(_01064_),
    .A2(_01065_),
    .B1_N(_01062_),
    .X(_01067_));
 sky130_fd_sc_hd__o22a_1 _07915_ (.A1(net226),
    .A2(net51),
    .B1(net49),
    .B2(net162),
    .X(_01068_));
 sky130_fd_sc_hd__xor2_1 _07916_ (.A(net107),
    .B(_01068_),
    .X(_01069_));
 sky130_fd_sc_hd__a21o_1 _07917_ (.A1(_01062_),
    .A2(_01066_),
    .B1(_01069_),
    .X(_01070_));
 sky130_fd_sc_hd__o22a_1 _07918_ (.A1(net301),
    .A2(net67),
    .B1(net253),
    .B2(net73),
    .X(_01071_));
 sky130_fd_sc_hd__xnor2_1 _07919_ (.A(net255),
    .B(_01071_),
    .Y(_01072_));
 sky130_fd_sc_hd__o22a_1 _07920_ (.A1(net118),
    .A2(net166),
    .B1(net99),
    .B2(net168),
    .X(_01073_));
 sky130_fd_sc_hd__xnor2_1 _07921_ (.A(net209),
    .B(_01073_),
    .Y(_01074_));
 sky130_fd_sc_hd__nor2_1 _07922_ (.A(_01072_),
    .B(_01074_),
    .Y(_01075_));
 sky130_fd_sc_hd__o22a_1 _07923_ (.A1(net70),
    .A2(net173),
    .B1(net170),
    .B2(net76),
    .X(_01076_));
 sky130_fd_sc_hd__xnor2_1 _07924_ (.A(net207),
    .B(_01076_),
    .Y(_01077_));
 sky130_fd_sc_hd__xor2_1 _07925_ (.A(_01072_),
    .B(_01074_),
    .X(_01078_));
 sky130_fd_sc_hd__and2b_1 _07926_ (.A_N(_01077_),
    .B(_01078_),
    .X(_01079_));
 sky130_fd_sc_hd__xnor2_1 _07927_ (.A(_01067_),
    .B(_01069_),
    .Y(_01080_));
 sky130_fd_sc_hd__o21ai_1 _07928_ (.A1(_01075_),
    .A2(_01079_),
    .B1(_01080_),
    .Y(_01081_));
 sky130_fd_sc_hd__xnor2_1 _07929_ (.A(_00990_),
    .B(_00992_),
    .Y(_01082_));
 sky130_fd_sc_hd__xor2_1 _07930_ (.A(_01026_),
    .B(_01028_),
    .X(_01083_));
 sky130_fd_sc_hd__nand2_1 _07931_ (.A(_01082_),
    .B(_01083_),
    .Y(_01084_));
 sky130_fd_sc_hd__xnor2_1 _07932_ (.A(_01021_),
    .B(_01023_),
    .Y(_01085_));
 sky130_fd_sc_hd__xnor2_1 _07933_ (.A(_01082_),
    .B(_01083_),
    .Y(_01086_));
 sky130_fd_sc_hd__o21a_1 _07934_ (.A1(_01085_),
    .A2(_01086_),
    .B1(_01084_),
    .X(_01087_));
 sky130_fd_sc_hd__a21oi_1 _07935_ (.A1(_01070_),
    .A2(_01081_),
    .B1(_01087_),
    .Y(_01088_));
 sky130_fd_sc_hd__o22a_1 _07936_ (.A1(net143),
    .A2(net43),
    .B1(net95),
    .B2(net141),
    .X(_01089_));
 sky130_fd_sc_hd__xor2_2 _07937_ (.A(net139),
    .B(_01089_),
    .X(_01090_));
 sky130_fd_sc_hd__o22a_1 _07938_ (.A1(net83),
    .A2(net132),
    .B1(net89),
    .B2(net131),
    .X(_01091_));
 sky130_fd_sc_hd__xnor2_1 _07939_ (.A(net159),
    .B(_01091_),
    .Y(_01092_));
 sky130_fd_sc_hd__nor2_1 _07940_ (.A(_01090_),
    .B(_01092_),
    .Y(_01093_));
 sky130_fd_sc_hd__nand2_1 _07941_ (.A(_01090_),
    .B(_01092_),
    .Y(_01094_));
 sky130_fd_sc_hd__xnor2_1 _07942_ (.A(_01090_),
    .B(_01092_),
    .Y(_01095_));
 sky130_fd_sc_hd__o22a_1 _07943_ (.A1(net79),
    .A2(net146),
    .B1(net145),
    .B2(net124),
    .X(_01096_));
 sky130_fd_sc_hd__xnor2_1 _07944_ (.A(net156),
    .B(_01096_),
    .Y(_01097_));
 sky130_fd_sc_hd__a21o_1 _07945_ (.A1(_01094_),
    .A2(_01097_),
    .B1(_01093_),
    .X(_01098_));
 sky130_fd_sc_hd__and2_1 _07946_ (.A(_01000_),
    .B(_01001_),
    .X(_01099_));
 sky130_fd_sc_hd__nor2_2 _07947_ (.A(_01002_),
    .B(_01099_),
    .Y(_01100_));
 sky130_fd_sc_hd__o22a_1 _07948_ (.A1(net165),
    .A2(net37),
    .B1(net35),
    .B2(net149),
    .X(_01101_));
 sky130_fd_sc_hd__xnor2_2 _07949_ (.A(net136),
    .B(_01101_),
    .Y(_01102_));
 sky130_fd_sc_hd__o22a_1 _07950_ (.A1(net162),
    .A2(net41),
    .B1(net39),
    .B2(net161),
    .X(_01103_));
 sky130_fd_sc_hd__xnor2_2 _07951_ (.A(net104),
    .B(_01103_),
    .Y(_01104_));
 sky130_fd_sc_hd__nand2_1 _07952_ (.A(_01102_),
    .B(_01104_),
    .Y(_01105_));
 sky130_fd_sc_hd__xor2_2 _07953_ (.A(_01098_),
    .B(_01100_),
    .X(_01106_));
 sky130_fd_sc_hd__a32o_1 _07954_ (.A1(_01102_),
    .A2(_01104_),
    .A3(_01106_),
    .B1(_01100_),
    .B2(_01098_),
    .X(_01107_));
 sky130_fd_sc_hd__and3_1 _07955_ (.A(_01070_),
    .B(_01081_),
    .C(_01087_),
    .X(_01108_));
 sky130_fd_sc_hd__nor2_1 _07956_ (.A(_01088_),
    .B(_01108_),
    .Y(_01109_));
 sky130_fd_sc_hd__a21oi_2 _07957_ (.A1(_01107_),
    .A2(_01109_),
    .B1(_01088_),
    .Y(_01110_));
 sky130_fd_sc_hd__nor2_1 _07958_ (.A(_01055_),
    .B(_01110_),
    .Y(_01111_));
 sky130_fd_sc_hd__or3_1 _07959_ (.A(_00998_),
    .B(_01002_),
    .C(_01003_),
    .X(_01112_));
 sky130_fd_sc_hd__nand2_1 _07960_ (.A(_01004_),
    .B(_01112_),
    .Y(_01113_));
 sky130_fd_sc_hd__xnor2_1 _07961_ (.A(_01011_),
    .B(_01012_),
    .Y(_01114_));
 sky130_fd_sc_hd__or2_1 _07962_ (.A(_01113_),
    .B(_01114_),
    .X(_01115_));
 sky130_fd_sc_hd__xnor2_1 _07963_ (.A(_01029_),
    .B(_01030_),
    .Y(_01116_));
 sky130_fd_sc_hd__nand2_1 _07964_ (.A(_01113_),
    .B(_01114_),
    .Y(_01117_));
 sky130_fd_sc_hd__and3_1 _07965_ (.A(_01115_),
    .B(_01116_),
    .C(_01117_),
    .X(_01118_));
 sky130_fd_sc_hd__a21bo_1 _07966_ (.A1(_01116_),
    .A2(_01117_),
    .B1_N(_01115_),
    .X(_01119_));
 sky130_fd_sc_hd__xor2_1 _07967_ (.A(_01055_),
    .B(_01110_),
    .X(_01120_));
 sky130_fd_sc_hd__a21o_1 _07968_ (.A1(_01119_),
    .A2(_01120_),
    .B1(_01111_),
    .X(_01121_));
 sky130_fd_sc_hd__xnor2_1 _07969_ (.A(_01052_),
    .B(_01053_),
    .Y(_01122_));
 sky130_fd_sc_hd__nand2b_1 _07970_ (.A_N(_01122_),
    .B(_01121_),
    .Y(_01123_));
 sky130_fd_sc_hd__nand2_1 _07971_ (.A(_01054_),
    .B(_01123_),
    .Y(_01124_));
 sky130_fd_sc_hd__xor2_2 _07972_ (.A(_01044_),
    .B(_01045_),
    .X(_01125_));
 sky130_fd_sc_hd__and2b_1 _07973_ (.A_N(_01125_),
    .B(_01124_),
    .X(_01126_));
 sky130_fd_sc_hd__and3_1 _07974_ (.A(_01054_),
    .B(_01123_),
    .C(_01125_),
    .X(_01127_));
 sky130_fd_sc_hd__xor2_2 _07975_ (.A(_01124_),
    .B(_01125_),
    .X(_01128_));
 sky130_fd_sc_hd__xor2_1 _07976_ (.A(_01119_),
    .B(_01120_),
    .X(_01129_));
 sky130_fd_sc_hd__inv_2 _07977_ (.A(_01129_),
    .Y(_01130_));
 sky130_fd_sc_hd__nand2_1 _07978_ (.A(_01038_),
    .B(_01039_),
    .Y(_01131_));
 sky130_fd_sc_hd__nand2_1 _07979_ (.A(_01040_),
    .B(_01131_),
    .Y(_01132_));
 sky130_fd_sc_hd__nor2_1 _07980_ (.A(_01130_),
    .B(_01132_),
    .Y(_01133_));
 sky130_fd_sc_hd__xor2_2 _07981_ (.A(_01107_),
    .B(_01109_),
    .X(_01134_));
 sky130_fd_sc_hd__xor2_1 _07982_ (.A(_01102_),
    .B(_01104_),
    .X(_01135_));
 sky130_fd_sc_hd__a21o_1 _07983_ (.A1(_01062_),
    .A2(_01065_),
    .B1(_01064_),
    .X(_01136_));
 sky130_fd_sc_hd__nand3_2 _07984_ (.A(_01066_),
    .B(_01135_),
    .C(_01136_),
    .Y(_01137_));
 sky130_fd_sc_hd__xnor2_1 _07985_ (.A(_01095_),
    .B(_01097_),
    .Y(_01138_));
 sky130_fd_sc_hd__a21o_1 _07986_ (.A1(_01066_),
    .A2(_01136_),
    .B1(_01135_),
    .X(_01139_));
 sky130_fd_sc_hd__nand3_1 _07987_ (.A(_01137_),
    .B(_01138_),
    .C(_01139_),
    .Y(_01140_));
 sky130_fd_sc_hd__nor2_1 _07988_ (.A(net223),
    .B(net48),
    .Y(_01141_));
 sky130_fd_sc_hd__o22a_2 _07989_ (.A1(net301),
    .A2(net73),
    .B1(net252),
    .B2(net76),
    .X(_01142_));
 sky130_fd_sc_hd__xnor2_4 _07990_ (.A(net254),
    .B(_01142_),
    .Y(_01143_));
 sky130_fd_sc_hd__o22a_2 _07991_ (.A1(net129),
    .A2(net168),
    .B1(net166),
    .B2(net99),
    .X(_01144_));
 sky130_fd_sc_hd__xnor2_4 _07992_ (.A(net209),
    .B(_01144_),
    .Y(_01145_));
 sky130_fd_sc_hd__nor2_1 _07993_ (.A(_01143_),
    .B(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hd__o22a_1 _07994_ (.A1(net118),
    .A2(net172),
    .B1(net170),
    .B2(net70),
    .X(_01147_));
 sky130_fd_sc_hd__xnor2_1 _07995_ (.A(net207),
    .B(_01147_),
    .Y(_01148_));
 sky130_fd_sc_hd__inv_2 _07996_ (.A(_01148_),
    .Y(_01149_));
 sky130_fd_sc_hd__xor2_4 _07997_ (.A(_01143_),
    .B(_01145_),
    .X(_01150_));
 sky130_fd_sc_hd__a21oi_1 _07998_ (.A1(_01149_),
    .A2(_01150_),
    .B1(_01146_),
    .Y(_01151_));
 sky130_fd_sc_hd__nor2_1 _07999_ (.A(net105),
    .B(_01141_),
    .Y(_01152_));
 sky130_fd_sc_hd__a21o_1 _08000_ (.A1(_01141_),
    .A2(_01151_),
    .B1(_01152_),
    .X(_01153_));
 sky130_fd_sc_hd__a21oi_1 _08001_ (.A1(_01137_),
    .A2(_01140_),
    .B1(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__o22a_2 _08002_ (.A1(net117),
    .A2(net89),
    .B1(net87),
    .B2(net115),
    .X(_01155_));
 sky130_fd_sc_hd__xnor2_4 _08003_ (.A(net181),
    .B(_01155_),
    .Y(_01156_));
 sky130_fd_sc_hd__o22a_2 _08004_ (.A1(net122),
    .A2(net176),
    .B1(net174),
    .B2(net81),
    .X(_01157_));
 sky130_fd_sc_hd__xnor2_4 _08005_ (.A(net188),
    .B(_01157_),
    .Y(_01158_));
 sky130_fd_sc_hd__nor2_1 _08006_ (.A(_01156_),
    .B(_01158_),
    .Y(_01159_));
 sky130_fd_sc_hd__o22a_1 _08007_ (.A1(net125),
    .A2(net151),
    .B1(net93),
    .B2(net153),
    .X(_01160_));
 sky130_fd_sc_hd__xnor2_1 _08008_ (.A(net192),
    .B(_01160_),
    .Y(_01161_));
 sky130_fd_sc_hd__inv_2 _08009_ (.A(_01161_),
    .Y(_01162_));
 sky130_fd_sc_hd__xor2_4 _08010_ (.A(_01156_),
    .B(_01158_),
    .X(_01163_));
 sky130_fd_sc_hd__a21o_1 _08011_ (.A1(_01162_),
    .A2(_01163_),
    .B1(_01159_),
    .X(_01164_));
 sky130_fd_sc_hd__xor2_1 _08012_ (.A(_01077_),
    .B(_01078_),
    .X(_01165_));
 sky130_fd_sc_hd__nand2b_1 _08013_ (.A_N(_01165_),
    .B(_01164_),
    .Y(_01166_));
 sky130_fd_sc_hd__o22a_1 _08014_ (.A1(net83),
    .A2(net145),
    .B1(net132),
    .B2(net131),
    .X(_01167_));
 sky130_fd_sc_hd__xnor2_1 _08015_ (.A(net159),
    .B(_01167_),
    .Y(_01168_));
 sky130_fd_sc_hd__o22a_1 _08016_ (.A1(net124),
    .A2(net146),
    .B1(net140),
    .B2(net79),
    .X(_01169_));
 sky130_fd_sc_hd__xor2_1 _08017_ (.A(net156),
    .B(_01169_),
    .X(_01170_));
 sky130_fd_sc_hd__nor2_1 _08018_ (.A(_01168_),
    .B(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hd__xnor2_1 _08019_ (.A(_01164_),
    .B(_01165_),
    .Y(_01172_));
 sky130_fd_sc_hd__nand2_1 _08020_ (.A(_01171_),
    .B(_01172_),
    .Y(_01173_));
 sky130_fd_sc_hd__nand2_1 _08021_ (.A(_01166_),
    .B(_01173_),
    .Y(_01174_));
 sky130_fd_sc_hd__and3_1 _08022_ (.A(_01137_),
    .B(_01140_),
    .C(_01153_),
    .X(_01175_));
 sky130_fd_sc_hd__nor2_1 _08023_ (.A(_01154_),
    .B(_01175_),
    .Y(_01176_));
 sky130_fd_sc_hd__a21oi_2 _08024_ (.A1(_01174_),
    .A2(_01176_),
    .B1(_01154_),
    .Y(_01177_));
 sky130_fd_sc_hd__nand2b_1 _08025_ (.A_N(_01177_),
    .B(_01134_),
    .Y(_01178_));
 sky130_fd_sc_hd__or3_1 _08026_ (.A(_01075_),
    .B(_01079_),
    .C(_01080_),
    .X(_01179_));
 sky130_fd_sc_hd__nand2_1 _08027_ (.A(_01081_),
    .B(_01179_),
    .Y(_01180_));
 sky130_fd_sc_hd__xnor2_1 _08028_ (.A(_01085_),
    .B(_01086_),
    .Y(_01181_));
 sky130_fd_sc_hd__nor2_1 _08029_ (.A(_01180_),
    .B(_01181_),
    .Y(_01182_));
 sky130_fd_sc_hd__xnor2_2 _08030_ (.A(_01105_),
    .B(_01106_),
    .Y(_01183_));
 sky130_fd_sc_hd__nand2_1 _08031_ (.A(_01180_),
    .B(_01181_),
    .Y(_01184_));
 sky130_fd_sc_hd__and2b_1 _08032_ (.A_N(_01182_),
    .B(_01184_),
    .X(_01185_));
 sky130_fd_sc_hd__a21o_1 _08033_ (.A1(_01183_),
    .A2(_01184_),
    .B1(_01182_),
    .X(_01186_));
 sky130_fd_sc_hd__xor2_2 _08034_ (.A(_01134_),
    .B(_01177_),
    .X(_01187_));
 sky130_fd_sc_hd__nand2b_1 _08035_ (.A_N(_01187_),
    .B(_01186_),
    .Y(_01188_));
 sky130_fd_sc_hd__nand2_1 _08036_ (.A(_01178_),
    .B(_01188_),
    .Y(_01189_));
 sky130_fd_sc_hd__xnor2_1 _08037_ (.A(_01129_),
    .B(_01132_),
    .Y(_01190_));
 sky130_fd_sc_hd__and2_1 _08038_ (.A(_01189_),
    .B(_01190_),
    .X(_01191_));
 sky130_fd_sc_hd__xnor2_1 _08039_ (.A(_01121_),
    .B(_01122_),
    .Y(_01192_));
 sky130_fd_sc_hd__o21a_1 _08040_ (.A1(_01133_),
    .A2(_01191_),
    .B1(_01192_),
    .X(_01193_));
 sky130_fd_sc_hd__inv_2 _08041_ (.A(_01193_),
    .Y(_01194_));
 sky130_fd_sc_hd__nor3_1 _08042_ (.A(_01133_),
    .B(_01191_),
    .C(_01192_),
    .Y(_01195_));
 sky130_fd_sc_hd__or2_2 _08043_ (.A(_01193_),
    .B(_01195_),
    .X(_01196_));
 sky130_fd_sc_hd__inv_2 _08044_ (.A(_01196_),
    .Y(_01197_));
 sky130_fd_sc_hd__nor2_1 _08045_ (.A(_01128_),
    .B(_01196_),
    .Y(_01198_));
 sky130_fd_sc_hd__o22a_1 _08046_ (.A1(net117),
    .A2(net145),
    .B1(net132),
    .B2(net115),
    .X(_01199_));
 sky130_fd_sc_hd__xnor2_1 _08047_ (.A(net181),
    .B(_01199_),
    .Y(_01200_));
 sky130_fd_sc_hd__o22a_1 _08048_ (.A1(net79),
    .A2(net148),
    .B1(net142),
    .B2(net124),
    .X(_01201_));
 sky130_fd_sc_hd__xor2_1 _08049_ (.A(net156),
    .B(_01201_),
    .X(_01202_));
 sky130_fd_sc_hd__xnor2_1 _08050_ (.A(_01200_),
    .B(_01202_),
    .Y(_01203_));
 sky130_fd_sc_hd__o22a_1 _08051_ (.A1(net131),
    .A2(net146),
    .B1(net140),
    .B2(net83),
    .X(_01204_));
 sky130_fd_sc_hd__xnor2_1 _08052_ (.A(net159),
    .B(_01204_),
    .Y(_01205_));
 sky130_fd_sc_hd__nor2_1 _08053_ (.A(_01203_),
    .B(_01205_),
    .Y(_01206_));
 sky130_fd_sc_hd__o21bai_1 _08054_ (.A1(_01200_),
    .A2(_01202_),
    .B1_N(_01206_),
    .Y(_01207_));
 sky130_fd_sc_hd__o22a_1 _08055_ (.A1(net153),
    .A2(net132),
    .B1(net89),
    .B2(net151),
    .X(_01208_));
 sky130_fd_sc_hd__xnor2_1 _08056_ (.A(net192),
    .B(_01208_),
    .Y(_01209_));
 sky130_fd_sc_hd__o22a_1 _08057_ (.A1(net174),
    .A2(net93),
    .B1(net87),
    .B2(net176),
    .X(_01210_));
 sky130_fd_sc_hd__xnor2_1 _08058_ (.A(net188),
    .B(_01210_),
    .Y(_01211_));
 sky130_fd_sc_hd__nor2_1 _08059_ (.A(_01209_),
    .B(_01211_),
    .Y(_01212_));
 sky130_fd_sc_hd__o22a_1 _08060_ (.A1(net153),
    .A2(net89),
    .B1(net87),
    .B2(net151),
    .X(_01213_));
 sky130_fd_sc_hd__xnor2_1 _08061_ (.A(net192),
    .B(_01213_),
    .Y(_01214_));
 sky130_fd_sc_hd__o22a_1 _08062_ (.A1(net125),
    .A2(net174),
    .B1(net93),
    .B2(net176),
    .X(_01215_));
 sky130_fd_sc_hd__xnor2_1 _08063_ (.A(net188),
    .B(_01215_),
    .Y(_01216_));
 sky130_fd_sc_hd__nor2_1 _08064_ (.A(_01214_),
    .B(_01216_),
    .Y(_01217_));
 sky130_fd_sc_hd__xor2_1 _08065_ (.A(_01214_),
    .B(_01216_),
    .X(_01218_));
 sky130_fd_sc_hd__nand2_1 _08066_ (.A(_01212_),
    .B(_01218_),
    .Y(_01219_));
 sky130_fd_sc_hd__o22a_1 _08067_ (.A1(net129),
    .A2(net172),
    .B1(net170),
    .B2(net99),
    .X(_01220_));
 sky130_fd_sc_hd__xnor2_1 _08068_ (.A(net207),
    .B(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__o22a_1 _08069_ (.A1(net122),
    .A2(net168),
    .B1(net166),
    .B2(net81),
    .X(_01222_));
 sky130_fd_sc_hd__xnor2_1 _08070_ (.A(net209),
    .B(_01222_),
    .Y(_01223_));
 sky130_fd_sc_hd__o22a_1 _08071_ (.A1(net301),
    .A2(net70),
    .B1(net252),
    .B2(net118),
    .X(_01224_));
 sky130_fd_sc_hd__xnor2_1 _08072_ (.A(net254),
    .B(_01224_),
    .Y(_01225_));
 sky130_fd_sc_hd__or2_1 _08073_ (.A(_01223_),
    .B(_01225_),
    .X(_01226_));
 sky130_fd_sc_hd__xor2_1 _08074_ (.A(_01223_),
    .B(_01225_),
    .X(_01227_));
 sky130_fd_sc_hd__nand2b_1 _08075_ (.A_N(_01221_),
    .B(_01227_),
    .Y(_01228_));
 sky130_fd_sc_hd__xor2_1 _08076_ (.A(_01221_),
    .B(_01227_),
    .X(_01229_));
 sky130_fd_sc_hd__or2_1 _08077_ (.A(_01212_),
    .B(_01218_),
    .X(_01230_));
 sky130_fd_sc_hd__nand2_1 _08078_ (.A(_01219_),
    .B(_01230_),
    .Y(_01231_));
 sky130_fd_sc_hd__nor2_1 _08079_ (.A(_01229_),
    .B(_01231_),
    .Y(_01232_));
 sky130_fd_sc_hd__o21ai_1 _08080_ (.A1(_01229_),
    .A2(_01231_),
    .B1(_01219_),
    .Y(_01233_));
 sky130_fd_sc_hd__o22a_1 _08081_ (.A1(net301),
    .A2(net118),
    .B1(net252),
    .B2(net99),
    .X(_01234_));
 sky130_fd_sc_hd__xnor2_1 _08082_ (.A(net254),
    .B(_01234_),
    .Y(_01235_));
 sky130_fd_sc_hd__o22a_1 _08083_ (.A1(net125),
    .A2(net168),
    .B1(net166),
    .B2(net122),
    .X(_01236_));
 sky130_fd_sc_hd__xnor2_1 _08084_ (.A(net209),
    .B(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__o22a_1 _08085_ (.A1(net81),
    .A2(net172),
    .B1(net170),
    .B2(net129),
    .X(_01238_));
 sky130_fd_sc_hd__xnor2_1 _08086_ (.A(net207),
    .B(_01238_),
    .Y(_01239_));
 sky130_fd_sc_hd__xor2_1 _08087_ (.A(_01235_),
    .B(_01237_),
    .X(_01240_));
 sky130_fd_sc_hd__and2b_1 _08088_ (.A_N(_01239_),
    .B(_01240_),
    .X(_01241_));
 sky130_fd_sc_hd__o21bai_1 _08089_ (.A1(_01235_),
    .A2(_01237_),
    .B1_N(_01241_),
    .Y(_01242_));
 sky130_fd_sc_hd__o22a_1 _08090_ (.A1(net164),
    .A2(net95),
    .B1(net160),
    .B2(net43),
    .X(_01243_));
 sky130_fd_sc_hd__xnor2_1 _08091_ (.A(net139),
    .B(_01243_),
    .Y(_01244_));
 sky130_fd_sc_hd__nand2_1 _08092_ (.A(_01242_),
    .B(_01244_),
    .Y(_01245_));
 sky130_fd_sc_hd__xnor2_1 _08093_ (.A(_01242_),
    .B(_01244_),
    .Y(_01246_));
 sky130_fd_sc_hd__o22a_1 _08094_ (.A1(net223),
    .A2(net37),
    .B1(net35),
    .B2(net162),
    .X(_01247_));
 sky130_fd_sc_hd__xnor2_1 _08095_ (.A(net136),
    .B(_01247_),
    .Y(_01248_));
 sky130_fd_sc_hd__inv_2 _08096_ (.A(_01248_),
    .Y(_01249_));
 sky130_fd_sc_hd__o21ai_1 _08097_ (.A1(_01246_),
    .A2(_01249_),
    .B1(_01245_),
    .Y(_01250_));
 sky130_fd_sc_hd__xnor2_1 _08098_ (.A(_01207_),
    .B(_01233_),
    .Y(_01251_));
 sky130_fd_sc_hd__nand2b_1 _08099_ (.A_N(_01251_),
    .B(_01250_),
    .Y(_01252_));
 sky130_fd_sc_hd__a21bo_2 _08100_ (.A1(_01207_),
    .A2(_01233_),
    .B1_N(_01252_),
    .X(_01253_));
 sky130_fd_sc_hd__xnor2_1 _08101_ (.A(net104),
    .B(_01217_),
    .Y(_01254_));
 sky130_fd_sc_hd__a21oi_1 _08102_ (.A1(_01226_),
    .A2(_01228_),
    .B1(_01254_),
    .Y(_01255_));
 sky130_fd_sc_hd__a21o_1 _08103_ (.A1(net104),
    .A2(_01217_),
    .B1(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__o22a_1 _08104_ (.A1(net79),
    .A2(net142),
    .B1(net140),
    .B2(net124),
    .X(_01257_));
 sky130_fd_sc_hd__xnor2_2 _08105_ (.A(net156),
    .B(_01257_),
    .Y(_01258_));
 sky130_fd_sc_hd__inv_2 _08106_ (.A(_01258_),
    .Y(_01259_));
 sky130_fd_sc_hd__o22a_2 _08107_ (.A1(net83),
    .A2(net146),
    .B1(net145),
    .B2(net131),
    .X(_01260_));
 sky130_fd_sc_hd__xnor2_4 _08108_ (.A(net159),
    .B(_01260_),
    .Y(_01261_));
 sky130_fd_sc_hd__nor2_2 _08109_ (.A(_01259_),
    .B(_01261_),
    .Y(_01262_));
 sky130_fd_sc_hd__xnor2_2 _08110_ (.A(_01258_),
    .B(_01261_),
    .Y(_01263_));
 sky130_fd_sc_hd__o22a_1 _08111_ (.A1(net118),
    .A2(net170),
    .B1(net99),
    .B2(net172),
    .X(_01264_));
 sky130_fd_sc_hd__xnor2_2 _08112_ (.A(net207),
    .B(_01264_),
    .Y(_01265_));
 sky130_fd_sc_hd__inv_2 _08113_ (.A(_01265_),
    .Y(_01266_));
 sky130_fd_sc_hd__o22a_2 _08114_ (.A1(net81),
    .A2(net168),
    .B1(net166),
    .B2(net129),
    .X(_01267_));
 sky130_fd_sc_hd__xnor2_4 _08115_ (.A(net209),
    .B(_01267_),
    .Y(_01268_));
 sky130_fd_sc_hd__o22a_2 _08116_ (.A1(net301),
    .A2(net76),
    .B1(net70),
    .B2(net252),
    .X(_01269_));
 sky130_fd_sc_hd__xnor2_4 _08117_ (.A(net254),
    .B(_01269_),
    .Y(_01270_));
 sky130_fd_sc_hd__nor2_1 _08118_ (.A(_01268_),
    .B(_01270_),
    .Y(_01271_));
 sky130_fd_sc_hd__xor2_4 _08119_ (.A(_01268_),
    .B(_01270_),
    .X(_01272_));
 sky130_fd_sc_hd__xnor2_2 _08120_ (.A(_01265_),
    .B(_01272_),
    .Y(_01273_));
 sky130_fd_sc_hd__and2_1 _08121_ (.A(_01263_),
    .B(_01273_),
    .X(_01274_));
 sky130_fd_sc_hd__o22a_1 _08122_ (.A1(net151),
    .A2(net93),
    .B1(net87),
    .B2(net153),
    .X(_01275_));
 sky130_fd_sc_hd__xnor2_2 _08123_ (.A(net192),
    .B(_01275_),
    .Y(_01276_));
 sky130_fd_sc_hd__o22a_1 _08124_ (.A1(net117),
    .A2(net132),
    .B1(net89),
    .B2(net115),
    .X(_01277_));
 sky130_fd_sc_hd__xnor2_2 _08125_ (.A(net181),
    .B(_01277_),
    .Y(_01278_));
 sky130_fd_sc_hd__o22a_1 _08126_ (.A1(net125),
    .A2(net176),
    .B1(net174),
    .B2(net122),
    .X(_01279_));
 sky130_fd_sc_hd__xnor2_2 _08127_ (.A(net188),
    .B(_01279_),
    .Y(_01280_));
 sky130_fd_sc_hd__xor2_2 _08128_ (.A(_01278_),
    .B(_01280_),
    .X(_01281_));
 sky130_fd_sc_hd__and2b_1 _08129_ (.A_N(_01276_),
    .B(_01281_),
    .X(_01282_));
 sky130_fd_sc_hd__xnor2_2 _08130_ (.A(_01276_),
    .B(_01281_),
    .Y(_01283_));
 sky130_fd_sc_hd__xor2_2 _08131_ (.A(_01263_),
    .B(_01273_),
    .X(_01284_));
 sky130_fd_sc_hd__a21oi_2 _08132_ (.A1(_01283_),
    .A2(_01284_),
    .B1(_01274_),
    .Y(_01285_));
 sky130_fd_sc_hd__o22a_1 _08133_ (.A1(net164),
    .A2(net43),
    .B1(net95),
    .B2(net148),
    .X(_01286_));
 sky130_fd_sc_hd__xnor2_1 _08134_ (.A(net139),
    .B(_01286_),
    .Y(_01287_));
 sky130_fd_sc_hd__or2_1 _08135_ (.A(net226),
    .B(net39),
    .X(_01288_));
 sky130_fd_sc_hd__xnor2_1 _08136_ (.A(net104),
    .B(_01288_),
    .Y(_01289_));
 sky130_fd_sc_hd__xnor2_1 _08137_ (.A(_01287_),
    .B(_01289_),
    .Y(_01290_));
 sky130_fd_sc_hd__o22a_1 _08138_ (.A1(net162),
    .A2(net37),
    .B1(net35),
    .B2(net160),
    .X(_01291_));
 sky130_fd_sc_hd__xnor2_1 _08139_ (.A(_00436_),
    .B(_01291_),
    .Y(_01292_));
 sky130_fd_sc_hd__nor2_1 _08140_ (.A(_01290_),
    .B(_01292_),
    .Y(_01293_));
 sky130_fd_sc_hd__a21oi_2 _08141_ (.A1(_01287_),
    .A2(_01289_),
    .B1(_01293_),
    .Y(_01294_));
 sky130_fd_sc_hd__nor2_1 _08142_ (.A(_01285_),
    .B(_01294_),
    .Y(_01295_));
 sky130_fd_sc_hd__xor2_2 _08143_ (.A(_01285_),
    .B(_01294_),
    .X(_01296_));
 sky130_fd_sc_hd__xnor2_2 _08144_ (.A(_01256_),
    .B(_01296_),
    .Y(_01297_));
 sky130_fd_sc_hd__and2b_1 _08145_ (.A_N(_01297_),
    .B(_01253_),
    .X(_01298_));
 sky130_fd_sc_hd__xnor2_2 _08146_ (.A(_01283_),
    .B(_01284_),
    .Y(_01299_));
 sky130_fd_sc_hd__and2_1 _08147_ (.A(_01290_),
    .B(_01292_),
    .X(_01300_));
 sky130_fd_sc_hd__or2_2 _08148_ (.A(_01293_),
    .B(_01300_),
    .X(_01301_));
 sky130_fd_sc_hd__and3_1 _08149_ (.A(_01226_),
    .B(_01228_),
    .C(_01254_),
    .X(_01302_));
 sky130_fd_sc_hd__or2_1 _08150_ (.A(_01255_),
    .B(_01302_),
    .X(_01303_));
 sky130_fd_sc_hd__xor2_1 _08151_ (.A(_01299_),
    .B(_01301_),
    .X(_01304_));
 sky130_fd_sc_hd__and2b_1 _08152_ (.A_N(_01303_),
    .B(_01304_),
    .X(_01305_));
 sky130_fd_sc_hd__o21bai_4 _08153_ (.A1(_01299_),
    .A2(_01301_),
    .B1_N(_01305_),
    .Y(_01306_));
 sky130_fd_sc_hd__xnor2_4 _08154_ (.A(_01253_),
    .B(_01297_),
    .Y(_01307_));
 sky130_fd_sc_hd__a21o_2 _08155_ (.A1(_01306_),
    .A2(_01307_),
    .B1(_01298_),
    .X(_01308_));
 sky130_fd_sc_hd__or2_1 _08156_ (.A(_01171_),
    .B(_01172_),
    .X(_01309_));
 sky130_fd_sc_hd__nand2_2 _08157_ (.A(_01173_),
    .B(_01309_),
    .Y(_01310_));
 sky130_fd_sc_hd__a21o_1 _08158_ (.A1(_01137_),
    .A2(_01139_),
    .B1(_01138_),
    .X(_01311_));
 sky130_fd_sc_hd__xnor2_1 _08159_ (.A(_01141_),
    .B(_01151_),
    .Y(_01312_));
 sky130_fd_sc_hd__and3_1 _08160_ (.A(_01140_),
    .B(_01311_),
    .C(_01312_),
    .X(_01313_));
 sky130_fd_sc_hd__a21oi_1 _08161_ (.A1(_01140_),
    .A2(_01311_),
    .B1(_01312_),
    .Y(_01314_));
 sky130_fd_sc_hd__nor2_2 _08162_ (.A(_01313_),
    .B(_01314_),
    .Y(_01315_));
 sky130_fd_sc_hd__xnor2_4 _08163_ (.A(_01310_),
    .B(_01315_),
    .Y(_01316_));
 sky130_fd_sc_hd__xnor2_4 _08164_ (.A(_01162_),
    .B(_01163_),
    .Y(_01317_));
 sky130_fd_sc_hd__xnor2_4 _08165_ (.A(_01149_),
    .B(_01150_),
    .Y(_01318_));
 sky130_fd_sc_hd__and2_1 _08166_ (.A(_01168_),
    .B(_01170_),
    .X(_01319_));
 sky130_fd_sc_hd__or2_2 _08167_ (.A(_01171_),
    .B(_01319_),
    .X(_01320_));
 sky130_fd_sc_hd__or2_1 _08168_ (.A(_01318_),
    .B(_01320_),
    .X(_01321_));
 sky130_fd_sc_hd__xnor2_4 _08169_ (.A(_01318_),
    .B(_01320_),
    .Y(_01322_));
 sky130_fd_sc_hd__xnor2_4 _08170_ (.A(_01317_),
    .B(_01322_),
    .Y(_01323_));
 sky130_fd_sc_hd__o22a_1 _08171_ (.A1(net148),
    .A2(net43),
    .B1(net95),
    .B2(net142),
    .X(_01324_));
 sky130_fd_sc_hd__xnor2_1 _08172_ (.A(net139),
    .B(_01324_),
    .Y(_01325_));
 sky130_fd_sc_hd__o22a_1 _08173_ (.A1(net223),
    .A2(net41),
    .B1(net39),
    .B2(net162),
    .X(_01326_));
 sky130_fd_sc_hd__xnor2_1 _08174_ (.A(net104),
    .B(_01326_),
    .Y(_01327_));
 sky130_fd_sc_hd__and2_1 _08175_ (.A(_01325_),
    .B(_01327_),
    .X(_01328_));
 sky130_fd_sc_hd__nor2_1 _08176_ (.A(_01325_),
    .B(_01327_),
    .Y(_01329_));
 sky130_fd_sc_hd__nor2_1 _08177_ (.A(_01328_),
    .B(_01329_),
    .Y(_01330_));
 sky130_fd_sc_hd__o22a_1 _08178_ (.A1(net160),
    .A2(net37),
    .B1(net35),
    .B2(net164),
    .X(_01331_));
 sky130_fd_sc_hd__xnor2_1 _08179_ (.A(net136),
    .B(_01331_),
    .Y(_01332_));
 sky130_fd_sc_hd__and2_1 _08180_ (.A(_01330_),
    .B(_01332_),
    .X(_01333_));
 sky130_fd_sc_hd__nor2_1 _08181_ (.A(_01330_),
    .B(_01332_),
    .Y(_01334_));
 sky130_fd_sc_hd__nor2_2 _08182_ (.A(_01333_),
    .B(_01334_),
    .Y(_01335_));
 sky130_fd_sc_hd__and2b_1 _08183_ (.A_N(_01323_),
    .B(_01335_),
    .X(_01336_));
 sky130_fd_sc_hd__o21ba_2 _08184_ (.A1(_01278_),
    .A2(_01280_),
    .B1_N(_01282_),
    .X(_01337_));
 sky130_fd_sc_hd__a21oi_4 _08185_ (.A1(_01266_),
    .A2(_01272_),
    .B1(_01271_),
    .Y(_01338_));
 sky130_fd_sc_hd__xnor2_4 _08186_ (.A(_01262_),
    .B(_01338_),
    .Y(_01339_));
 sky130_fd_sc_hd__nand2b_1 _08187_ (.A_N(_01337_),
    .B(_01339_),
    .Y(_01340_));
 sky130_fd_sc_hd__xnor2_4 _08188_ (.A(_01337_),
    .B(_01339_),
    .Y(_01341_));
 sky130_fd_sc_hd__xnor2_4 _08189_ (.A(_01323_),
    .B(_01335_),
    .Y(_01342_));
 sky130_fd_sc_hd__a21o_2 _08190_ (.A1(_01341_),
    .A2(_01342_),
    .B1(_01336_),
    .X(_01343_));
 sky130_fd_sc_hd__o31ai_4 _08191_ (.A1(_01259_),
    .A2(_01261_),
    .A3(_01338_),
    .B1(_01340_),
    .Y(_01344_));
 sky130_fd_sc_hd__o21ai_2 _08192_ (.A1(_01317_),
    .A2(_01322_),
    .B1(_01321_),
    .Y(_01345_));
 sky130_fd_sc_hd__nor2_1 _08193_ (.A(_01328_),
    .B(_01333_),
    .Y(_01346_));
 sky130_fd_sc_hd__o21ai_1 _08194_ (.A1(_01328_),
    .A2(_01333_),
    .B1(_01345_),
    .Y(_01347_));
 sky130_fd_sc_hd__xnor2_2 _08195_ (.A(_01345_),
    .B(_01346_),
    .Y(_01348_));
 sky130_fd_sc_hd__xnor2_2 _08196_ (.A(_01344_),
    .B(_01348_),
    .Y(_01349_));
 sky130_fd_sc_hd__a21oi_2 _08197_ (.A1(_01256_),
    .A2(_01296_),
    .B1(_01295_),
    .Y(_01350_));
 sky130_fd_sc_hd__xnor2_2 _08198_ (.A(_01349_),
    .B(_01350_),
    .Y(_01351_));
 sky130_fd_sc_hd__nand2b_1 _08199_ (.A_N(_01351_),
    .B(_01343_),
    .Y(_01352_));
 sky130_fd_sc_hd__xnor2_4 _08200_ (.A(_01343_),
    .B(_01351_),
    .Y(_01353_));
 sky130_fd_sc_hd__and2_1 _08201_ (.A(_01316_),
    .B(_01353_),
    .X(_01354_));
 sky130_fd_sc_hd__xor2_4 _08202_ (.A(_01316_),
    .B(_01353_),
    .X(_01355_));
 sky130_fd_sc_hd__xnor2_4 _08203_ (.A(_01308_),
    .B(_01355_),
    .Y(_01356_));
 sky130_fd_sc_hd__xnor2_4 _08204_ (.A(_01306_),
    .B(_01307_),
    .Y(_01357_));
 sky130_fd_sc_hd__xnor2_4 _08205_ (.A(_01341_),
    .B(_01342_),
    .Y(_01358_));
 sky130_fd_sc_hd__nor2_1 _08206_ (.A(_01357_),
    .B(_01358_),
    .Y(_01359_));
 sky130_fd_sc_hd__xnor2_1 _08207_ (.A(_01250_),
    .B(_01251_),
    .Y(_01360_));
 sky130_fd_sc_hd__o22a_1 _08208_ (.A1(net117),
    .A2(net146),
    .B1(net145),
    .B2(net115),
    .X(_01361_));
 sky130_fd_sc_hd__xnor2_1 _08209_ (.A(net181),
    .B(_01361_),
    .Y(_01362_));
 sky130_fd_sc_hd__o22a_1 _08210_ (.A1(net79),
    .A2(net164),
    .B1(net148),
    .B2(net124),
    .X(_01363_));
 sky130_fd_sc_hd__xor2_1 _08211_ (.A(net156),
    .B(_01363_),
    .X(_01364_));
 sky130_fd_sc_hd__nor2_1 _08212_ (.A(_01362_),
    .B(_01364_),
    .Y(_01365_));
 sky130_fd_sc_hd__xnor2_1 _08213_ (.A(_01362_),
    .B(_01364_),
    .Y(_01366_));
 sky130_fd_sc_hd__o22a_1 _08214_ (.A1(net83),
    .A2(net142),
    .B1(net140),
    .B2(net131),
    .X(_01367_));
 sky130_fd_sc_hd__xnor2_1 _08215_ (.A(net159),
    .B(_01367_),
    .Y(_01368_));
 sky130_fd_sc_hd__o21ba_1 _08216_ (.A1(_01366_),
    .A2(_01368_),
    .B1_N(_01365_),
    .X(_01369_));
 sky130_fd_sc_hd__o22a_1 _08217_ (.A1(net129),
    .A2(net252),
    .B1(net101),
    .B2(net302),
    .X(_01370_));
 sky130_fd_sc_hd__xnor2_1 _08218_ (.A(_00187_),
    .B(_01370_),
    .Y(_01371_));
 sky130_fd_sc_hd__or2_1 _08219_ (.A(net122),
    .B(net172),
    .X(_01372_));
 sky130_fd_sc_hd__a21o_1 _08220_ (.A1(_06456_),
    .A2(_06457_),
    .B1(net170),
    .X(_01373_));
 sky130_fd_sc_hd__a21o_1 _08221_ (.A1(_01372_),
    .A2(_01373_),
    .B1(net207),
    .X(_01374_));
 sky130_fd_sc_hd__nand3_1 _08222_ (.A(net207),
    .B(_01372_),
    .C(_01373_),
    .Y(_01375_));
 sky130_fd_sc_hd__nand3_2 _08223_ (.A(_01371_),
    .B(_01374_),
    .C(_01375_),
    .Y(_01376_));
 sky130_fd_sc_hd__xor2_1 _08224_ (.A(_01209_),
    .B(_01211_),
    .X(_01377_));
 sky130_fd_sc_hd__and2b_1 _08225_ (.A_N(_01376_),
    .B(_01377_),
    .X(_01378_));
 sky130_fd_sc_hd__xnor2_1 _08226_ (.A(_01239_),
    .B(_01240_),
    .Y(_01379_));
 sky130_fd_sc_hd__xnor2_1 _08227_ (.A(_01376_),
    .B(_01377_),
    .Y(_01380_));
 sky130_fd_sc_hd__a21oi_1 _08228_ (.A1(_01379_),
    .A2(_01380_),
    .B1(_01378_),
    .Y(_01381_));
 sky130_fd_sc_hd__xor2_1 _08229_ (.A(_01369_),
    .B(_01381_),
    .X(_01382_));
 sky130_fd_sc_hd__nor2_1 _08230_ (.A(net223),
    .B(net35),
    .Y(_01383_));
 sky130_fd_sc_hd__o22a_1 _08231_ (.A1(net163),
    .A2(net43),
    .B1(net95),
    .B2(net161),
    .X(_01384_));
 sky130_fd_sc_hd__xnor2_1 _08232_ (.A(net139),
    .B(_01384_),
    .Y(_01385_));
 sky130_fd_sc_hd__or3_1 _08233_ (.A(net223),
    .B(net35),
    .C(_01385_),
    .X(_01386_));
 sky130_fd_sc_hd__o21a_1 _08234_ (.A1(net136),
    .A2(_01383_),
    .B1(_01386_),
    .X(_01387_));
 sky130_fd_sc_hd__o21ai_1 _08235_ (.A1(net136),
    .A2(_01383_),
    .B1(_01386_),
    .Y(_01388_));
 sky130_fd_sc_hd__o2bb2a_1 _08236_ (.A1_N(_01382_),
    .A2_N(_01387_),
    .B1(_01369_),
    .B2(_01381_),
    .X(_01389_));
 sky130_fd_sc_hd__nand2b_1 _08237_ (.A_N(_01389_),
    .B(_01360_),
    .Y(_01390_));
 sky130_fd_sc_hd__and2_1 _08238_ (.A(_01203_),
    .B(_01205_),
    .X(_01391_));
 sky130_fd_sc_hd__or2_1 _08239_ (.A(_01206_),
    .B(_01391_),
    .X(_01392_));
 sky130_fd_sc_hd__and2_1 _08240_ (.A(_01229_),
    .B(_01231_),
    .X(_01393_));
 sky130_fd_sc_hd__or3_1 _08241_ (.A(_01232_),
    .B(_01392_),
    .C(_01393_),
    .X(_01394_));
 sky130_fd_sc_hd__xnor2_1 _08242_ (.A(_01246_),
    .B(_01248_),
    .Y(_01395_));
 sky130_fd_sc_hd__o21ai_1 _08243_ (.A1(_01232_),
    .A2(_01393_),
    .B1(_01392_),
    .Y(_01396_));
 sky130_fd_sc_hd__and3_1 _08244_ (.A(_01394_),
    .B(_01395_),
    .C(_01396_),
    .X(_01397_));
 sky130_fd_sc_hd__a21bo_1 _08245_ (.A1(_01395_),
    .A2(_01396_),
    .B1_N(_01394_),
    .X(_01398_));
 sky130_fd_sc_hd__xor2_1 _08246_ (.A(_01360_),
    .B(_01389_),
    .X(_01399_));
 sky130_fd_sc_hd__nand2b_1 _08247_ (.A_N(_01399_),
    .B(_01398_),
    .Y(_01400_));
 sky130_fd_sc_hd__nand2_2 _08248_ (.A(_01390_),
    .B(_01400_),
    .Y(_01401_));
 sky130_fd_sc_hd__xor2_4 _08249_ (.A(_01357_),
    .B(_01358_),
    .X(_01402_));
 sky130_fd_sc_hd__a21oi_4 _08250_ (.A1(_01401_),
    .A2(_01402_),
    .B1(_01359_),
    .Y(_01403_));
 sky130_fd_sc_hd__nor2_1 _08251_ (.A(_01356_),
    .B(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__xor2_4 _08252_ (.A(_01356_),
    .B(_01403_),
    .X(_01405_));
 sky130_fd_sc_hd__a21oi_2 _08253_ (.A1(_01308_),
    .A2(_01355_),
    .B1(_01354_),
    .Y(_01406_));
 sky130_fd_sc_hd__o21ai_2 _08254_ (.A1(_01349_),
    .A2(_01350_),
    .B1(_01352_),
    .Y(_01407_));
 sky130_fd_sc_hd__o21ba_1 _08255_ (.A1(_01310_),
    .A2(_01314_),
    .B1_N(_01313_),
    .X(_01408_));
 sky130_fd_sc_hd__a21bo_1 _08256_ (.A1(_01344_),
    .A2(_01348_),
    .B1_N(_01347_),
    .X(_01409_));
 sky130_fd_sc_hd__xnor2_1 _08257_ (.A(_01174_),
    .B(_01176_),
    .Y(_01410_));
 sky130_fd_sc_hd__nand2b_1 _08258_ (.A_N(_01410_),
    .B(_01409_),
    .Y(_01411_));
 sky130_fd_sc_hd__xnor2_2 _08259_ (.A(_01409_),
    .B(_01410_),
    .Y(_01412_));
 sky130_fd_sc_hd__nand2b_1 _08260_ (.A_N(_01408_),
    .B(_01412_),
    .Y(_01413_));
 sky130_fd_sc_hd__xnor2_2 _08261_ (.A(_01408_),
    .B(_01412_),
    .Y(_01414_));
 sky130_fd_sc_hd__xor2_2 _08262_ (.A(_01183_),
    .B(_01185_),
    .X(_01415_));
 sky130_fd_sc_hd__nand2_1 _08263_ (.A(_01414_),
    .B(_01415_),
    .Y(_01416_));
 sky130_fd_sc_hd__xnor2_2 _08264_ (.A(_01414_),
    .B(_01415_),
    .Y(_01417_));
 sky130_fd_sc_hd__nand2b_1 _08265_ (.A_N(_01417_),
    .B(_01407_),
    .Y(_01418_));
 sky130_fd_sc_hd__xor2_2 _08266_ (.A(_01407_),
    .B(_01417_),
    .X(_01419_));
 sky130_fd_sc_hd__xor2_2 _08267_ (.A(_01406_),
    .B(_01419_),
    .X(_01420_));
 sky130_fd_sc_hd__xnor2_1 _08268_ (.A(_01382_),
    .B(_01388_),
    .Y(_01421_));
 sky130_fd_sc_hd__a21o_1 _08269_ (.A1(_01374_),
    .A2(_01375_),
    .B1(_01371_),
    .X(_01422_));
 sky130_fd_sc_hd__o22a_1 _08270_ (.A1(net225),
    .A2(net43),
    .B1(net95),
    .B2(net163),
    .X(_01423_));
 sky130_fd_sc_hd__xnor2_1 _08271_ (.A(net139),
    .B(_01423_),
    .Y(_01424_));
 sky130_fd_sc_hd__and3_1 _08272_ (.A(_01376_),
    .B(_01422_),
    .C(_01424_),
    .X(_01425_));
 sky130_fd_sc_hd__a21oi_1 _08273_ (.A1(_06456_),
    .A2(_06457_),
    .B1(net253),
    .Y(_01426_));
 sky130_fd_sc_hd__nor2_1 _08274_ (.A(net301),
    .B(net129),
    .Y(_01427_));
 sky130_fd_sc_hd__o21a_1 _08275_ (.A1(_01426_),
    .A2(_01427_),
    .B1(_00187_),
    .X(_01428_));
 sky130_fd_sc_hd__nor3_1 _08276_ (.A(_00187_),
    .B(_01426_),
    .C(_01427_),
    .Y(_01429_));
 sky130_fd_sc_hd__o22a_1 _08277_ (.A1(net127),
    .A2(net172),
    .B1(net171),
    .B2(net122),
    .X(_01430_));
 sky130_fd_sc_hd__xnor2_1 _08278_ (.A(net207),
    .B(_01430_),
    .Y(_01431_));
 sky130_fd_sc_hd__nor3_1 _08279_ (.A(_01428_),
    .B(_01429_),
    .C(_01431_),
    .Y(_01432_));
 sky130_fd_sc_hd__or3_1 _08280_ (.A(_01428_),
    .B(_01429_),
    .C(_01431_),
    .X(_01433_));
 sky130_fd_sc_hd__a21oi_1 _08281_ (.A1(_01376_),
    .A2(_01422_),
    .B1(_01424_),
    .Y(_01434_));
 sky130_fd_sc_hd__a21o_1 _08282_ (.A1(_01376_),
    .A2(_01422_),
    .B1(_01424_),
    .X(_01435_));
 sky130_fd_sc_hd__and3b_1 _08283_ (.A_N(_01425_),
    .B(_01432_),
    .C(_01435_),
    .X(_01436_));
 sky130_fd_sc_hd__a21o_1 _08284_ (.A1(_01432_),
    .A2(_01435_),
    .B1(_01425_),
    .X(_01437_));
 sky130_fd_sc_hd__o22a_1 _08285_ (.A1(net127),
    .A2(net167),
    .B1(net93),
    .B2(net169),
    .X(_01438_));
 sky130_fd_sc_hd__xnor2_1 _08286_ (.A(net211),
    .B(_01438_),
    .Y(_01439_));
 sky130_fd_sc_hd__o22a_1 _08287_ (.A1(net153),
    .A2(net145),
    .B1(net134),
    .B2(net151),
    .X(_01440_));
 sky130_fd_sc_hd__xnor2_1 _08288_ (.A(net192),
    .B(_01440_),
    .Y(_01441_));
 sky130_fd_sc_hd__o22a_1 _08289_ (.A1(net176),
    .A2(net91),
    .B1(net88),
    .B2(net175),
    .X(_01442_));
 sky130_fd_sc_hd__xnor2_1 _08290_ (.A(net190),
    .B(_01442_),
    .Y(_01443_));
 sky130_fd_sc_hd__xor2_1 _08291_ (.A(_01439_),
    .B(_01441_),
    .X(_01444_));
 sky130_fd_sc_hd__nand2b_1 _08292_ (.A_N(_01443_),
    .B(_01444_),
    .Y(_01445_));
 sky130_fd_sc_hd__o21a_1 _08293_ (.A1(_01439_),
    .A2(_01441_),
    .B1(_01445_),
    .X(_01446_));
 sky130_fd_sc_hd__o21ba_1 _08294_ (.A1(_01425_),
    .A2(_01436_),
    .B1_N(_01446_),
    .X(_01447_));
 sky130_fd_sc_hd__o22a_1 _08295_ (.A1(net115),
    .A2(net146),
    .B1(net140),
    .B2(net117),
    .X(_01448_));
 sky130_fd_sc_hd__xnor2_1 _08296_ (.A(net181),
    .B(_01448_),
    .Y(_01449_));
 sky130_fd_sc_hd__o22a_1 _08297_ (.A1(net124),
    .A2(net164),
    .B1(net161),
    .B2(net79),
    .X(_01450_));
 sky130_fd_sc_hd__xor2_1 _08298_ (.A(net156),
    .B(_01450_),
    .X(_01451_));
 sky130_fd_sc_hd__xnor2_1 _08299_ (.A(_01449_),
    .B(_01451_),
    .Y(_01452_));
 sky130_fd_sc_hd__o22a_1 _08300_ (.A1(net83),
    .A2(net148),
    .B1(net142),
    .B2(net131),
    .X(_01453_));
 sky130_fd_sc_hd__xnor2_1 _08301_ (.A(net159),
    .B(_01453_),
    .Y(_01454_));
 sky130_fd_sc_hd__or2_1 _08302_ (.A(_01452_),
    .B(_01454_),
    .X(_01455_));
 sky130_fd_sc_hd__o21ai_1 _08303_ (.A1(_01449_),
    .A2(_01451_),
    .B1(_01455_),
    .Y(_01456_));
 sky130_fd_sc_hd__xnor2_1 _08304_ (.A(_01437_),
    .B(_01446_),
    .Y(_01457_));
 sky130_fd_sc_hd__a21o_1 _08305_ (.A1(_01456_),
    .A2(_01457_),
    .B1(_01447_),
    .X(_01458_));
 sky130_fd_sc_hd__xnor2_1 _08306_ (.A(_01366_),
    .B(_01368_),
    .Y(_01459_));
 sky130_fd_sc_hd__xnor2_1 _08307_ (.A(_01379_),
    .B(_01380_),
    .Y(_01460_));
 sky130_fd_sc_hd__xor2_1 _08308_ (.A(_01459_),
    .B(_01460_),
    .X(_01461_));
 sky130_fd_sc_hd__xnor2_1 _08309_ (.A(_01383_),
    .B(_01385_),
    .Y(_01462_));
 sky130_fd_sc_hd__and2b_1 _08310_ (.A_N(_01462_),
    .B(_01461_),
    .X(_01463_));
 sky130_fd_sc_hd__o21ba_1 _08311_ (.A1(_01459_),
    .A2(_01460_),
    .B1_N(_01463_),
    .X(_01464_));
 sky130_fd_sc_hd__xor2_1 _08312_ (.A(_01421_),
    .B(_01458_),
    .X(_01465_));
 sky130_fd_sc_hd__nand2b_1 _08313_ (.A_N(_01464_),
    .B(_01465_),
    .Y(_01466_));
 sky130_fd_sc_hd__a21bo_1 _08314_ (.A1(_01421_),
    .A2(_01458_),
    .B1_N(_01466_),
    .X(_01467_));
 sky130_fd_sc_hd__xnor2_1 _08315_ (.A(_01398_),
    .B(_01399_),
    .Y(_01468_));
 sky130_fd_sc_hd__xnor2_1 _08316_ (.A(_01303_),
    .B(_01304_),
    .Y(_01469_));
 sky130_fd_sc_hd__and2_1 _08317_ (.A(_01468_),
    .B(_01469_),
    .X(_01470_));
 sky130_fd_sc_hd__xor2_1 _08318_ (.A(_01468_),
    .B(_01469_),
    .X(_01471_));
 sky130_fd_sc_hd__xnor2_1 _08319_ (.A(_01467_),
    .B(_01471_),
    .Y(_01472_));
 sky130_fd_sc_hd__xnor2_1 _08320_ (.A(_01464_),
    .B(_01465_),
    .Y(_01473_));
 sky130_fd_sc_hd__a21oi_1 _08321_ (.A1(_01394_),
    .A2(_01396_),
    .B1(_01395_),
    .Y(_01474_));
 sky130_fd_sc_hd__nor2_1 _08322_ (.A(_01397_),
    .B(_01474_),
    .Y(_01475_));
 sky130_fd_sc_hd__xnor2_1 _08323_ (.A(_01456_),
    .B(_01457_),
    .Y(_01476_));
 sky130_fd_sc_hd__o22a_1 _08324_ (.A1(net153),
    .A2(net146),
    .B1(net145),
    .B2(net151),
    .X(_01477_));
 sky130_fd_sc_hd__xnor2_1 _08325_ (.A(net192),
    .B(_01477_),
    .Y(_01478_));
 sky130_fd_sc_hd__o22a_1 _08326_ (.A1(net166),
    .A2(net93),
    .B1(net88),
    .B2(net169),
    .X(_01479_));
 sky130_fd_sc_hd__xnor2_1 _08327_ (.A(net211),
    .B(_01479_),
    .Y(_01480_));
 sky130_fd_sc_hd__nor2_1 _08328_ (.A(_01478_),
    .B(_01480_),
    .Y(_01481_));
 sky130_fd_sc_hd__o22a_1 _08329_ (.A1(net176),
    .A2(net132),
    .B1(net89),
    .B2(net174),
    .X(_01482_));
 sky130_fd_sc_hd__xnor2_1 _08330_ (.A(net188),
    .B(_01482_),
    .Y(_01483_));
 sky130_fd_sc_hd__xor2_1 _08331_ (.A(_01478_),
    .B(_01480_),
    .X(_01484_));
 sky130_fd_sc_hd__and2b_1 _08332_ (.A_N(_01483_),
    .B(_01484_),
    .X(_01485_));
 sky130_fd_sc_hd__or2_1 _08333_ (.A(net225),
    .B(net95),
    .X(_01486_));
 sky130_fd_sc_hd__o21ai_1 _08334_ (.A1(_01428_),
    .A2(_01429_),
    .B1(_01431_),
    .Y(_01487_));
 sky130_fd_sc_hd__and2_1 _08335_ (.A(_01433_),
    .B(_01487_),
    .X(_01488_));
 sky130_fd_sc_hd__a21o_1 _08336_ (.A1(_01433_),
    .A2(_01487_),
    .B1(_01486_),
    .X(_01489_));
 sky130_fd_sc_hd__nand2b_1 _08337_ (.A_N(net139),
    .B(_01486_),
    .Y(_01490_));
 sky130_fd_sc_hd__o211ai_2 _08338_ (.A1(_01481_),
    .A2(_01485_),
    .B1(_01489_),
    .C1(_01490_),
    .Y(_01491_));
 sky130_fd_sc_hd__o22a_1 _08339_ (.A1(net117),
    .A2(net142),
    .B1(net140),
    .B2(net115),
    .X(_01492_));
 sky130_fd_sc_hd__xnor2_1 _08340_ (.A(net181),
    .B(_01492_),
    .Y(_01493_));
 sky130_fd_sc_hd__o22a_1 _08341_ (.A1(net79),
    .A2(net163),
    .B1(net161),
    .B2(net124),
    .X(_01494_));
 sky130_fd_sc_hd__xor2_1 _08342_ (.A(net156),
    .B(_01494_),
    .X(_01495_));
 sky130_fd_sc_hd__or2_1 _08343_ (.A(_01493_),
    .B(_01495_),
    .X(_01496_));
 sky130_fd_sc_hd__xnor2_1 _08344_ (.A(_01493_),
    .B(_01495_),
    .Y(_01497_));
 sky130_fd_sc_hd__o22a_1 _08345_ (.A1(net83),
    .A2(net164),
    .B1(net148),
    .B2(net131),
    .X(_01498_));
 sky130_fd_sc_hd__xnor2_1 _08346_ (.A(net159),
    .B(_01498_),
    .Y(_01499_));
 sky130_fd_sc_hd__o21ai_1 _08347_ (.A1(_01497_),
    .A2(_01499_),
    .B1(_01496_),
    .Y(_01500_));
 sky130_fd_sc_hd__a211o_1 _08348_ (.A1(_01489_),
    .A2(_01490_),
    .B1(_01481_),
    .C1(_01485_),
    .X(_01501_));
 sky130_fd_sc_hd__nand3_1 _08349_ (.A(_01491_),
    .B(_01500_),
    .C(_01501_),
    .Y(_01502_));
 sky130_fd_sc_hd__and2_1 _08350_ (.A(_01491_),
    .B(_01502_),
    .X(_01503_));
 sky130_fd_sc_hd__o21a_1 _08351_ (.A1(_01425_),
    .A2(_01434_),
    .B1(_01433_),
    .X(_01504_));
 sky130_fd_sc_hd__xor2_1 _08352_ (.A(_01443_),
    .B(_01444_),
    .X(_01505_));
 sky130_fd_sc_hd__or3_1 _08353_ (.A(_01436_),
    .B(_01504_),
    .C(_01505_),
    .X(_01506_));
 sky130_fd_sc_hd__nand2_1 _08354_ (.A(_01452_),
    .B(_01454_),
    .Y(_01507_));
 sky130_fd_sc_hd__and2_1 _08355_ (.A(_01455_),
    .B(_01507_),
    .X(_01508_));
 sky130_fd_sc_hd__o21ai_1 _08356_ (.A1(_01436_),
    .A2(_01504_),
    .B1(_01505_),
    .Y(_01509_));
 sky130_fd_sc_hd__nand3_1 _08357_ (.A(_01506_),
    .B(_01508_),
    .C(_01509_),
    .Y(_01510_));
 sky130_fd_sc_hd__nand2_1 _08358_ (.A(_01506_),
    .B(_01510_),
    .Y(_01511_));
 sky130_fd_sc_hd__xnor2_1 _08359_ (.A(_01476_),
    .B(_01503_),
    .Y(_01512_));
 sky130_fd_sc_hd__nand2b_1 _08360_ (.A_N(_01512_),
    .B(_01511_),
    .Y(_01513_));
 sky130_fd_sc_hd__o21ai_1 _08361_ (.A1(_01476_),
    .A2(_01503_),
    .B1(_01513_),
    .Y(_01514_));
 sky130_fd_sc_hd__xnor2_1 _08362_ (.A(_01473_),
    .B(_01475_),
    .Y(_01515_));
 sky130_fd_sc_hd__and2b_1 _08363_ (.A_N(_01515_),
    .B(_01514_),
    .X(_01516_));
 sky130_fd_sc_hd__a21oi_1 _08364_ (.A1(_01473_),
    .A2(_01475_),
    .B1(_01516_),
    .Y(_01517_));
 sky130_fd_sc_hd__nor2_1 _08365_ (.A(_01472_),
    .B(_01517_),
    .Y(_01518_));
 sky130_fd_sc_hd__and2_1 _08366_ (.A(_01472_),
    .B(_01517_),
    .X(_01519_));
 sky130_fd_sc_hd__nor2_2 _08367_ (.A(_01518_),
    .B(_01519_),
    .Y(_01520_));
 sky130_fd_sc_hd__a21o_1 _08368_ (.A1(_01467_),
    .A2(_01471_),
    .B1(_01470_),
    .X(_01521_));
 sky130_fd_sc_hd__xor2_2 _08369_ (.A(_01401_),
    .B(_01402_),
    .X(_01522_));
 sky130_fd_sc_hd__xor2_2 _08370_ (.A(_01521_),
    .B(_01522_),
    .X(_01523_));
 sky130_fd_sc_hd__nand4_1 _08371_ (.A(_01405_),
    .B(_01420_),
    .C(_01520_),
    .D(_01523_),
    .Y(_01524_));
 sky130_fd_sc_hd__xnor2_1 _08372_ (.A(_01511_),
    .B(_01512_),
    .Y(_01525_));
 sky130_fd_sc_hd__and2b_1 _08373_ (.A_N(_01461_),
    .B(_01462_),
    .X(_01526_));
 sky130_fd_sc_hd__nor2_1 _08374_ (.A(_01463_),
    .B(_01526_),
    .Y(_01527_));
 sky130_fd_sc_hd__nand2_1 _08375_ (.A(_01525_),
    .B(_01527_),
    .Y(_01528_));
 sky130_fd_sc_hd__a21o_1 _08376_ (.A1(_01491_),
    .A2(_01501_),
    .B1(_01500_),
    .X(_01529_));
 sky130_fd_sc_hd__o22a_1 _08377_ (.A1(net131),
    .A2(net164),
    .B1(net160),
    .B2(net83),
    .X(_01530_));
 sky130_fd_sc_hd__xnor2_1 _08378_ (.A(net159),
    .B(_01530_),
    .Y(_01531_));
 sky130_fd_sc_hd__o22a_1 _08379_ (.A1(net223),
    .A2(net79),
    .B1(net124),
    .B2(net162),
    .X(_01532_));
 sky130_fd_sc_hd__xor2_1 _08380_ (.A(net156),
    .B(_01532_),
    .X(_01533_));
 sky130_fd_sc_hd__or2_1 _08381_ (.A(_01531_),
    .B(_01533_),
    .X(_01534_));
 sky130_fd_sc_hd__o22a_1 _08382_ (.A1(net168),
    .A2(net89),
    .B1(net87),
    .B2(net166),
    .X(_01535_));
 sky130_fd_sc_hd__xor2_1 _08383_ (.A(net209),
    .B(_01535_),
    .X(_01536_));
 sky130_fd_sc_hd__nand2_2 _08384_ (.A(_06483_),
    .B(_00215_),
    .Y(_01537_));
 sky130_fd_sc_hd__a21o_1 _08385_ (.A1(_06456_),
    .A2(_06457_),
    .B1(net302),
    .X(_01538_));
 sky130_fd_sc_hd__a21o_1 _08386_ (.A1(_01537_),
    .A2(_01538_),
    .B1(net255),
    .X(_01539_));
 sky130_fd_sc_hd__nand3_1 _08387_ (.A(net255),
    .B(_01537_),
    .C(_01538_),
    .Y(_01540_));
 sky130_fd_sc_hd__and3_1 _08388_ (.A(_01536_),
    .B(_01539_),
    .C(_01540_),
    .X(_01541_));
 sky130_fd_sc_hd__o22a_1 _08389_ (.A1(net125),
    .A2(net171),
    .B1(net93),
    .B2(net173),
    .X(_01542_));
 sky130_fd_sc_hd__xnor2_1 _08390_ (.A(_00180_),
    .B(_01542_),
    .Y(_01543_));
 sky130_fd_sc_hd__a21o_1 _08391_ (.A1(_01539_),
    .A2(_01540_),
    .B1(_01536_),
    .X(_01544_));
 sky130_fd_sc_hd__and2b_1 _08392_ (.A_N(_01541_),
    .B(_01544_),
    .X(_01545_));
 sky130_fd_sc_hd__a21o_1 _08393_ (.A1(_01543_),
    .A2(_01544_),
    .B1(_01541_),
    .X(_01546_));
 sky130_fd_sc_hd__and2b_1 _08394_ (.A_N(_01534_),
    .B(_01546_),
    .X(_01547_));
 sky130_fd_sc_hd__o22a_1 _08395_ (.A1(net117),
    .A2(net148),
    .B1(net142),
    .B2(net115),
    .X(_01548_));
 sky130_fd_sc_hd__xnor2_1 _08396_ (.A(net181),
    .B(_01548_),
    .Y(_01549_));
 sky130_fd_sc_hd__o22a_1 _08397_ (.A1(net176),
    .A2(net145),
    .B1(net132),
    .B2(net174),
    .X(_01550_));
 sky130_fd_sc_hd__xnor2_1 _08398_ (.A(net188),
    .B(_01550_),
    .Y(_01551_));
 sky130_fd_sc_hd__o22a_1 _08399_ (.A1(net151),
    .A2(net146),
    .B1(net140),
    .B2(net153),
    .X(_01552_));
 sky130_fd_sc_hd__xnor2_1 _08400_ (.A(net192),
    .B(_01552_),
    .Y(_01553_));
 sky130_fd_sc_hd__xor2_1 _08401_ (.A(_01549_),
    .B(_01551_),
    .X(_01554_));
 sky130_fd_sc_hd__and2b_1 _08402_ (.A_N(_01553_),
    .B(_01554_),
    .X(_01555_));
 sky130_fd_sc_hd__o21ba_1 _08403_ (.A1(_01549_),
    .A2(_01551_),
    .B1_N(_01555_),
    .X(_01556_));
 sky130_fd_sc_hd__xnor2_1 _08404_ (.A(_01534_),
    .B(_01546_),
    .Y(_01557_));
 sky130_fd_sc_hd__and2b_1 _08405_ (.A_N(_01556_),
    .B(_01557_),
    .X(_01558_));
 sky130_fd_sc_hd__o211ai_2 _08406_ (.A1(_01547_),
    .A2(_01558_),
    .B1(_01502_),
    .C1(_01529_),
    .Y(_01559_));
 sky130_fd_sc_hd__xnor2_1 _08407_ (.A(_01483_),
    .B(_01484_),
    .Y(_01560_));
 sky130_fd_sc_hd__xnor2_1 _08408_ (.A(_01486_),
    .B(_01488_),
    .Y(_01561_));
 sky130_fd_sc_hd__and2_1 _08409_ (.A(_01560_),
    .B(_01561_),
    .X(_01562_));
 sky130_fd_sc_hd__xnor2_1 _08410_ (.A(_01497_),
    .B(_01499_),
    .Y(_01563_));
 sky130_fd_sc_hd__nor2_1 _08411_ (.A(_01560_),
    .B(_01561_),
    .Y(_01564_));
 sky130_fd_sc_hd__or2_1 _08412_ (.A(_01562_),
    .B(_01564_),
    .X(_01565_));
 sky130_fd_sc_hd__nor2_1 _08413_ (.A(_01563_),
    .B(_01565_),
    .Y(_01566_));
 sky130_fd_sc_hd__a211o_1 _08414_ (.A1(_01502_),
    .A2(_01529_),
    .B1(_01547_),
    .C1(_01558_),
    .X(_01567_));
 sky130_fd_sc_hd__o211ai_2 _08415_ (.A1(_01562_),
    .A2(_01566_),
    .B1(_01567_),
    .C1(_01559_),
    .Y(_01568_));
 sky130_fd_sc_hd__nand2_1 _08416_ (.A(_01559_),
    .B(_01568_),
    .Y(_01569_));
 sky130_fd_sc_hd__xor2_1 _08417_ (.A(_01525_),
    .B(_01527_),
    .X(_01570_));
 sky130_fd_sc_hd__nand2_1 _08418_ (.A(_01569_),
    .B(_01570_),
    .Y(_01571_));
 sky130_fd_sc_hd__xor2_1 _08419_ (.A(_01514_),
    .B(_01515_),
    .X(_01572_));
 sky130_fd_sc_hd__a21o_1 _08420_ (.A1(_01528_),
    .A2(_01571_),
    .B1(_01572_),
    .X(_01573_));
 sky130_fd_sc_hd__nand3_1 _08421_ (.A(_01528_),
    .B(_01571_),
    .C(_01572_),
    .Y(_01574_));
 sky130_fd_sc_hd__nand2_1 _08422_ (.A(_01573_),
    .B(_01574_),
    .Y(_01575_));
 sky130_fd_sc_hd__or2_1 _08423_ (.A(_01569_),
    .B(_01570_),
    .X(_01576_));
 sky130_fd_sc_hd__and2_1 _08424_ (.A(_01571_),
    .B(_01576_),
    .X(_01577_));
 sky130_fd_sc_hd__a211o_1 _08425_ (.A1(_01559_),
    .A2(_01567_),
    .B1(_01566_),
    .C1(_01562_),
    .X(_01578_));
 sky130_fd_sc_hd__a21o_1 _08426_ (.A1(_01506_),
    .A2(_01509_),
    .B1(_01508_),
    .X(_01579_));
 sky130_fd_sc_hd__and4_1 _08427_ (.A(_01510_),
    .B(_01568_),
    .C(_01578_),
    .D(_01579_),
    .X(_01580_));
 sky130_fd_sc_hd__o22a_1 _08428_ (.A1(net83),
    .A2(net162),
    .B1(net160),
    .B2(net131),
    .X(_01581_));
 sky130_fd_sc_hd__xnor2_1 _08429_ (.A(net159),
    .B(_01581_),
    .Y(_01582_));
 sky130_fd_sc_hd__nor2_1 _08430_ (.A(net223),
    .B(net124),
    .Y(_01583_));
 sky130_fd_sc_hd__xnor2_1 _08431_ (.A(net156),
    .B(_01583_),
    .Y(_01584_));
 sky130_fd_sc_hd__or2_1 _08432_ (.A(_01582_),
    .B(_01584_),
    .X(_01585_));
 sky130_fd_sc_hd__o22a_1 _08433_ (.A1(net168),
    .A2(net132),
    .B1(net89),
    .B2(net166),
    .X(_01586_));
 sky130_fd_sc_hd__xnor2_1 _08434_ (.A(net209),
    .B(_01586_),
    .Y(_01587_));
 sky130_fd_sc_hd__o22a_1 _08435_ (.A1(net301),
    .A2(net122),
    .B1(net252),
    .B2(net125),
    .X(_01588_));
 sky130_fd_sc_hd__xnor2_1 _08436_ (.A(net254),
    .B(_01588_),
    .Y(_01589_));
 sky130_fd_sc_hd__nor2_1 _08437_ (.A(_01587_),
    .B(_01589_),
    .Y(_01590_));
 sky130_fd_sc_hd__o22a_1 _08438_ (.A1(net170),
    .A2(net93),
    .B1(net87),
    .B2(net172),
    .X(_01591_));
 sky130_fd_sc_hd__xnor2_1 _08439_ (.A(_00180_),
    .B(_01591_),
    .Y(_01592_));
 sky130_fd_sc_hd__xor2_1 _08440_ (.A(_01587_),
    .B(_01589_),
    .X(_01593_));
 sky130_fd_sc_hd__a21oi_1 _08441_ (.A1(_01592_),
    .A2(_01593_),
    .B1(_01590_),
    .Y(_01594_));
 sky130_fd_sc_hd__nor2_1 _08442_ (.A(_01585_),
    .B(_01594_),
    .Y(_01595_));
 sky130_fd_sc_hd__o22a_1 _08443_ (.A1(net117),
    .A2(net164),
    .B1(net148),
    .B2(net115),
    .X(_01596_));
 sky130_fd_sc_hd__xnor2_1 _08444_ (.A(net181),
    .B(_01596_),
    .Y(_01597_));
 sky130_fd_sc_hd__o22a_1 _08445_ (.A1(net176),
    .A2(net146),
    .B1(net145),
    .B2(net174),
    .X(_01598_));
 sky130_fd_sc_hd__xnor2_1 _08446_ (.A(net188),
    .B(_01598_),
    .Y(_01599_));
 sky130_fd_sc_hd__o22a_1 _08447_ (.A1(net153),
    .A2(net142),
    .B1(net140),
    .B2(net151),
    .X(_01600_));
 sky130_fd_sc_hd__xnor2_1 _08448_ (.A(net192),
    .B(_01600_),
    .Y(_01601_));
 sky130_fd_sc_hd__xor2_1 _08449_ (.A(_01597_),
    .B(_01599_),
    .X(_01602_));
 sky130_fd_sc_hd__and2b_1 _08450_ (.A_N(_01601_),
    .B(_01602_),
    .X(_01603_));
 sky130_fd_sc_hd__o21ba_1 _08451_ (.A1(_01597_),
    .A2(_01599_),
    .B1_N(_01603_),
    .X(_01604_));
 sky130_fd_sc_hd__xnor2_1 _08452_ (.A(_01585_),
    .B(_01594_),
    .Y(_01605_));
 sky130_fd_sc_hd__nor2_1 _08453_ (.A(_01604_),
    .B(_01605_),
    .Y(_01606_));
 sky130_fd_sc_hd__xnor2_1 _08454_ (.A(_01556_),
    .B(_01557_),
    .Y(_01607_));
 sky130_fd_sc_hd__o21ai_1 _08455_ (.A1(_01595_),
    .A2(_01606_),
    .B1(_01607_),
    .Y(_01608_));
 sky130_fd_sc_hd__xnor2_1 _08456_ (.A(_01531_),
    .B(_01533_),
    .Y(_01609_));
 sky130_fd_sc_hd__inv_2 _08457_ (.A(_01609_),
    .Y(_01610_));
 sky130_fd_sc_hd__xor2_1 _08458_ (.A(_01543_),
    .B(_01545_),
    .X(_01611_));
 sky130_fd_sc_hd__and2_1 _08459_ (.A(_01610_),
    .B(_01611_),
    .X(_01612_));
 sky130_fd_sc_hd__xnor2_1 _08460_ (.A(_01553_),
    .B(_01554_),
    .Y(_01613_));
 sky130_fd_sc_hd__or2_1 _08461_ (.A(_01610_),
    .B(_01611_),
    .X(_01614_));
 sky130_fd_sc_hd__nand2b_1 _08462_ (.A_N(_01612_),
    .B(_01614_),
    .Y(_01615_));
 sky130_fd_sc_hd__a21o_1 _08463_ (.A1(_01613_),
    .A2(_01614_),
    .B1(_01612_),
    .X(_01616_));
 sky130_fd_sc_hd__or3_1 _08464_ (.A(_01595_),
    .B(_01606_),
    .C(_01607_),
    .X(_01617_));
 sky130_fd_sc_hd__and2_1 _08465_ (.A(_01608_),
    .B(_01617_),
    .X(_01618_));
 sky130_fd_sc_hd__nand2_1 _08466_ (.A(_01616_),
    .B(_01618_),
    .Y(_01619_));
 sky130_fd_sc_hd__a22oi_2 _08467_ (.A1(_01568_),
    .A2(_01578_),
    .B1(_01579_),
    .B2(_01510_),
    .Y(_01620_));
 sky130_fd_sc_hd__a211o_1 _08468_ (.A1(_01608_),
    .A2(_01619_),
    .B1(_01620_),
    .C1(_01580_),
    .X(_01621_));
 sky130_fd_sc_hd__and2b_1 _08469_ (.A_N(_01580_),
    .B(_01621_),
    .X(_01622_));
 sky130_fd_sc_hd__and2b_1 _08470_ (.A_N(_01622_),
    .B(_01577_),
    .X(_01623_));
 sky130_fd_sc_hd__xnor2_2 _08471_ (.A(_01577_),
    .B(_01622_),
    .Y(_01624_));
 sky130_fd_sc_hd__nand2b_1 _08472_ (.A_N(_01575_),
    .B(_01624_),
    .Y(_01625_));
 sky130_fd_sc_hd__xnor2_1 _08473_ (.A(_01616_),
    .B(_01618_),
    .Y(_01626_));
 sky130_fd_sc_hd__and2_1 _08474_ (.A(_01563_),
    .B(_01565_),
    .X(_01627_));
 sky130_fd_sc_hd__or2_1 _08475_ (.A(_01566_),
    .B(_01627_),
    .X(_01628_));
 sky130_fd_sc_hd__nor2_1 _08476_ (.A(_01626_),
    .B(_01628_),
    .Y(_01629_));
 sky130_fd_sc_hd__xnor2_1 _08477_ (.A(_01604_),
    .B(_01605_),
    .Y(_01630_));
 sky130_fd_sc_hd__o22a_1 _08478_ (.A1(net153),
    .A2(net148),
    .B1(net142),
    .B2(net151),
    .X(_01631_));
 sky130_fd_sc_hd__xnor2_1 _08479_ (.A(net192),
    .B(_01631_),
    .Y(_01632_));
 sky130_fd_sc_hd__o22a_1 _08480_ (.A1(net174),
    .A2(net146),
    .B1(net140),
    .B2(net176),
    .X(_01633_));
 sky130_fd_sc_hd__xnor2_1 _08481_ (.A(net188),
    .B(_01633_),
    .Y(_01634_));
 sky130_fd_sc_hd__nor2_1 _08482_ (.A(_01632_),
    .B(_01634_),
    .Y(_01635_));
 sky130_fd_sc_hd__o22a_1 _08483_ (.A1(net168),
    .A2(net145),
    .B1(net132),
    .B2(net166),
    .X(_01636_));
 sky130_fd_sc_hd__xnor2_1 _08484_ (.A(net209),
    .B(_01636_),
    .Y(_01637_));
 sky130_fd_sc_hd__o22a_1 _08485_ (.A1(net301),
    .A2(net125),
    .B1(net252),
    .B2(net93),
    .X(_01638_));
 sky130_fd_sc_hd__xnor2_1 _08486_ (.A(net254),
    .B(_01638_),
    .Y(_01639_));
 sky130_fd_sc_hd__or2_1 _08487_ (.A(_01637_),
    .B(_01639_),
    .X(_01640_));
 sky130_fd_sc_hd__o22a_1 _08488_ (.A1(net172),
    .A2(net89),
    .B1(net87),
    .B2(net170),
    .X(_01641_));
 sky130_fd_sc_hd__xnor2_1 _08489_ (.A(net207),
    .B(_01641_),
    .Y(_01642_));
 sky130_fd_sc_hd__xor2_1 _08490_ (.A(_01637_),
    .B(_01639_),
    .X(_01643_));
 sky130_fd_sc_hd__nand2b_1 _08491_ (.A_N(_01642_),
    .B(_01643_),
    .Y(_01644_));
 sky130_fd_sc_hd__xnor2_1 _08492_ (.A(net156),
    .B(_01635_),
    .Y(_01645_));
 sky130_fd_sc_hd__a21oi_1 _08493_ (.A1(_01640_),
    .A2(_01644_),
    .B1(_01645_),
    .Y(_01646_));
 sky130_fd_sc_hd__a21oi_1 _08494_ (.A1(net156),
    .A2(_01635_),
    .B1(_01646_),
    .Y(_01647_));
 sky130_fd_sc_hd__or2_1 _08495_ (.A(_01630_),
    .B(_01647_),
    .X(_01648_));
 sky130_fd_sc_hd__xnor2_1 _08496_ (.A(_01630_),
    .B(_01647_),
    .Y(_01649_));
 sky130_fd_sc_hd__xor2_1 _08497_ (.A(_01582_),
    .B(_01584_),
    .X(_01650_));
 sky130_fd_sc_hd__xor2_1 _08498_ (.A(_01592_),
    .B(_01593_),
    .X(_01651_));
 sky130_fd_sc_hd__nand2_1 _08499_ (.A(_01650_),
    .B(_01651_),
    .Y(_01652_));
 sky130_fd_sc_hd__xnor2_1 _08500_ (.A(_01601_),
    .B(_01602_),
    .Y(_01653_));
 sky130_fd_sc_hd__inv_2 _08501_ (.A(_01653_),
    .Y(_01654_));
 sky130_fd_sc_hd__or2_1 _08502_ (.A(_01650_),
    .B(_01651_),
    .X(_01655_));
 sky130_fd_sc_hd__nand2_1 _08503_ (.A(_01652_),
    .B(_01655_),
    .Y(_01656_));
 sky130_fd_sc_hd__o21a_1 _08504_ (.A1(_01654_),
    .A2(_01656_),
    .B1(_01652_),
    .X(_01657_));
 sky130_fd_sc_hd__o21ai_1 _08505_ (.A1(_01649_),
    .A2(_01657_),
    .B1(_01648_),
    .Y(_01658_));
 sky130_fd_sc_hd__and2_1 _08506_ (.A(_01626_),
    .B(_01628_),
    .X(_01659_));
 sky130_fd_sc_hd__nor2_1 _08507_ (.A(_01629_),
    .B(_01659_),
    .Y(_01660_));
 sky130_fd_sc_hd__a21oi_1 _08508_ (.A1(_01658_),
    .A2(_01660_),
    .B1(_01629_),
    .Y(_01661_));
 sky130_fd_sc_hd__o211ai_1 _08509_ (.A1(_01580_),
    .A2(_01620_),
    .B1(_01619_),
    .C1(_01608_),
    .Y(_01662_));
 sky130_fd_sc_hd__nand2_1 _08510_ (.A(_01621_),
    .B(_01662_),
    .Y(_01663_));
 sky130_fd_sc_hd__and2_1 _08511_ (.A(_01661_),
    .B(_01663_),
    .X(_01664_));
 sky130_fd_sc_hd__xnor2_1 _08512_ (.A(_01658_),
    .B(_01660_),
    .Y(_01665_));
 sky130_fd_sc_hd__xor2_1 _08513_ (.A(_01649_),
    .B(_01657_),
    .X(_01666_));
 sky130_fd_sc_hd__xnor2_1 _08514_ (.A(_01613_),
    .B(_01615_),
    .Y(_01667_));
 sky130_fd_sc_hd__nand2_1 _08515_ (.A(_01666_),
    .B(_01667_),
    .Y(_01668_));
 sky130_fd_sc_hd__or2_1 _08516_ (.A(_01666_),
    .B(_01667_),
    .X(_01669_));
 sky130_fd_sc_hd__nand2_1 _08517_ (.A(_01668_),
    .B(_01669_),
    .Y(_01670_));
 sky130_fd_sc_hd__and3_1 _08518_ (.A(_01640_),
    .B(_01644_),
    .C(_01645_),
    .X(_01671_));
 sky130_fd_sc_hd__nor2_1 _08519_ (.A(_01646_),
    .B(_01671_),
    .Y(_01672_));
 sky130_fd_sc_hd__o22a_1 _08520_ (.A1(net301),
    .A2(net93),
    .B1(net87),
    .B2(net252),
    .X(_01673_));
 sky130_fd_sc_hd__xnor2_1 _08521_ (.A(net254),
    .B(_01673_),
    .Y(_01674_));
 sky130_fd_sc_hd__o22a_1 _08522_ (.A1(net168),
    .A2(net146),
    .B1(net145),
    .B2(net166),
    .X(_01675_));
 sky130_fd_sc_hd__xnor2_1 _08523_ (.A(net209),
    .B(_01675_),
    .Y(_01676_));
 sky130_fd_sc_hd__or2_1 _08524_ (.A(_01674_),
    .B(_01676_),
    .X(_01677_));
 sky130_fd_sc_hd__o22a_1 _08525_ (.A1(net172),
    .A2(net132),
    .B1(net89),
    .B2(net170),
    .X(_01678_));
 sky130_fd_sc_hd__xnor2_1 _08526_ (.A(net207),
    .B(_01678_),
    .Y(_01679_));
 sky130_fd_sc_hd__and2_1 _08527_ (.A(_01674_),
    .B(_01676_),
    .X(_01680_));
 sky130_fd_sc_hd__xor2_1 _08528_ (.A(_01674_),
    .B(_01676_),
    .X(_01681_));
 sky130_fd_sc_hd__o21a_1 _08529_ (.A1(_01679_),
    .A2(_01680_),
    .B1(_01677_),
    .X(_01682_));
 sky130_fd_sc_hd__o22a_1 _08530_ (.A1(net115),
    .A2(net164),
    .B1(net160),
    .B2(net117),
    .X(_01683_));
 sky130_fd_sc_hd__xnor2_2 _08531_ (.A(net181),
    .B(_01683_),
    .Y(_01684_));
 sky130_fd_sc_hd__or2_1 _08532_ (.A(_01682_),
    .B(_01684_),
    .X(_01685_));
 sky130_fd_sc_hd__xnor2_2 _08533_ (.A(_01682_),
    .B(_01684_),
    .Y(_01686_));
 sky130_fd_sc_hd__o22a_1 _08534_ (.A1(net223),
    .A2(net83),
    .B1(net131),
    .B2(net162),
    .X(_01687_));
 sky130_fd_sc_hd__xnor2_2 _08535_ (.A(net159),
    .B(_01687_),
    .Y(_01688_));
 sky130_fd_sc_hd__o21a_1 _08536_ (.A1(_01686_),
    .A2(_01688_),
    .B1(_01685_),
    .X(_01689_));
 sky130_fd_sc_hd__and2b_1 _08537_ (.A_N(_01689_),
    .B(_01672_),
    .X(_01690_));
 sky130_fd_sc_hd__and2_1 _08538_ (.A(_01632_),
    .B(_01634_),
    .X(_01691_));
 sky130_fd_sc_hd__nor2_1 _08539_ (.A(_01635_),
    .B(_01691_),
    .Y(_01692_));
 sky130_fd_sc_hd__o22a_1 _08540_ (.A1(net153),
    .A2(net164),
    .B1(net148),
    .B2(net151),
    .X(_01693_));
 sky130_fd_sc_hd__xnor2_1 _08541_ (.A(net192),
    .B(_01693_),
    .Y(_01694_));
 sky130_fd_sc_hd__o22a_1 _08542_ (.A1(net176),
    .A2(net142),
    .B1(net140),
    .B2(net174),
    .X(_01695_));
 sky130_fd_sc_hd__xnor2_1 _08543_ (.A(net188),
    .B(_01695_),
    .Y(_01696_));
 sky130_fd_sc_hd__nor2_1 _08544_ (.A(_01694_),
    .B(_01696_),
    .Y(_01697_));
 sky130_fd_sc_hd__xor2_1 _08545_ (.A(_01642_),
    .B(_01643_),
    .X(_01698_));
 sky130_fd_sc_hd__xnor2_1 _08546_ (.A(_01692_),
    .B(_01697_),
    .Y(_01699_));
 sky130_fd_sc_hd__or2_1 _08547_ (.A(_01698_),
    .B(_01699_),
    .X(_01700_));
 sky130_fd_sc_hd__a21bo_1 _08548_ (.A1(_01692_),
    .A2(_01697_),
    .B1_N(_01700_),
    .X(_01701_));
 sky130_fd_sc_hd__xnor2_1 _08549_ (.A(_01672_),
    .B(_01689_),
    .Y(_01702_));
 sky130_fd_sc_hd__a21oi_1 _08550_ (.A1(_01701_),
    .A2(_01702_),
    .B1(_01690_),
    .Y(_01703_));
 sky130_fd_sc_hd__or2_1 _08551_ (.A(_01670_),
    .B(_01703_),
    .X(_01704_));
 sky130_fd_sc_hd__a21oi_1 _08552_ (.A1(_01668_),
    .A2(_01704_),
    .B1(_01665_),
    .Y(_01705_));
 sky130_fd_sc_hd__nor2_1 _08553_ (.A(_01661_),
    .B(_01663_),
    .Y(_01706_));
 sky130_fd_sc_hd__o21bai_2 _08554_ (.A1(_01705_),
    .A2(_01706_),
    .B1_N(_01664_),
    .Y(_01707_));
 sky130_fd_sc_hd__inv_2 _08555_ (.A(_01707_),
    .Y(_01708_));
 sky130_fd_sc_hd__nand2_1 _08556_ (.A(_01574_),
    .B(_01623_),
    .Y(_01709_));
 sky130_fd_sc_hd__o211ai_2 _08557_ (.A1(_01625_),
    .A2(_01707_),
    .B1(_01709_),
    .C1(_01573_),
    .Y(_01710_));
 sky130_fd_sc_hd__nand2_1 _08558_ (.A(_01670_),
    .B(_01703_),
    .Y(_01711_));
 sky130_fd_sc_hd__and2_1 _08559_ (.A(_01704_),
    .B(_01711_),
    .X(_01712_));
 sky130_fd_sc_hd__xnor2_1 _08560_ (.A(_01701_),
    .B(_01702_),
    .Y(_01713_));
 sky130_fd_sc_hd__xnor2_1 _08561_ (.A(_01654_),
    .B(_01656_),
    .Y(_01714_));
 sky130_fd_sc_hd__nor2_1 _08562_ (.A(_01713_),
    .B(_01714_),
    .Y(_01715_));
 sky130_fd_sc_hd__xor2_2 _08563_ (.A(_01686_),
    .B(_01688_),
    .X(_01716_));
 sky130_fd_sc_hd__inv_2 _08564_ (.A(_01716_),
    .Y(_01717_));
 sky130_fd_sc_hd__or2_1 _08565_ (.A(net223),
    .B(net131),
    .X(_01718_));
 sky130_fd_sc_hd__o22a_1 _08566_ (.A1(net117),
    .A2(net162),
    .B1(net160),
    .B2(net115),
    .X(_01719_));
 sky130_fd_sc_hd__xnor2_1 _08567_ (.A(net181),
    .B(_01719_),
    .Y(_01720_));
 sky130_fd_sc_hd__mux2_1 _08568_ (.A0(_01720_),
    .A1(net159),
    .S(_01718_),
    .X(_01721_));
 sky130_fd_sc_hd__xor2_1 _08569_ (.A(_01716_),
    .B(_01721_),
    .X(_01722_));
 sky130_fd_sc_hd__o22a_1 _08570_ (.A1(net252),
    .A2(net89),
    .B1(net87),
    .B2(net301),
    .X(_01723_));
 sky130_fd_sc_hd__xnor2_1 _08571_ (.A(net254),
    .B(_01723_),
    .Y(_01724_));
 sky130_fd_sc_hd__o22a_1 _08572_ (.A1(net172),
    .A2(net145),
    .B1(net132),
    .B2(net170),
    .X(_01725_));
 sky130_fd_sc_hd__xnor2_1 _08573_ (.A(net207),
    .B(_01725_),
    .Y(_01726_));
 sky130_fd_sc_hd__nor2_1 _08574_ (.A(_01724_),
    .B(_01726_),
    .Y(_01727_));
 sky130_fd_sc_hd__and2_1 _08575_ (.A(_01694_),
    .B(_01696_),
    .X(_01728_));
 sky130_fd_sc_hd__nor2_1 _08576_ (.A(_01697_),
    .B(_01728_),
    .Y(_01729_));
 sky130_fd_sc_hd__xnor2_1 _08577_ (.A(_01679_),
    .B(_01681_),
    .Y(_01730_));
 sky130_fd_sc_hd__inv_2 _08578_ (.A(_01730_),
    .Y(_01731_));
 sky130_fd_sc_hd__xnor2_1 _08579_ (.A(_01727_),
    .B(_01729_),
    .Y(_01732_));
 sky130_fd_sc_hd__nor2_1 _08580_ (.A(_01731_),
    .B(_01732_),
    .Y(_01733_));
 sky130_fd_sc_hd__a21oi_1 _08581_ (.A1(_01727_),
    .A2(_01729_),
    .B1(_01733_),
    .Y(_01734_));
 sky130_fd_sc_hd__or2_1 _08582_ (.A(_01722_),
    .B(_01734_),
    .X(_01735_));
 sky130_fd_sc_hd__o21a_1 _08583_ (.A1(_01717_),
    .A2(_01721_),
    .B1(_01735_),
    .X(_01736_));
 sky130_fd_sc_hd__and2_1 _08584_ (.A(_01713_),
    .B(_01714_),
    .X(_01737_));
 sky130_fd_sc_hd__nor2_1 _08585_ (.A(_01715_),
    .B(_01737_),
    .Y(_01738_));
 sky130_fd_sc_hd__and2b_1 _08586_ (.A_N(_01736_),
    .B(_01738_),
    .X(_01739_));
 sky130_fd_sc_hd__o21a_1 _08587_ (.A1(_01715_),
    .A2(_01739_),
    .B1(_01712_),
    .X(_01740_));
 sky130_fd_sc_hd__or3_1 _08588_ (.A(_01712_),
    .B(_01715_),
    .C(_01739_),
    .X(_01741_));
 sky130_fd_sc_hd__xnor2_1 _08589_ (.A(_01722_),
    .B(_01734_),
    .Y(_01742_));
 sky130_fd_sc_hd__nand2_1 _08590_ (.A(_01698_),
    .B(_01699_),
    .Y(_01743_));
 sky130_fd_sc_hd__nand2_1 _08591_ (.A(_01700_),
    .B(_01743_),
    .Y(_01744_));
 sky130_fd_sc_hd__nor2_1 _08592_ (.A(_01742_),
    .B(_01744_),
    .Y(_01745_));
 sky130_fd_sc_hd__xnor2_1 _08593_ (.A(_01742_),
    .B(_01744_),
    .Y(_01746_));
 sky130_fd_sc_hd__o22a_1 _08594_ (.A1(net166),
    .A2(net146),
    .B1(net140),
    .B2(net168),
    .X(_01747_));
 sky130_fd_sc_hd__xnor2_1 _08595_ (.A(net209),
    .B(_01747_),
    .Y(_01748_));
 sky130_fd_sc_hd__o22a_1 _08596_ (.A1(net151),
    .A2(net164),
    .B1(net160),
    .B2(net153),
    .X(_01749_));
 sky130_fd_sc_hd__xnor2_1 _08597_ (.A(net192),
    .B(_01749_),
    .Y(_01750_));
 sky130_fd_sc_hd__nor2_1 _08598_ (.A(_01748_),
    .B(_01750_),
    .Y(_01751_));
 sky130_fd_sc_hd__o22a_1 _08599_ (.A1(net176),
    .A2(net148),
    .B1(net142),
    .B2(net174),
    .X(_01752_));
 sky130_fd_sc_hd__xnor2_1 _08600_ (.A(net188),
    .B(_01752_),
    .Y(_01753_));
 sky130_fd_sc_hd__xnor2_1 _08601_ (.A(_01748_),
    .B(_01750_),
    .Y(_01754_));
 sky130_fd_sc_hd__nor2_1 _08602_ (.A(_01753_),
    .B(_01754_),
    .Y(_01755_));
 sky130_fd_sc_hd__xor2_1 _08603_ (.A(_01718_),
    .B(_01720_),
    .X(_01756_));
 sky130_fd_sc_hd__o21a_1 _08604_ (.A1(_01751_),
    .A2(_01755_),
    .B1(_01756_),
    .X(_01757_));
 sky130_fd_sc_hd__xnor2_1 _08605_ (.A(_01724_),
    .B(_01726_),
    .Y(_01758_));
 sky130_fd_sc_hd__o22a_1 _08606_ (.A1(net223),
    .A2(net117),
    .B1(net115),
    .B2(net162),
    .X(_01759_));
 sky130_fd_sc_hd__xnor2_1 _08607_ (.A(net181),
    .B(_01759_),
    .Y(_01760_));
 sky130_fd_sc_hd__o22a_1 _08608_ (.A1(net172),
    .A2(net146),
    .B1(net145),
    .B2(net170),
    .X(_01761_));
 sky130_fd_sc_hd__xnor2_2 _08609_ (.A(net207),
    .B(_01761_),
    .Y(_01762_));
 sky130_fd_sc_hd__o22a_1 _08610_ (.A1(net252),
    .A2(net132),
    .B1(net89),
    .B2(net301),
    .X(_01763_));
 sky130_fd_sc_hd__xnor2_2 _08611_ (.A(net254),
    .B(_01763_),
    .Y(_01764_));
 sky130_fd_sc_hd__or2_1 _08612_ (.A(_01762_),
    .B(_01764_),
    .X(_01765_));
 sky130_fd_sc_hd__xnor2_1 _08613_ (.A(_01758_),
    .B(_01760_),
    .Y(_01766_));
 sky130_fd_sc_hd__nor2_1 _08614_ (.A(_01765_),
    .B(_01766_),
    .Y(_01767_));
 sky130_fd_sc_hd__o21bai_1 _08615_ (.A1(_01758_),
    .A2(_01760_),
    .B1_N(_01767_),
    .Y(_01768_));
 sky130_fd_sc_hd__nor3_1 _08616_ (.A(_01751_),
    .B(_01755_),
    .C(_01756_),
    .Y(_01769_));
 sky130_fd_sc_hd__nor2_1 _08617_ (.A(_01757_),
    .B(_01769_),
    .Y(_01770_));
 sky130_fd_sc_hd__a21oi_1 _08618_ (.A1(_01768_),
    .A2(_01770_),
    .B1(_01757_),
    .Y(_01771_));
 sky130_fd_sc_hd__nor2_1 _08619_ (.A(_01746_),
    .B(_01771_),
    .Y(_01772_));
 sky130_fd_sc_hd__xnor2_1 _08620_ (.A(_01736_),
    .B(_01738_),
    .Y(_01773_));
 sky130_fd_sc_hd__o21a_1 _08621_ (.A1(_01745_),
    .A2(_01772_),
    .B1(_01773_),
    .X(_01774_));
 sky130_fd_sc_hd__or3_1 _08622_ (.A(_01745_),
    .B(_01772_),
    .C(_01773_),
    .X(_01775_));
 sky130_fd_sc_hd__and2_1 _08623_ (.A(_01746_),
    .B(_01771_),
    .X(_01776_));
 sky130_fd_sc_hd__nor2_1 _08624_ (.A(_01772_),
    .B(_01776_),
    .Y(_01777_));
 sky130_fd_sc_hd__xnor2_1 _08625_ (.A(_01768_),
    .B(_01770_),
    .Y(_01778_));
 sky130_fd_sc_hd__and2_1 _08626_ (.A(_01731_),
    .B(_01732_),
    .X(_01779_));
 sky130_fd_sc_hd__or2_1 _08627_ (.A(_01733_),
    .B(_01779_),
    .X(_01780_));
 sky130_fd_sc_hd__nor2_1 _08628_ (.A(_01778_),
    .B(_01780_),
    .Y(_01781_));
 sky130_fd_sc_hd__o22a_1 _08629_ (.A1(net168),
    .A2(net142),
    .B1(net140),
    .B2(net166),
    .X(_01782_));
 sky130_fd_sc_hd__xnor2_1 _08630_ (.A(net209),
    .B(_01782_),
    .Y(_01783_));
 sky130_fd_sc_hd__o22a_1 _08631_ (.A1(net153),
    .A2(net162),
    .B1(net160),
    .B2(net151),
    .X(_01784_));
 sky130_fd_sc_hd__xnor2_1 _08632_ (.A(net192),
    .B(_01784_),
    .Y(_01785_));
 sky130_fd_sc_hd__nor2_1 _08633_ (.A(_01783_),
    .B(_01785_),
    .Y(_01786_));
 sky130_fd_sc_hd__xnor2_1 _08634_ (.A(_01783_),
    .B(_01785_),
    .Y(_01787_));
 sky130_fd_sc_hd__o22a_1 _08635_ (.A1(net176),
    .A2(net164),
    .B1(net148),
    .B2(net174),
    .X(_01788_));
 sky130_fd_sc_hd__xnor2_1 _08636_ (.A(net188),
    .B(_01788_),
    .Y(_01789_));
 sky130_fd_sc_hd__nor2_1 _08637_ (.A(_01787_),
    .B(_01789_),
    .Y(_01790_));
 sky130_fd_sc_hd__xor2_1 _08638_ (.A(_01753_),
    .B(_01754_),
    .X(_01791_));
 sky130_fd_sc_hd__o21ai_1 _08639_ (.A1(_01786_),
    .A2(_01790_),
    .B1(_01791_),
    .Y(_01792_));
 sky130_fd_sc_hd__or3_1 _08640_ (.A(_01786_),
    .B(_01790_),
    .C(_01791_),
    .X(_01793_));
 sky130_fd_sc_hd__nand2_1 _08641_ (.A(_01792_),
    .B(_01793_),
    .Y(_01794_));
 sky130_fd_sc_hd__or2_1 _08642_ (.A(net223),
    .B(net115),
    .X(_01795_));
 sky130_fd_sc_hd__xor2_2 _08643_ (.A(_01762_),
    .B(_01764_),
    .X(_01796_));
 sky130_fd_sc_hd__inv_2 _08644_ (.A(_01796_),
    .Y(_01797_));
 sky130_fd_sc_hd__mux2_1 _08645_ (.A0(_01797_),
    .A1(net181),
    .S(_01795_),
    .X(_01798_));
 sky130_fd_sc_hd__o21ai_2 _08646_ (.A1(_01794_),
    .A2(_01798_),
    .B1(_01792_),
    .Y(_01799_));
 sky130_fd_sc_hd__nand2_1 _08647_ (.A(_01778_),
    .B(_01780_),
    .Y(_01800_));
 sky130_fd_sc_hd__nand2b_1 _08648_ (.A_N(_01781_),
    .B(_01800_),
    .Y(_01801_));
 sky130_fd_sc_hd__a21oi_2 _08649_ (.A1(_01799_),
    .A2(_01800_),
    .B1(_01781_),
    .Y(_01802_));
 sky130_fd_sc_hd__and2b_1 _08650_ (.A_N(_01802_),
    .B(_01777_),
    .X(_01803_));
 sky130_fd_sc_hd__xnor2_2 _08651_ (.A(_01777_),
    .B(_01802_),
    .Y(_01804_));
 sky130_fd_sc_hd__xnor2_1 _08652_ (.A(_01794_),
    .B(_01798_),
    .Y(_01805_));
 sky130_fd_sc_hd__and2_1 _08653_ (.A(_01765_),
    .B(_01766_),
    .X(_01806_));
 sky130_fd_sc_hd__or2_1 _08654_ (.A(_01767_),
    .B(_01806_),
    .X(_01807_));
 sky130_fd_sc_hd__xor2_1 _08655_ (.A(_01805_),
    .B(_01807_),
    .X(_01808_));
 sky130_fd_sc_hd__and2_1 _08656_ (.A(_01787_),
    .B(_01789_),
    .X(_01809_));
 sky130_fd_sc_hd__or2_1 _08657_ (.A(_01790_),
    .B(_01809_),
    .X(_01810_));
 sky130_fd_sc_hd__o22a_1 _08658_ (.A1(net168),
    .A2(net148),
    .B1(net142),
    .B2(net166),
    .X(_01811_));
 sky130_fd_sc_hd__xnor2_1 _08659_ (.A(net209),
    .B(_01811_),
    .Y(_01812_));
 sky130_fd_sc_hd__o22a_1 _08660_ (.A1(net252),
    .A2(net145),
    .B1(net132),
    .B2(net301),
    .X(_01813_));
 sky130_fd_sc_hd__xnor2_1 _08661_ (.A(net254),
    .B(_01813_),
    .Y(_01814_));
 sky130_fd_sc_hd__xor2_1 _08662_ (.A(_01812_),
    .B(_01814_),
    .X(_01815_));
 sky130_fd_sc_hd__o22a_1 _08663_ (.A1(net170),
    .A2(net146),
    .B1(net140),
    .B2(net172),
    .X(_01816_));
 sky130_fd_sc_hd__xnor2_1 _08664_ (.A(net207),
    .B(_01816_),
    .Y(_01817_));
 sky130_fd_sc_hd__inv_2 _08665_ (.A(_01817_),
    .Y(_01818_));
 sky130_fd_sc_hd__nand2_1 _08666_ (.A(_01815_),
    .B(_01818_),
    .Y(_01819_));
 sky130_fd_sc_hd__o21ai_1 _08667_ (.A1(_01812_),
    .A2(_01814_),
    .B1(_01819_),
    .Y(_01820_));
 sky130_fd_sc_hd__nand2b_1 _08668_ (.A_N(_01810_),
    .B(_01820_),
    .Y(_01821_));
 sky130_fd_sc_hd__xor2_1 _08669_ (.A(_01810_),
    .B(_01820_),
    .X(_01822_));
 sky130_fd_sc_hd__o22a_1 _08670_ (.A1(net223),
    .A2(net153),
    .B1(net151),
    .B2(net162),
    .X(_01823_));
 sky130_fd_sc_hd__xnor2_1 _08671_ (.A(net192),
    .B(_01823_),
    .Y(_01824_));
 sky130_fd_sc_hd__o22a_1 _08672_ (.A1(net174),
    .A2(net164),
    .B1(net160),
    .B2(net176),
    .X(_01825_));
 sky130_fd_sc_hd__xnor2_1 _08673_ (.A(net188),
    .B(_01825_),
    .Y(_01826_));
 sky130_fd_sc_hd__nor2_1 _08674_ (.A(_01824_),
    .B(_01826_),
    .Y(_01827_));
 sky130_fd_sc_hd__o31a_1 _08675_ (.A1(_01822_),
    .A2(_01824_),
    .A3(_01826_),
    .B1(_01821_),
    .X(_01828_));
 sky130_fd_sc_hd__nand2b_1 _08676_ (.A_N(_01828_),
    .B(_01808_),
    .Y(_01829_));
 sky130_fd_sc_hd__o21a_1 _08677_ (.A1(_01805_),
    .A2(_01807_),
    .B1(_01829_),
    .X(_01830_));
 sky130_fd_sc_hd__xnor2_2 _08678_ (.A(_01799_),
    .B(_01801_),
    .Y(_01831_));
 sky130_fd_sc_hd__and2b_1 _08679_ (.A_N(_01830_),
    .B(_01831_),
    .X(_01832_));
 sky130_fd_sc_hd__xnor2_2 _08680_ (.A(_01830_),
    .B(_01831_),
    .Y(_01833_));
 sky130_fd_sc_hd__xor2_1 _08681_ (.A(_01808_),
    .B(_01828_),
    .X(_01834_));
 sky130_fd_sc_hd__xnor2_1 _08682_ (.A(_01822_),
    .B(_01827_),
    .Y(_01835_));
 sky130_fd_sc_hd__xnor2_1 _08683_ (.A(_01795_),
    .B(_01796_),
    .Y(_01836_));
 sky130_fd_sc_hd__nand2_1 _08684_ (.A(_01835_),
    .B(_01836_),
    .Y(_01837_));
 sky130_fd_sc_hd__or2_1 _08685_ (.A(_01815_),
    .B(_01818_),
    .X(_01838_));
 sky130_fd_sc_hd__nand2_1 _08686_ (.A(_01819_),
    .B(_01838_),
    .Y(_01839_));
 sky130_fd_sc_hd__o22a_1 _08687_ (.A1(net168),
    .A2(net164),
    .B1(net148),
    .B2(net166),
    .X(_01840_));
 sky130_fd_sc_hd__xnor2_1 _08688_ (.A(net211),
    .B(_01840_),
    .Y(_01841_));
 sky130_fd_sc_hd__o22a_1 _08689_ (.A1(net252),
    .A2(net146),
    .B1(net145),
    .B2(net301),
    .X(_01842_));
 sky130_fd_sc_hd__xnor2_1 _08690_ (.A(net254),
    .B(_01842_),
    .Y(_01843_));
 sky130_fd_sc_hd__o22a_1 _08691_ (.A1(net172),
    .A2(net142),
    .B1(net140),
    .B2(net170),
    .X(_01844_));
 sky130_fd_sc_hd__xnor2_1 _08692_ (.A(net207),
    .B(_01844_),
    .Y(_01845_));
 sky130_fd_sc_hd__xor2_1 _08693_ (.A(_01841_),
    .B(_01843_),
    .X(_01846_));
 sky130_fd_sc_hd__nand2b_1 _08694_ (.A_N(_01845_),
    .B(_01846_),
    .Y(_01847_));
 sky130_fd_sc_hd__o21a_1 _08695_ (.A1(_01841_),
    .A2(_01843_),
    .B1(_01847_),
    .X(_01848_));
 sky130_fd_sc_hd__xnor2_1 _08696_ (.A(_01839_),
    .B(_01848_),
    .Y(_01849_));
 sky130_fd_sc_hd__o22a_1 _08697_ (.A1(net176),
    .A2(net162),
    .B1(net160),
    .B2(net174),
    .X(_01850_));
 sky130_fd_sc_hd__xor2_1 _08698_ (.A(net190),
    .B(_01850_),
    .X(_01851_));
 sky130_fd_sc_hd__o21a_1 _08699_ (.A1(net223),
    .A2(net151),
    .B1(_06490_),
    .X(_01852_));
 sky130_fd_sc_hd__and3_2 _08700_ (.A(net227),
    .B(net191),
    .C(_00138_),
    .X(_01853_));
 sky130_fd_sc_hd__o21ai_2 _08701_ (.A1(_01852_),
    .A2(_01853_),
    .B1(_01851_),
    .Y(_01854_));
 sky130_fd_sc_hd__nor2_1 _08702_ (.A(_01849_),
    .B(_01854_),
    .Y(_01855_));
 sky130_fd_sc_hd__o21bai_1 _08703_ (.A1(_01839_),
    .A2(_01848_),
    .B1_N(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__xor2_1 _08704_ (.A(_01835_),
    .B(_01836_),
    .X(_01857_));
 sky130_fd_sc_hd__nand2_1 _08705_ (.A(_01856_),
    .B(_01857_),
    .Y(_01858_));
 sky130_fd_sc_hd__and3_1 _08706_ (.A(_01834_),
    .B(_01837_),
    .C(_01858_),
    .X(_01859_));
 sky130_fd_sc_hd__xor2_1 _08707_ (.A(_01849_),
    .B(_01854_),
    .X(_01860_));
 sky130_fd_sc_hd__and2_1 _08708_ (.A(_01824_),
    .B(_01826_),
    .X(_01861_));
 sky130_fd_sc_hd__nor2_1 _08709_ (.A(_01827_),
    .B(_01861_),
    .Y(_01862_));
 sky130_fd_sc_hd__nand2_1 _08710_ (.A(_01860_),
    .B(_01862_),
    .Y(_01863_));
 sky130_fd_sc_hd__xnor2_1 _08711_ (.A(_01860_),
    .B(_01862_),
    .Y(_01864_));
 sky130_fd_sc_hd__xnor2_1 _08712_ (.A(_01845_),
    .B(_01846_),
    .Y(_01865_));
 sky130_fd_sc_hd__nand2_1 _08713_ (.A(_06490_),
    .B(_01865_),
    .Y(_01866_));
 sky130_fd_sc_hd__xnor2_1 _08714_ (.A(net192),
    .B(_01865_),
    .Y(_01867_));
 sky130_fd_sc_hd__o22a_1 _08715_ (.A1(net301),
    .A2(net146),
    .B1(net140),
    .B2(net252),
    .X(_01868_));
 sky130_fd_sc_hd__xnor2_1 _08716_ (.A(net254),
    .B(_01868_),
    .Y(_01869_));
 sky130_fd_sc_hd__o22a_1 _08717_ (.A1(net172),
    .A2(net148),
    .B1(net142),
    .B2(net170),
    .X(_01870_));
 sky130_fd_sc_hd__xnor2_1 _08718_ (.A(net207),
    .B(_01870_),
    .Y(_01871_));
 sky130_fd_sc_hd__nor2_1 _08719_ (.A(_01869_),
    .B(_01871_),
    .Y(_01872_));
 sky130_fd_sc_hd__a21bo_1 _08720_ (.A1(_01867_),
    .A2(_01872_),
    .B1_N(_01866_),
    .X(_01873_));
 sky130_fd_sc_hd__nand2b_1 _08721_ (.A_N(_01864_),
    .B(_01873_),
    .Y(_01874_));
 sky130_fd_sc_hd__xnor2_1 _08722_ (.A(_01856_),
    .B(_01857_),
    .Y(_01875_));
 sky130_fd_sc_hd__a21oi_1 _08723_ (.A1(_01863_),
    .A2(_01874_),
    .B1(_01875_),
    .Y(_01876_));
 sky130_fd_sc_hd__a21o_1 _08724_ (.A1(_01863_),
    .A2(_01874_),
    .B1(_01875_),
    .X(_01877_));
 sky130_fd_sc_hd__a21o_1 _08725_ (.A1(_01837_),
    .A2(_01858_),
    .B1(_01834_),
    .X(_01878_));
 sky130_fd_sc_hd__and3_1 _08726_ (.A(_01863_),
    .B(_01874_),
    .C(_01875_),
    .X(_01879_));
 sky130_fd_sc_hd__nor2_1 _08727_ (.A(_01876_),
    .B(_01879_),
    .Y(_01880_));
 sky130_fd_sc_hd__xor2_1 _08728_ (.A(_01864_),
    .B(_01873_),
    .X(_01881_));
 sky130_fd_sc_hd__xnor2_1 _08729_ (.A(_01867_),
    .B(_01872_),
    .Y(_01882_));
 sky130_fd_sc_hd__or3_1 _08730_ (.A(_01851_),
    .B(_01852_),
    .C(_01853_),
    .X(_01883_));
 sky130_fd_sc_hd__nand2_1 _08731_ (.A(_01854_),
    .B(_01883_),
    .Y(_01884_));
 sky130_fd_sc_hd__xnor2_1 _08732_ (.A(_01882_),
    .B(_01884_),
    .Y(_01885_));
 sky130_fd_sc_hd__o22a_1 _08733_ (.A1(net172),
    .A2(net164),
    .B1(net148),
    .B2(net170),
    .X(_01886_));
 sky130_fd_sc_hd__xnor2_2 _08734_ (.A(net207),
    .B(_01886_),
    .Y(_01887_));
 sky130_fd_sc_hd__o22a_1 _08735_ (.A1(net252),
    .A2(net142),
    .B1(net140),
    .B2(net301),
    .X(_01888_));
 sky130_fd_sc_hd__xnor2_2 _08736_ (.A(net254),
    .B(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__o22a_1 _08737_ (.A1(net166),
    .A2(net164),
    .B1(net160),
    .B2(net168),
    .X(_01890_));
 sky130_fd_sc_hd__xor2_1 _08738_ (.A(net209),
    .B(_01890_),
    .X(_01891_));
 sky130_fd_sc_hd__or3b_1 _08739_ (.A(_01887_),
    .B(_01889_),
    .C_N(_01891_),
    .X(_01892_));
 sky130_fd_sc_hd__o22a_1 _08740_ (.A1(net223),
    .A2(net176),
    .B1(net174),
    .B2(net162),
    .X(_01893_));
 sky130_fd_sc_hd__xor2_1 _08741_ (.A(net188),
    .B(_01893_),
    .X(_01894_));
 sky130_fd_sc_hd__o21bai_1 _08742_ (.A1(_01887_),
    .A2(_01889_),
    .B1_N(_01891_),
    .Y(_01895_));
 sky130_fd_sc_hd__nand3_1 _08743_ (.A(_01892_),
    .B(_01894_),
    .C(_01895_),
    .Y(_01896_));
 sky130_fd_sc_hd__nand2_1 _08744_ (.A(_01892_),
    .B(_01896_),
    .Y(_01897_));
 sky130_fd_sc_hd__and2b_1 _08745_ (.A_N(_01885_),
    .B(_01897_),
    .X(_01898_));
 sky130_fd_sc_hd__o21bai_1 _08746_ (.A1(_01882_),
    .A2(_01884_),
    .B1_N(_01898_),
    .Y(_01899_));
 sky130_fd_sc_hd__and2b_1 _08747_ (.A_N(_01881_),
    .B(_01899_),
    .X(_01900_));
 sky130_fd_sc_hd__xnor2_1 _08748_ (.A(_01881_),
    .B(_01899_),
    .Y(_01901_));
 sky130_fd_sc_hd__xnor2_1 _08749_ (.A(_01885_),
    .B(_01897_),
    .Y(_01902_));
 sky130_fd_sc_hd__a21o_1 _08750_ (.A1(_01892_),
    .A2(_01895_),
    .B1(_01894_),
    .X(_01903_));
 sky130_fd_sc_hd__and2_1 _08751_ (.A(_01869_),
    .B(_01871_),
    .X(_01904_));
 sky130_fd_sc_hd__nor2_1 _08752_ (.A(_01872_),
    .B(_01904_),
    .Y(_01905_));
 sky130_fd_sc_hd__and3_1 _08753_ (.A(_01896_),
    .B(_01903_),
    .C(_01905_),
    .X(_01906_));
 sky130_fd_sc_hd__a21oi_1 _08754_ (.A1(_01896_),
    .A2(_01903_),
    .B1(_01905_),
    .Y(_01907_));
 sky130_fd_sc_hd__or2_1 _08755_ (.A(net223),
    .B(net174),
    .X(_01908_));
 sky130_fd_sc_hd__o22a_1 _08756_ (.A1(net168),
    .A2(net162),
    .B1(net160),
    .B2(net166),
    .X(_01909_));
 sky130_fd_sc_hd__xnor2_2 _08757_ (.A(net209),
    .B(_01909_),
    .Y(_01910_));
 sky130_fd_sc_hd__mux2_1 _08758_ (.A0(_01910_),
    .A1(net188),
    .S(_01908_),
    .X(_01911_));
 sky130_fd_sc_hd__or3_1 _08759_ (.A(_01906_),
    .B(_01907_),
    .C(_01911_),
    .X(_01912_));
 sky130_fd_sc_hd__and2b_1 _08760_ (.A_N(_01906_),
    .B(_01912_),
    .X(_01913_));
 sky130_fd_sc_hd__and2b_1 _08761_ (.A_N(_01913_),
    .B(_01902_),
    .X(_01914_));
 sky130_fd_sc_hd__xnor2_1 _08762_ (.A(_01902_),
    .B(_01913_),
    .Y(_01915_));
 sky130_fd_sc_hd__xor2_2 _08763_ (.A(_01887_),
    .B(_01889_),
    .X(_01916_));
 sky130_fd_sc_hd__xor2_2 _08764_ (.A(_01908_),
    .B(_01910_),
    .X(_01917_));
 sky130_fd_sc_hd__or3_2 _08765_ (.A(net253),
    .B(_00260_),
    .C(_00262_),
    .X(_01918_));
 sky130_fd_sc_hd__a21o_1 _08766_ (.A1(_00297_),
    .A2(_00298_),
    .B1(net302),
    .X(_01919_));
 sky130_fd_sc_hd__a21o_1 _08767_ (.A1(_01918_),
    .A2(_01919_),
    .B1(net255),
    .X(_01920_));
 sky130_fd_sc_hd__nand3_2 _08768_ (.A(net255),
    .B(_01918_),
    .C(_01919_),
    .Y(_01921_));
 sky130_fd_sc_hd__o22a_1 _08769_ (.A1(net171),
    .A2(net165),
    .B1(net161),
    .B2(net173),
    .X(_01922_));
 sky130_fd_sc_hd__xnor2_1 _08770_ (.A(net208),
    .B(_01922_),
    .Y(_01923_));
 sky130_fd_sc_hd__nand3b_4 _08771_ (.A_N(_01923_),
    .B(_01921_),
    .C(_01920_),
    .Y(_01924_));
 sky130_fd_sc_hd__xor2_2 _08772_ (.A(_01916_),
    .B(_01917_),
    .X(_01925_));
 sky130_fd_sc_hd__and2b_1 _08773_ (.A_N(_01924_),
    .B(_01925_),
    .X(_01926_));
 sky130_fd_sc_hd__a21o_1 _08774_ (.A1(_01916_),
    .A2(_01917_),
    .B1(_01926_),
    .X(_01927_));
 sky130_fd_sc_hd__o21ai_1 _08775_ (.A1(_01906_),
    .A2(_01907_),
    .B1(_01911_),
    .Y(_01928_));
 sky130_fd_sc_hd__nand3_1 _08776_ (.A(_01912_),
    .B(_01927_),
    .C(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__a21oi_1 _08777_ (.A1(_01912_),
    .A2(_01928_),
    .B1(_01927_),
    .Y(_01930_));
 sky130_fd_sc_hd__a21o_1 _08778_ (.A1(_01912_),
    .A2(_01928_),
    .B1(_01927_),
    .X(_01931_));
 sky130_fd_sc_hd__and2_1 _08779_ (.A(_01929_),
    .B(_01931_),
    .X(_01932_));
 sky130_fd_sc_hd__xor2_2 _08780_ (.A(_01924_),
    .B(_01925_),
    .X(_01933_));
 sky130_fd_sc_hd__a21bo_1 _08781_ (.A1(_01920_),
    .A2(_01921_),
    .B1_N(_01923_),
    .X(_01934_));
 sky130_fd_sc_hd__o22a_1 _08782_ (.A1(net223),
    .A2(net168),
    .B1(net167),
    .B2(net162),
    .X(_01935_));
 sky130_fd_sc_hd__xor2_1 _08783_ (.A(net209),
    .B(_01935_),
    .X(_01936_));
 sky130_fd_sc_hd__and3_1 _08784_ (.A(_01924_),
    .B(_01934_),
    .C(_01936_),
    .X(_01937_));
 sky130_fd_sc_hd__o22a_1 _08785_ (.A1(net173),
    .A2(net163),
    .B1(net160),
    .B2(net171),
    .X(_01938_));
 sky130_fd_sc_hd__xnor2_1 _08786_ (.A(net208),
    .B(_01938_),
    .Y(_01939_));
 sky130_fd_sc_hd__o32a_2 _08787_ (.A1(_04416_),
    .A2(_00260_),
    .A3(_00262_),
    .B1(net253),
    .B2(net165),
    .X(_01940_));
 sky130_fd_sc_hd__xnor2_1 _08788_ (.A(net254),
    .B(_01940_),
    .Y(_01941_));
 sky130_fd_sc_hd__nor2_1 _08789_ (.A(_01939_),
    .B(_01941_),
    .Y(_01942_));
 sky130_fd_sc_hd__inv_2 _08790_ (.A(_01942_),
    .Y(_01943_));
 sky130_fd_sc_hd__a21oi_1 _08791_ (.A1(_01924_),
    .A2(_01934_),
    .B1(_01936_),
    .Y(_01944_));
 sky130_fd_sc_hd__or3_1 _08792_ (.A(_01937_),
    .B(_01943_),
    .C(_01944_),
    .X(_01945_));
 sky130_fd_sc_hd__nand2b_1 _08793_ (.A_N(_01937_),
    .B(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__and2b_1 _08794_ (.A_N(_01933_),
    .B(_01946_),
    .X(_01947_));
 sky130_fd_sc_hd__xor2_1 _08795_ (.A(_01933_),
    .B(_01946_),
    .X(_01948_));
 sky130_fd_sc_hd__o21ai_1 _08796_ (.A1(_01937_),
    .A2(_01944_),
    .B1(_01943_),
    .Y(_01949_));
 sky130_fd_sc_hd__nand2_1 _08797_ (.A(_01945_),
    .B(_01949_),
    .Y(_01950_));
 sky130_fd_sc_hd__or2_1 _08798_ (.A(net225),
    .B(net167),
    .X(_01951_));
 sky130_fd_sc_hd__xor2_1 _08799_ (.A(_01939_),
    .B(_01941_),
    .X(_01952_));
 sky130_fd_sc_hd__nor2_1 _08800_ (.A(_01951_),
    .B(_01952_),
    .Y(_01953_));
 sky130_fd_sc_hd__and2_1 _08801_ (.A(net209),
    .B(_01951_),
    .X(_01954_));
 sky130_fd_sc_hd__nor2_1 _08802_ (.A(_01953_),
    .B(_01954_),
    .Y(_01955_));
 sky130_fd_sc_hd__or3_1 _08803_ (.A(_01950_),
    .B(_01953_),
    .C(_01954_),
    .X(_01956_));
 sky130_fd_sc_hd__xor2_1 _08804_ (.A(_01950_),
    .B(_01955_),
    .X(_01957_));
 sky130_fd_sc_hd__o22a_1 _08805_ (.A1(net302),
    .A2(net165),
    .B1(net160),
    .B2(net252),
    .X(_01958_));
 sky130_fd_sc_hd__xnor2_1 _08806_ (.A(net255),
    .B(_01958_),
    .Y(_01959_));
 sky130_fd_sc_hd__o22a_1 _08807_ (.A1(net225),
    .A2(net172),
    .B1(net171),
    .B2(net163),
    .X(_01960_));
 sky130_fd_sc_hd__xnor2_1 _08808_ (.A(net208),
    .B(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__nor2_1 _08809_ (.A(_01959_),
    .B(_01961_),
    .Y(_01962_));
 sky130_fd_sc_hd__xnor2_1 _08810_ (.A(_01951_),
    .B(_01952_),
    .Y(_01963_));
 sky130_fd_sc_hd__xor2_1 _08811_ (.A(_01962_),
    .B(_01963_),
    .X(_01964_));
 sky130_fd_sc_hd__xnor2_1 _08812_ (.A(_01959_),
    .B(_01961_),
    .Y(_01965_));
 sky130_fd_sc_hd__o22a_1 _08813_ (.A1(net252),
    .A2(net163),
    .B1(net160),
    .B2(net302),
    .X(_01966_));
 sky130_fd_sc_hd__xnor2_2 _08814_ (.A(net254),
    .B(_01966_),
    .Y(_01967_));
 sky130_fd_sc_hd__or2_1 _08815_ (.A(net225),
    .B(net170),
    .X(_01968_));
 sky130_fd_sc_hd__xnor2_1 _08816_ (.A(net208),
    .B(_01968_),
    .Y(_01969_));
 sky130_fd_sc_hd__or2_1 _08817_ (.A(_01967_),
    .B(_01969_),
    .X(_01970_));
 sky130_fd_sc_hd__nor2_1 _08818_ (.A(_01965_),
    .B(_01970_),
    .Y(_01971_));
 sky130_fd_sc_hd__xnor2_1 _08819_ (.A(_01965_),
    .B(_01970_),
    .Y(_01972_));
 sky130_fd_sc_hd__xor2_1 _08820_ (.A(_01967_),
    .B(_01969_),
    .X(_01973_));
 sky130_fd_sc_hd__xor2_2 _08821_ (.A(_01967_),
    .B(_01968_),
    .X(_01974_));
 sky130_fd_sc_hd__a22o_1 _08822_ (.A1(_06308_),
    .A2(_00215_),
    .B1(_00338_),
    .B2(net304),
    .X(_01975_));
 sky130_fd_sc_hd__nand2b_2 _08823_ (.A_N(_01975_),
    .B(_06371_),
    .Y(_01976_));
 sky130_fd_sc_hd__nor2_1 _08824_ (.A(net255),
    .B(_01976_),
    .Y(_01977_));
 sky130_fd_sc_hd__a22oi_1 _08825_ (.A1(_00180_),
    .A2(_01973_),
    .B1(_01974_),
    .B2(_01977_),
    .Y(_01978_));
 sky130_fd_sc_hd__nor2_1 _08826_ (.A(_01972_),
    .B(_01978_),
    .Y(_01979_));
 sky130_fd_sc_hd__o21ai_1 _08827_ (.A1(_01971_),
    .A2(_01979_),
    .B1(_01964_),
    .Y(_01980_));
 sky130_fd_sc_hd__a21boi_1 _08828_ (.A1(_01962_),
    .A2(_01963_),
    .B1_N(_01980_),
    .Y(_01981_));
 sky130_fd_sc_hd__o21a_1 _08829_ (.A1(_01957_),
    .A2(_01981_),
    .B1(_01956_),
    .X(_01982_));
 sky130_fd_sc_hd__o21ba_1 _08830_ (.A1(_01948_),
    .A2(_01982_),
    .B1_N(_01947_),
    .X(_01983_));
 sky130_fd_sc_hd__o21ai_1 _08831_ (.A1(_01930_),
    .A2(_01983_),
    .B1(_01929_),
    .Y(_01984_));
 sky130_fd_sc_hd__a21o_1 _08832_ (.A1(_01915_),
    .A2(_01984_),
    .B1(_01914_),
    .X(_01985_));
 sky130_fd_sc_hd__a21o_1 _08833_ (.A1(_01901_),
    .A2(_01985_),
    .B1(_01900_),
    .X(_01986_));
 sky130_fd_sc_hd__a21oi_1 _08834_ (.A1(_01877_),
    .A2(_01878_),
    .B1(_01859_),
    .Y(_01987_));
 sky130_fd_sc_hd__and2b_1 _08835_ (.A_N(_01859_),
    .B(_01878_),
    .X(_01988_));
 sky130_fd_sc_hd__a31o_1 _08836_ (.A1(_01880_),
    .A2(_01986_),
    .A3(_01988_),
    .B1(_01987_),
    .X(_01989_));
 sky130_fd_sc_hd__a21o_1 _08837_ (.A1(_01833_),
    .A2(_01989_),
    .B1(_01832_),
    .X(_01990_));
 sky130_fd_sc_hd__a21o_1 _08838_ (.A1(_01804_),
    .A2(_01990_),
    .B1(_01803_),
    .X(_01991_));
 sky130_fd_sc_hd__a21o_1 _08839_ (.A1(_01775_),
    .A2(_01991_),
    .B1(_01774_),
    .X(_01992_));
 sky130_fd_sc_hd__a21o_2 _08840_ (.A1(_01741_),
    .A2(_01992_),
    .B1(_01740_),
    .X(_01993_));
 sky130_fd_sc_hd__and3_1 _08841_ (.A(_01665_),
    .B(_01668_),
    .C(_01704_),
    .X(_01994_));
 sky130_fd_sc_hd__nor2_1 _08842_ (.A(_01705_),
    .B(_01994_),
    .Y(_01995_));
 sky130_fd_sc_hd__nor2_1 _08843_ (.A(_01664_),
    .B(_01706_),
    .Y(_01996_));
 sky130_fd_sc_hd__and3b_1 _08844_ (.A_N(_01625_),
    .B(_01995_),
    .C(_01996_),
    .X(_01997_));
 sky130_fd_sc_hd__a21o_1 _08845_ (.A1(_01993_),
    .A2(_01997_),
    .B1(_01710_),
    .X(_01998_));
 sky130_fd_sc_hd__nand2b_1 _08846_ (.A_N(_01524_),
    .B(_01710_),
    .Y(_01999_));
 sky130_fd_sc_hd__nand3b_2 _08847_ (.A_N(_01524_),
    .B(_01993_),
    .C(_01997_),
    .Y(_02000_));
 sky130_fd_sc_hd__a21o_1 _08848_ (.A1(_01521_),
    .A2(_01522_),
    .B1(_01518_),
    .X(_02001_));
 sky130_fd_sc_hd__o21a_1 _08849_ (.A1(_01521_),
    .A2(_01522_),
    .B1(_02001_),
    .X(_02002_));
 sky130_fd_sc_hd__a211o_1 _08850_ (.A1(_01406_),
    .A2(_01419_),
    .B1(_01356_),
    .C1(_01403_),
    .X(_02003_));
 sky130_fd_sc_hd__o21ai_2 _08851_ (.A1(_01406_),
    .A2(_01419_),
    .B1(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__a31oi_4 _08852_ (.A1(_01405_),
    .A2(_01420_),
    .A3(_02002_),
    .B1(_02004_),
    .Y(_02005_));
 sky130_fd_sc_hd__xnor2_2 _08853_ (.A(_01186_),
    .B(_01187_),
    .Y(_02006_));
 sky130_fd_sc_hd__a21oi_1 _08854_ (.A1(_01115_),
    .A2(_01117_),
    .B1(_01116_),
    .Y(_02007_));
 sky130_fd_sc_hd__nor2_2 _08855_ (.A(_01118_),
    .B(_02007_),
    .Y(_02008_));
 sky130_fd_sc_hd__nand2_1 _08856_ (.A(_02006_),
    .B(_02008_),
    .Y(_02009_));
 sky130_fd_sc_hd__nand2_1 _08857_ (.A(_01411_),
    .B(_01413_),
    .Y(_02010_));
 sky130_fd_sc_hd__xnor2_1 _08858_ (.A(_02006_),
    .B(_02008_),
    .Y(_02011_));
 sky130_fd_sc_hd__nand2b_1 _08859_ (.A_N(_02011_),
    .B(_02010_),
    .Y(_02012_));
 sky130_fd_sc_hd__xnor2_1 _08860_ (.A(_01189_),
    .B(_01190_),
    .Y(_02013_));
 sky130_fd_sc_hd__and3_1 _08861_ (.A(_02009_),
    .B(_02012_),
    .C(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__a21o_1 _08862_ (.A1(_02009_),
    .A2(_02012_),
    .B1(_02013_),
    .X(_02015_));
 sky130_fd_sc_hd__and2b_1 _08863_ (.A_N(_02014_),
    .B(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__nand2_1 _08864_ (.A(_01416_),
    .B(_01418_),
    .Y(_02017_));
 sky130_fd_sc_hd__nand2b_1 _08865_ (.A_N(_02010_),
    .B(_02011_),
    .Y(_02018_));
 sky130_fd_sc_hd__nand2_1 _08866_ (.A(_02012_),
    .B(_02018_),
    .Y(_02019_));
 sky130_fd_sc_hd__a21o_1 _08867_ (.A1(_01416_),
    .A2(_01418_),
    .B1(_02019_),
    .X(_02020_));
 sky130_fd_sc_hd__xnor2_1 _08868_ (.A(_02017_),
    .B(_02019_),
    .Y(_02021_));
 sky130_fd_sc_hd__inv_2 _08869_ (.A(_02021_),
    .Y(_02022_));
 sky130_fd_sc_hd__nand2_1 _08870_ (.A(_02016_),
    .B(_02021_),
    .Y(_02023_));
 sky130_fd_sc_hd__a31oi_2 _08871_ (.A1(_01999_),
    .A2(_02000_),
    .A3(_02005_),
    .B1(_02023_),
    .Y(_02024_));
 sky130_fd_sc_hd__a21o_1 _08872_ (.A1(_02015_),
    .A2(_02020_),
    .B1(_02014_),
    .X(_02025_));
 sky130_fd_sc_hd__o32ai_1 _08873_ (.A1(_01128_),
    .A2(_01196_),
    .A3(_02025_),
    .B1(_01194_),
    .B2(_01127_),
    .Y(_02026_));
 sky130_fd_sc_hd__a211o_2 _08874_ (.A1(_01198_),
    .A2(_02024_),
    .B1(_02026_),
    .C1(_01126_),
    .X(_02027_));
 sky130_fd_sc_hd__a21bo_1 _08875_ (.A1(_01050_),
    .A2(_02027_),
    .B1_N(_01048_),
    .X(_02028_));
 sky130_fd_sc_hd__nor2_1 _08876_ (.A(_00976_),
    .B(_01048_),
    .Y(_02029_));
 sky130_fd_sc_hd__nor2_2 _08877_ (.A(_00975_),
    .B(_00976_),
    .Y(_02030_));
 sky130_fd_sc_hd__a311o_4 _08878_ (.A1(_01050_),
    .A2(_02027_),
    .A3(_02030_),
    .B1(_02029_),
    .C1(_00975_),
    .X(_02031_));
 sky130_fd_sc_hd__a21boi_2 _08879_ (.A1(_00897_),
    .A2(_02031_),
    .B1_N(_00895_),
    .Y(_02032_));
 sky130_fd_sc_hd__nor2_1 _08880_ (.A(_00813_),
    .B(_00895_),
    .Y(_02033_));
 sky130_fd_sc_hd__nor2_2 _08881_ (.A(_00812_),
    .B(_00813_),
    .Y(_02034_));
 sky130_fd_sc_hd__a311o_4 _08882_ (.A1(_00897_),
    .A2(_02031_),
    .A3(_02034_),
    .B1(_02033_),
    .C1(_00812_),
    .X(_02035_));
 sky130_fd_sc_hd__a21bo_2 _08883_ (.A1(_00799_),
    .A2(_00805_),
    .B1_N(_00807_),
    .X(_02036_));
 sky130_fd_sc_hd__o21ai_4 _08884_ (.A1(_00749_),
    .A2(_00776_),
    .B1(_00775_),
    .Y(_02037_));
 sky130_fd_sc_hd__o22a_1 _08885_ (.A1(net165),
    .A2(net12),
    .B1(net46),
    .B2(net149),
    .X(_02038_));
 sky130_fd_sc_hd__xnor2_1 _08886_ (.A(net97),
    .B(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__inv_2 _08887_ (.A(_02039_),
    .Y(_02040_));
 sky130_fd_sc_hd__o22a_1 _08888_ (.A1(net147),
    .A2(net13),
    .B1(net47),
    .B2(net144),
    .X(_02041_));
 sky130_fd_sc_hd__xnor2_1 _08889_ (.A(net109),
    .B(_02041_),
    .Y(_02042_));
 sky130_fd_sc_hd__xor2_1 _08890_ (.A(_02039_),
    .B(_02042_),
    .X(_02043_));
 sky130_fd_sc_hd__o22a_1 _08891_ (.A1(net15),
    .A2(net143),
    .B1(net141),
    .B2(net53),
    .X(_02044_));
 sky130_fd_sc_hd__xnor2_1 _08892_ (.A(net113),
    .B(_02044_),
    .Y(_02045_));
 sky130_fd_sc_hd__and2b_1 _08893_ (.A_N(_02043_),
    .B(_02045_),
    .X(_02046_));
 sky130_fd_sc_hd__and2b_1 _08894_ (.A_N(_02045_),
    .B(_02043_),
    .X(_02047_));
 sky130_fd_sc_hd__or2_1 _08895_ (.A(_02046_),
    .B(_02047_),
    .X(_02048_));
 sky130_fd_sc_hd__a21oi_1 _08896_ (.A1(_00721_),
    .A2(_00724_),
    .B1(_02048_),
    .Y(_02049_));
 sky130_fd_sc_hd__and3_1 _08897_ (.A(_00721_),
    .B(_00724_),
    .C(_02048_),
    .X(_02050_));
 sky130_fd_sc_hd__nor2_2 _08898_ (.A(_02049_),
    .B(_02050_),
    .Y(_02051_));
 sky130_fd_sc_hd__xor2_4 _08899_ (.A(_02037_),
    .B(_02051_),
    .X(_02052_));
 sky130_fd_sc_hd__a21o_1 _08900_ (.A1(_00741_),
    .A2(_00747_),
    .B1(_00746_),
    .X(_02053_));
 sky130_fd_sc_hd__xor2_1 _08901_ (.A(_00785_),
    .B(_02053_),
    .X(_02054_));
 sky130_fd_sc_hd__o21a_1 _08902_ (.A1(_00768_),
    .A2(_00772_),
    .B1(_02054_),
    .X(_02055_));
 sky130_fd_sc_hd__nor3_1 _08903_ (.A(_00768_),
    .B(_00772_),
    .C(_02054_),
    .Y(_02056_));
 sky130_fd_sc_hd__nor2_1 _08904_ (.A(_02055_),
    .B(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__o22a_1 _08905_ (.A1(net152),
    .A2(net65),
    .B1(net58),
    .B2(net150),
    .X(_02058_));
 sky130_fd_sc_hd__xnor2_1 _08906_ (.A(net191),
    .B(_02058_),
    .Y(_02059_));
 sky130_fd_sc_hd__o22a_1 _08907_ (.A1(net74),
    .A2(net116),
    .B1(net114),
    .B2(net68),
    .X(_02060_));
 sky130_fd_sc_hd__xnor2_1 _08908_ (.A(net179),
    .B(_02060_),
    .Y(_02061_));
 sky130_fd_sc_hd__o22a_1 _08909_ (.A1(net175),
    .A2(net63),
    .B1(net54),
    .B2(net177),
    .X(_02062_));
 sky130_fd_sc_hd__xnor2_1 _08910_ (.A(net189),
    .B(_02062_),
    .Y(_02063_));
 sky130_fd_sc_hd__nor2_1 _08911_ (.A(_02061_),
    .B(_02063_),
    .Y(_02064_));
 sky130_fd_sc_hd__and2_1 _08912_ (.A(_02061_),
    .B(_02063_),
    .X(_02065_));
 sky130_fd_sc_hd__nor2_1 _08913_ (.A(_02064_),
    .B(_02065_),
    .Y(_02066_));
 sky130_fd_sc_hd__xnor2_1 _08914_ (.A(_02059_),
    .B(_02066_),
    .Y(_02067_));
 sky130_fd_sc_hd__o22a_1 _08915_ (.A1(net130),
    .A2(net76),
    .B1(net71),
    .B2(net82),
    .X(_02068_));
 sky130_fd_sc_hd__xnor2_1 _08916_ (.A(net158),
    .B(_02068_),
    .Y(_02069_));
 sky130_fd_sc_hd__o22a_1 _08917_ (.A1(net80),
    .A2(net42),
    .B1(net94),
    .B2(net128),
    .X(_02070_));
 sky130_fd_sc_hd__xnor2_1 _08918_ (.A(net137),
    .B(_02070_),
    .Y(_02071_));
 sky130_fd_sc_hd__nand2b_1 _08919_ (.A_N(_02069_),
    .B(_02071_),
    .Y(_02072_));
 sky130_fd_sc_hd__xor2_1 _08920_ (.A(_02069_),
    .B(_02071_),
    .X(_02073_));
 sky130_fd_sc_hd__o22a_1 _08921_ (.A1(net123),
    .A2(net119),
    .B1(net100),
    .B2(net79),
    .X(_02074_));
 sky130_fd_sc_hd__xor2_1 _08922_ (.A(net154),
    .B(_02074_),
    .X(_02075_));
 sky130_fd_sc_hd__or2_1 _08923_ (.A(_02073_),
    .B(_02075_),
    .X(_02076_));
 sky130_fd_sc_hd__nand2_1 _08924_ (.A(_02073_),
    .B(_02075_),
    .Y(_02077_));
 sky130_fd_sc_hd__nand2_1 _08925_ (.A(_02076_),
    .B(_02077_),
    .Y(_02078_));
 sky130_fd_sc_hd__o22a_1 _08926_ (.A1(net173),
    .A2(net17),
    .B1(net9),
    .B2(net171),
    .X(_02079_));
 sky130_fd_sc_hd__xnor2_2 _08927_ (.A(_00180_),
    .B(_02079_),
    .Y(_02080_));
 sky130_fd_sc_hd__a32o_1 _08928_ (.A1(_00210_),
    .A2(_00219_),
    .A3(_00221_),
    .B1(_00208_),
    .B2(_00197_),
    .X(_02081_));
 sky130_fd_sc_hd__xnor2_2 _08929_ (.A(net210),
    .B(_02081_),
    .Y(_02082_));
 sky130_fd_sc_hd__a21oi_2 _08930_ (.A1(net302),
    .A2(_00756_),
    .B1(_00188_),
    .Y(_02083_));
 sky130_fd_sc_hd__and2_1 _08931_ (.A(_02082_),
    .B(_02083_),
    .X(_02084_));
 sky130_fd_sc_hd__xor2_2 _08932_ (.A(_02082_),
    .B(_02083_),
    .X(_02085_));
 sky130_fd_sc_hd__xor2_2 _08933_ (.A(_02080_),
    .B(_02085_),
    .X(_02086_));
 sky130_fd_sc_hd__xnor2_1 _08934_ (.A(_02078_),
    .B(_02086_),
    .Y(_02087_));
 sky130_fd_sc_hd__xnor2_1 _08935_ (.A(_02067_),
    .B(_02087_),
    .Y(_02088_));
 sky130_fd_sc_hd__nor2_1 _08936_ (.A(_06309_),
    .B(net32),
    .Y(_02089_));
 sky130_fd_sc_hd__a21o_1 _08937_ (.A1(_00752_),
    .A2(_00761_),
    .B1(_00760_),
    .X(_02090_));
 sky130_fd_sc_hd__o22a_1 _08938_ (.A1(net8),
    .A2(net161),
    .B1(net6),
    .B2(net163),
    .X(_02091_));
 sky130_fd_sc_hd__xnor2_1 _08939_ (.A(net33),
    .B(_02091_),
    .Y(_02092_));
 sky130_fd_sc_hd__nand2_1 _08940_ (.A(_02090_),
    .B(_02092_),
    .Y(_02093_));
 sky130_fd_sc_hd__xor2_1 _08941_ (.A(_02090_),
    .B(_02092_),
    .X(_02094_));
 sky130_fd_sc_hd__xnor2_1 _08942_ (.A(_02089_),
    .B(_02094_),
    .Y(_02095_));
 sky130_fd_sc_hd__nor2_1 _08943_ (.A(_02088_),
    .B(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__xor2_1 _08944_ (.A(_02088_),
    .B(_02095_),
    .X(_02097_));
 sky130_fd_sc_hd__xnor2_1 _08945_ (.A(_02057_),
    .B(_02097_),
    .Y(_02098_));
 sky130_fd_sc_hd__o21bai_2 _08946_ (.A1(_00712_),
    .A2(_00715_),
    .B1_N(_00711_),
    .Y(_02099_));
 sky130_fd_sc_hd__o22a_1 _08947_ (.A1(net51),
    .A2(net132),
    .B1(net89),
    .B2(net49),
    .X(_02100_));
 sky130_fd_sc_hd__xnor2_1 _08948_ (.A(net106),
    .B(_02100_),
    .Y(_02101_));
 sky130_fd_sc_hd__o22a_1 _08949_ (.A1(net125),
    .A2(net36),
    .B1(net34),
    .B2(net121),
    .X(_02102_));
 sky130_fd_sc_hd__xnor2_1 _08950_ (.A(net135),
    .B(_02102_),
    .Y(_02103_));
 sky130_fd_sc_hd__and2_1 _08951_ (.A(_02101_),
    .B(_02103_),
    .X(_02104_));
 sky130_fd_sc_hd__nor2_1 _08952_ (.A(_02101_),
    .B(_02103_),
    .Y(_02105_));
 sky130_fd_sc_hd__nor2_1 _08953_ (.A(_02104_),
    .B(_02105_),
    .Y(_02106_));
 sky130_fd_sc_hd__o22a_1 _08954_ (.A1(net92),
    .A2(net38),
    .B1(net87),
    .B2(net41),
    .X(_02107_));
 sky130_fd_sc_hd__xnor2_1 _08955_ (.A(net102),
    .B(_02107_),
    .Y(_02108_));
 sky130_fd_sc_hd__xor2_1 _08956_ (.A(_02106_),
    .B(_02108_),
    .X(_02109_));
 sky130_fd_sc_hd__o21a_1 _08957_ (.A1(_00732_),
    .A2(_00737_),
    .B1(_00736_),
    .X(_02110_));
 sky130_fd_sc_hd__and2b_1 _08958_ (.A_N(_02110_),
    .B(_02109_),
    .X(_02111_));
 sky130_fd_sc_hd__xnor2_1 _08959_ (.A(_02109_),
    .B(_02110_),
    .Y(_02112_));
 sky130_fd_sc_hd__xnor2_1 _08960_ (.A(_02099_),
    .B(_02112_),
    .Y(_02113_));
 sky130_fd_sc_hd__nor2_1 _08961_ (.A(_02098_),
    .B(_02113_),
    .Y(_02114_));
 sky130_fd_sc_hd__nand2_1 _08962_ (.A(_02098_),
    .B(_02113_),
    .Y(_02115_));
 sky130_fd_sc_hd__and2b_1 _08963_ (.A_N(_02114_),
    .B(_02115_),
    .X(_02116_));
 sky130_fd_sc_hd__xor2_4 _08964_ (.A(_02052_),
    .B(_02116_),
    .X(_02117_));
 sky130_fd_sc_hd__o31ai_2 _08965_ (.A1(_00780_),
    .A2(_00791_),
    .A3(_00792_),
    .B1(_00795_),
    .Y(_02118_));
 sky130_fd_sc_hd__o21ai_4 _08966_ (.A1(_00706_),
    .A2(_00719_),
    .B1(_00717_),
    .Y(_02119_));
 sky130_fd_sc_hd__o21a_2 _08967_ (.A1(_00726_),
    .A2(_00779_),
    .B1(_00778_),
    .X(_02120_));
 sky130_fd_sc_hd__a21oi_2 _08968_ (.A1(_00787_),
    .A2(_00789_),
    .B1(_00791_),
    .Y(_02121_));
 sky130_fd_sc_hd__nor2_1 _08969_ (.A(_02120_),
    .B(_02121_),
    .Y(_02122_));
 sky130_fd_sc_hd__xor2_4 _08970_ (.A(_02120_),
    .B(_02121_),
    .X(_02123_));
 sky130_fd_sc_hd__xnor2_2 _08971_ (.A(_02119_),
    .B(_02123_),
    .Y(_02124_));
 sky130_fd_sc_hd__a21oi_2 _08972_ (.A1(_00800_),
    .A2(_00804_),
    .B1(_00803_),
    .Y(_02125_));
 sky130_fd_sc_hd__xnor2_1 _08973_ (.A(_02124_),
    .B(_02125_),
    .Y(_02126_));
 sky130_fd_sc_hd__nand2b_1 _08974_ (.A_N(_02126_),
    .B(_02118_),
    .Y(_02127_));
 sky130_fd_sc_hd__xnor2_2 _08975_ (.A(_02118_),
    .B(_02126_),
    .Y(_02128_));
 sky130_fd_sc_hd__and2_1 _08976_ (.A(_02117_),
    .B(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__xor2_4 _08977_ (.A(_02117_),
    .B(_02128_),
    .X(_02130_));
 sky130_fd_sc_hd__xnor2_4 _08978_ (.A(_02036_),
    .B(_02130_),
    .Y(_02131_));
 sky130_fd_sc_hd__a21oi_4 _08979_ (.A1(_00705_),
    .A2(_00810_),
    .B1(_00809_),
    .Y(_02132_));
 sky130_fd_sc_hd__nor2_1 _08980_ (.A(_02131_),
    .B(_02132_),
    .Y(_02133_));
 sky130_fd_sc_hd__xor2_4 _08981_ (.A(_02131_),
    .B(_02132_),
    .X(_02134_));
 sky130_fd_sc_hd__xor2_4 _08982_ (.A(_02035_),
    .B(_02134_),
    .X(_02135_));
 sky130_fd_sc_hd__nor2_1 _08983_ (.A(net299),
    .B(_04796_),
    .Y(_02136_));
 sky130_fd_sc_hd__nand2_2 _08984_ (.A(net306),
    .B(_04785_),
    .Y(_02137_));
 sky130_fd_sc_hd__xor2_4 _08985_ (.A(_00897_),
    .B(_02031_),
    .X(_02138_));
 sky130_fd_sc_hd__xnor2_2 _08986_ (.A(_01049_),
    .B(_02027_),
    .Y(_02139_));
 sky130_fd_sc_hd__nand2b_1 _08987_ (.A_N(_02024_),
    .B(_02025_),
    .Y(_02140_));
 sky130_fd_sc_hd__xnor2_2 _08988_ (.A(_01196_),
    .B(_02140_),
    .Y(_02141_));
 sky130_fd_sc_hd__a31o_1 _08989_ (.A1(_01999_),
    .A2(_02000_),
    .A3(_02005_),
    .B1(_02022_),
    .X(_02142_));
 sky130_fd_sc_hd__a21bo_1 _08990_ (.A1(_02020_),
    .A2(_02142_),
    .B1_N(_02016_),
    .X(_02143_));
 sky130_fd_sc_hd__nand3b_1 _08991_ (.A_N(_02016_),
    .B(_02020_),
    .C(_02142_),
    .Y(_02144_));
 sky130_fd_sc_hd__and2_1 _08992_ (.A(_02143_),
    .B(_02144_),
    .X(_02145_));
 sky130_fd_sc_hd__a31o_1 _08993_ (.A1(_01520_),
    .A2(_01523_),
    .A3(_01998_),
    .B1(_02002_),
    .X(_02146_));
 sky130_fd_sc_hd__a21oi_1 _08994_ (.A1(_01405_),
    .A2(_02146_),
    .B1(_01404_),
    .Y(_02147_));
 sky130_fd_sc_hd__xnor2_1 _08995_ (.A(_01420_),
    .B(_02147_),
    .Y(_02148_));
 sky130_fd_sc_hd__xor2_2 _08996_ (.A(_01405_),
    .B(_02146_),
    .X(_02149_));
 sky130_fd_sc_hd__a21oi_1 _08997_ (.A1(_01520_),
    .A2(_01998_),
    .B1(_01518_),
    .Y(_02150_));
 sky130_fd_sc_hd__xnor2_1 _08998_ (.A(_01523_),
    .B(_02150_),
    .Y(_02151_));
 sky130_fd_sc_hd__a31o_1 _08999_ (.A1(_01993_),
    .A2(_01995_),
    .A3(_01996_),
    .B1(_01708_),
    .X(_02152_));
 sky130_fd_sc_hd__xor2_2 _09000_ (.A(_01624_),
    .B(_02152_),
    .X(_02153_));
 sky130_fd_sc_hd__xnor2_1 _09001_ (.A(_01993_),
    .B(_01995_),
    .Y(_02154_));
 sky130_fd_sc_hd__xnor2_2 _09002_ (.A(_01804_),
    .B(_01990_),
    .Y(_02155_));
 sky130_fd_sc_hd__xnor2_2 _09003_ (.A(_01833_),
    .B(_01989_),
    .Y(_02156_));
 sky130_fd_sc_hd__xor2_1 _09004_ (.A(_01880_),
    .B(_01986_),
    .X(_02157_));
 sky130_fd_sc_hd__xnor2_1 _09005_ (.A(_01901_),
    .B(_01985_),
    .Y(_02158_));
 sky130_fd_sc_hd__xor2_1 _09006_ (.A(_01915_),
    .B(_01984_),
    .X(_02159_));
 sky130_fd_sc_hd__xnor2_1 _09007_ (.A(_01932_),
    .B(_01983_),
    .Y(_02160_));
 sky130_fd_sc_hd__xnor2_1 _09008_ (.A(_01948_),
    .B(_01982_),
    .Y(_02161_));
 sky130_fd_sc_hd__xor2_1 _09009_ (.A(_01957_),
    .B(_01981_),
    .X(_02162_));
 sky130_fd_sc_hd__or3_1 _09010_ (.A(_01964_),
    .B(_01971_),
    .C(_01979_),
    .X(_02163_));
 sky130_fd_sc_hd__and2_1 _09011_ (.A(_01980_),
    .B(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__and2_1 _09012_ (.A(_01972_),
    .B(_01978_),
    .X(_02165_));
 sky130_fd_sc_hd__or2_1 _09013_ (.A(_01979_),
    .B(_02165_),
    .X(_02166_));
 sky130_fd_sc_hd__xor2_1 _09014_ (.A(_01974_),
    .B(_01977_),
    .X(_02167_));
 sky130_fd_sc_hd__nor2_1 _09015_ (.A(_01976_),
    .B(_02167_),
    .Y(_02168_));
 sky130_fd_sc_hd__nand2_1 _09016_ (.A(_02166_),
    .B(_02168_),
    .Y(_02169_));
 sky130_fd_sc_hd__or2_1 _09017_ (.A(_02164_),
    .B(_02169_),
    .X(_02170_));
 sky130_fd_sc_hd__nor2_1 _09018_ (.A(_02162_),
    .B(_02170_),
    .Y(_02171_));
 sky130_fd_sc_hd__nand2_1 _09019_ (.A(_02161_),
    .B(_02171_),
    .Y(_02172_));
 sky130_fd_sc_hd__or2_1 _09020_ (.A(_02160_),
    .B(_02172_),
    .X(_02173_));
 sky130_fd_sc_hd__nor2_1 _09021_ (.A(_02159_),
    .B(_02173_),
    .Y(_02174_));
 sky130_fd_sc_hd__nand2_1 _09022_ (.A(_02158_),
    .B(_02174_),
    .Y(_02175_));
 sky130_fd_sc_hd__or2_1 _09023_ (.A(_02157_),
    .B(_02175_),
    .X(_02176_));
 sky130_fd_sc_hd__a21oi_1 _09024_ (.A1(_01880_),
    .A2(_01986_),
    .B1(_01876_),
    .Y(_02177_));
 sky130_fd_sc_hd__xnor2_2 _09025_ (.A(_01988_),
    .B(_02177_),
    .Y(_02178_));
 sky130_fd_sc_hd__nor2_1 _09026_ (.A(_02176_),
    .B(_02178_),
    .Y(_02179_));
 sky130_fd_sc_hd__nor3b_1 _09027_ (.A(_02176_),
    .B(_02178_),
    .C_N(_02156_),
    .Y(_02180_));
 sky130_fd_sc_hd__nand2_1 _09028_ (.A(_02155_),
    .B(_02180_),
    .Y(_02181_));
 sky130_fd_sc_hd__nand2b_1 _09029_ (.A_N(_01774_),
    .B(_01775_),
    .Y(_02182_));
 sky130_fd_sc_hd__xnor2_2 _09030_ (.A(_01991_),
    .B(_02182_),
    .Y(_02183_));
 sky130_fd_sc_hd__nor2_1 _09031_ (.A(_02181_),
    .B(_02183_),
    .Y(_02184_));
 sky130_fd_sc_hd__and2b_1 _09032_ (.A_N(_01740_),
    .B(_01741_),
    .X(_02185_));
 sky130_fd_sc_hd__xnor2_1 _09033_ (.A(_01992_),
    .B(_02185_),
    .Y(_02186_));
 sky130_fd_sc_hd__and2_1 _09034_ (.A(_02184_),
    .B(_02186_),
    .X(_02187_));
 sky130_fd_sc_hd__nand2_1 _09035_ (.A(_02154_),
    .B(_02187_),
    .Y(_02188_));
 sky130_fd_sc_hd__a21oi_1 _09036_ (.A1(_01993_),
    .A2(_01995_),
    .B1(_01705_),
    .Y(_02189_));
 sky130_fd_sc_hd__xnor2_2 _09037_ (.A(_01996_),
    .B(_02189_),
    .Y(_02190_));
 sky130_fd_sc_hd__or2_1 _09038_ (.A(_02188_),
    .B(_02190_),
    .X(_02191_));
 sky130_fd_sc_hd__or3_1 _09039_ (.A(_02153_),
    .B(_02188_),
    .C(_02190_),
    .X(_02192_));
 sky130_fd_sc_hd__a21o_1 _09040_ (.A1(_01624_),
    .A2(_02152_),
    .B1(_01623_),
    .X(_02193_));
 sky130_fd_sc_hd__xnor2_2 _09041_ (.A(_01575_),
    .B(_02193_),
    .Y(_02194_));
 sky130_fd_sc_hd__or2_1 _09042_ (.A(_02192_),
    .B(_02194_),
    .X(_02195_));
 sky130_fd_sc_hd__xor2_2 _09043_ (.A(_01520_),
    .B(_01998_),
    .X(_02196_));
 sky130_fd_sc_hd__or2_1 _09044_ (.A(_02195_),
    .B(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__or4_2 _09045_ (.A(_02151_),
    .B(_02192_),
    .C(_02194_),
    .D(_02196_),
    .X(_02198_));
 sky130_fd_sc_hd__or2_1 _09046_ (.A(_02149_),
    .B(_02198_),
    .X(_02199_));
 sky130_fd_sc_hd__or2_1 _09047_ (.A(_02148_),
    .B(_02199_),
    .X(_02200_));
 sky130_fd_sc_hd__nand4_1 _09048_ (.A(_01999_),
    .B(_02000_),
    .C(_02005_),
    .D(_02022_),
    .Y(_02201_));
 sky130_fd_sc_hd__and2_1 _09049_ (.A(_02142_),
    .B(_02201_),
    .X(_02202_));
 sky130_fd_sc_hd__or2_1 _09050_ (.A(_02200_),
    .B(_02202_),
    .X(_02203_));
 sky130_fd_sc_hd__a21o_1 _09051_ (.A1(_02143_),
    .A2(_02144_),
    .B1(_02202_),
    .X(_02204_));
 sky130_fd_sc_hd__or4_2 _09052_ (.A(_02148_),
    .B(_02149_),
    .C(_02198_),
    .D(_02204_),
    .X(_02205_));
 sky130_fd_sc_hd__nor2_1 _09053_ (.A(_02141_),
    .B(_02205_),
    .Y(_02206_));
 sky130_fd_sc_hd__a21oi_1 _09054_ (.A1(_01197_),
    .A2(_02140_),
    .B1(_01193_),
    .Y(_02207_));
 sky130_fd_sc_hd__xnor2_2 _09055_ (.A(_01128_),
    .B(_02207_),
    .Y(_02208_));
 sky130_fd_sc_hd__or4b_2 _09056_ (.A(_02139_),
    .B(_02141_),
    .C(_02205_),
    .D_N(_02208_),
    .X(_02209_));
 sky130_fd_sc_hd__xor2_4 _09057_ (.A(_02028_),
    .B(_02030_),
    .X(_02210_));
 sky130_fd_sc_hd__xnor2_4 _09058_ (.A(_02032_),
    .B(_02034_),
    .Y(_02211_));
 sky130_fd_sc_hd__or4_4 _09059_ (.A(_02138_),
    .B(_02209_),
    .C(_02210_),
    .D(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__nor2_2 _09060_ (.A(_06388_),
    .B(_06395_),
    .Y(_02213_));
 sky130_fd_sc_hd__or2_4 _09061_ (.A(_06388_),
    .B(_06395_),
    .X(_02214_));
 sky130_fd_sc_hd__a21oi_1 _09062_ (.A1(net22),
    .A2(_02212_),
    .B1(_02135_),
    .Y(_02215_));
 sky130_fd_sc_hd__a31o_1 _09063_ (.A1(_02135_),
    .A2(net22),
    .A3(_02212_),
    .B1(_02214_),
    .X(_02216_));
 sky130_fd_sc_hd__nor2_2 _09064_ (.A(net299),
    .B(_06417_),
    .Y(_02217_));
 sky130_fd_sc_hd__nand2_1 _09065_ (.A(net305),
    .B(_06416_),
    .Y(_02218_));
 sky130_fd_sc_hd__mux2_1 _09066_ (.A0(net304),
    .A1(reg1_val[31]),
    .S(net187),
    .X(_02219_));
 sky130_fd_sc_hd__mux2_1 _09067_ (.A0(reg1_val[1]),
    .A1(reg1_val[30]),
    .S(net187),
    .X(_02220_));
 sky130_fd_sc_hd__mux2_1 _09068_ (.A0(_02219_),
    .A1(_02220_),
    .S(net227),
    .X(_02221_));
 sky130_fd_sc_hd__mux2_1 _09069_ (.A0(reg1_val[3]),
    .A1(reg1_val[28]),
    .S(net187),
    .X(_02222_));
 sky130_fd_sc_hd__mux2_1 _09070_ (.A0(reg1_val[2]),
    .A1(reg1_val[29]),
    .S(net187),
    .X(_02223_));
 sky130_fd_sc_hd__mux2_1 _09071_ (.A0(_02222_),
    .A1(_02223_),
    .S(net224),
    .X(_02224_));
 sky130_fd_sc_hd__mux2_1 _09072_ (.A0(_02221_),
    .A1(_02224_),
    .S(net230),
    .X(_02225_));
 sky130_fd_sc_hd__mux2_1 _09073_ (.A0(reg1_val[7]),
    .A1(reg1_val[24]),
    .S(net187),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _09074_ (.A0(reg1_val[6]),
    .A1(reg1_val[25]),
    .S(net187),
    .X(_02227_));
 sky130_fd_sc_hd__mux2_1 _09075_ (.A0(_02226_),
    .A1(_02227_),
    .S(net224),
    .X(_02228_));
 sky130_fd_sc_hd__mux2_1 _09076_ (.A0(reg1_val[5]),
    .A1(reg1_val[26]),
    .S(net187),
    .X(_02229_));
 sky130_fd_sc_hd__mux2_1 _09077_ (.A0(reg1_val[4]),
    .A1(reg1_val[27]),
    .S(net187),
    .X(_02230_));
 sky130_fd_sc_hd__mux2_1 _09078_ (.A0(_02229_),
    .A1(_02230_),
    .S(net224),
    .X(_02231_));
 sky130_fd_sc_hd__mux2_1 _09079_ (.A0(_02228_),
    .A1(_02231_),
    .S(net228),
    .X(_02232_));
 sky130_fd_sc_hd__mux2_1 _09080_ (.A0(_02225_),
    .A1(_02232_),
    .S(net232),
    .X(_02233_));
 sky130_fd_sc_hd__mux2_1 _09081_ (.A0(reg1_val[15]),
    .A1(reg1_val[16]),
    .S(net187),
    .X(_02234_));
 sky130_fd_sc_hd__mux2_1 _09082_ (.A0(reg1_val[14]),
    .A1(reg1_val[17]),
    .S(net187),
    .X(_02235_));
 sky130_fd_sc_hd__mux2_1 _09083_ (.A0(_02234_),
    .A1(_02235_),
    .S(net225),
    .X(_02236_));
 sky130_fd_sc_hd__mux2_1 _09084_ (.A0(net303),
    .A1(reg1_val[18]),
    .S(net187),
    .X(_02237_));
 sky130_fd_sc_hd__mux2_1 _09085_ (.A0(reg1_val[12]),
    .A1(reg1_val[19]),
    .S(net187),
    .X(_02238_));
 sky130_fd_sc_hd__mux2_1 _09086_ (.A0(_02237_),
    .A1(_02238_),
    .S(net225),
    .X(_02239_));
 sky130_fd_sc_hd__mux2_1 _09087_ (.A0(_02236_),
    .A1(_02239_),
    .S(net229),
    .X(_02240_));
 sky130_fd_sc_hd__mux2_1 _09088_ (.A0(reg1_val[11]),
    .A1(reg1_val[20]),
    .S(net187),
    .X(_02241_));
 sky130_fd_sc_hd__mux2_1 _09089_ (.A0(reg1_val[10]),
    .A1(reg1_val[21]),
    .S(net187),
    .X(_02242_));
 sky130_fd_sc_hd__mux2_1 _09090_ (.A0(_02241_),
    .A1(_02242_),
    .S(net224),
    .X(_02243_));
 sky130_fd_sc_hd__mux2_1 _09091_ (.A0(reg1_val[9]),
    .A1(reg1_val[22]),
    .S(net187),
    .X(_02244_));
 sky130_fd_sc_hd__mux2_1 _09092_ (.A0(reg1_val[8]),
    .A1(reg1_val[23]),
    .S(net187),
    .X(_02245_));
 sky130_fd_sc_hd__mux2_1 _09093_ (.A0(_02244_),
    .A1(_02245_),
    .S(net224),
    .X(_02246_));
 sky130_fd_sc_hd__mux2_1 _09094_ (.A0(_02243_),
    .A1(_02246_),
    .S(net229),
    .X(_02247_));
 sky130_fd_sc_hd__mux2_1 _09095_ (.A0(_02247_),
    .A1(_02240_),
    .S(net232),
    .X(_02248_));
 sky130_fd_sc_hd__mux2_1 _09096_ (.A0(_02233_),
    .A1(_02248_),
    .S(net234),
    .X(_02249_));
 sky130_fd_sc_hd__mux2_1 _09097_ (.A0(reg1_val[8]),
    .A1(reg1_val[23]),
    .S(net184),
    .X(_02250_));
 sky130_fd_sc_hd__mux2_1 _09098_ (.A0(reg1_val[9]),
    .A1(reg1_val[22]),
    .S(net184),
    .X(_02251_));
 sky130_fd_sc_hd__mux2_1 _09099_ (.A0(_02250_),
    .A1(_02251_),
    .S(net225),
    .X(_02252_));
 sky130_fd_sc_hd__mux2_1 _09100_ (.A0(reg1_val[10]),
    .A1(reg1_val[21]),
    .S(net184),
    .X(_02253_));
 sky130_fd_sc_hd__mux2_1 _09101_ (.A0(reg1_val[11]),
    .A1(reg1_val[20]),
    .S(net184),
    .X(_02254_));
 sky130_fd_sc_hd__mux2_1 _09102_ (.A0(_02253_),
    .A1(_02254_),
    .S(net224),
    .X(_02255_));
 sky130_fd_sc_hd__mux2_1 _09103_ (.A0(_02252_),
    .A1(_02255_),
    .S(net228),
    .X(_02256_));
 sky130_fd_sc_hd__mux2_1 _09104_ (.A0(reg1_val[12]),
    .A1(reg1_val[19]),
    .S(net184),
    .X(_02257_));
 sky130_fd_sc_hd__mux2_1 _09105_ (.A0(net303),
    .A1(reg1_val[18]),
    .S(net184),
    .X(_02258_));
 sky130_fd_sc_hd__mux2_1 _09106_ (.A0(_02257_),
    .A1(_02258_),
    .S(net225),
    .X(_02259_));
 sky130_fd_sc_hd__mux2_1 _09107_ (.A0(reg1_val[14]),
    .A1(reg1_val[17]),
    .S(net184),
    .X(_02260_));
 sky130_fd_sc_hd__mux2_1 _09108_ (.A0(reg1_val[15]),
    .A1(reg1_val[16]),
    .S(net184),
    .X(_02261_));
 sky130_fd_sc_hd__mux2_1 _09109_ (.A0(_02260_),
    .A1(_02261_),
    .S(net225),
    .X(_02262_));
 sky130_fd_sc_hd__mux2_1 _09110_ (.A0(_02259_),
    .A1(_02262_),
    .S(net228),
    .X(_02263_));
 sky130_fd_sc_hd__mux2_1 _09111_ (.A0(_02263_),
    .A1(_02256_),
    .S(net232),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _09112_ (.A0(net304),
    .A1(reg1_val[31]),
    .S(net185),
    .X(_02265_));
 sky130_fd_sc_hd__inv_2 _09113_ (.A(_02265_),
    .Y(_02266_));
 sky130_fd_sc_hd__mux2_1 _09114_ (.A0(reg1_val[1]),
    .A1(reg1_val[30]),
    .S(net184),
    .X(_02267_));
 sky130_fd_sc_hd__mux2_1 _09115_ (.A0(_02265_),
    .A1(_02267_),
    .S(net224),
    .X(_02268_));
 sky130_fd_sc_hd__mux2_1 _09116_ (.A0(reg1_val[2]),
    .A1(reg1_val[29]),
    .S(net184),
    .X(_02269_));
 sky130_fd_sc_hd__mux2_1 _09117_ (.A0(reg1_val[3]),
    .A1(reg1_val[28]),
    .S(net184),
    .X(_02270_));
 sky130_fd_sc_hd__mux2_1 _09118_ (.A0(_02269_),
    .A1(_02270_),
    .S(net224),
    .X(_02271_));
 sky130_fd_sc_hd__mux2_1 _09119_ (.A0(_02268_),
    .A1(_02271_),
    .S(net228),
    .X(_02272_));
 sky130_fd_sc_hd__mux2_1 _09120_ (.A0(reg1_val[4]),
    .A1(reg1_val[27]),
    .S(net184),
    .X(_02273_));
 sky130_fd_sc_hd__mux2_1 _09121_ (.A0(reg1_val[5]),
    .A1(reg1_val[26]),
    .S(net185),
    .X(_02274_));
 sky130_fd_sc_hd__mux2_1 _09122_ (.A0(_02273_),
    .A1(_02274_),
    .S(net224),
    .X(_02275_));
 sky130_fd_sc_hd__mux2_1 _09123_ (.A0(reg1_val[6]),
    .A1(reg1_val[25]),
    .S(net185),
    .X(_02276_));
 sky130_fd_sc_hd__mux2_1 _09124_ (.A0(reg1_val[7]),
    .A1(reg1_val[24]),
    .S(net185),
    .X(_02277_));
 sky130_fd_sc_hd__mux2_1 _09125_ (.A0(_02276_),
    .A1(_02277_),
    .S(net224),
    .X(_02278_));
 sky130_fd_sc_hd__mux2_1 _09126_ (.A0(_02275_),
    .A1(_02278_),
    .S(net229),
    .X(_02279_));
 sky130_fd_sc_hd__mux2_1 _09127_ (.A0(_02279_),
    .A1(_02272_),
    .S(net232),
    .X(_02280_));
 sky130_fd_sc_hd__mux2_1 _09128_ (.A0(_02264_),
    .A1(_02280_),
    .S(net234),
    .X(_02281_));
 sky130_fd_sc_hd__or2_1 _09129_ (.A(net239),
    .B(_02249_),
    .X(_02282_));
 sky130_fd_sc_hd__o21ai_2 _09130_ (.A1(net237),
    .A2(_02281_),
    .B1(_02282_),
    .Y(_02283_));
 sky130_fd_sc_hd__nand2_1 _09131_ (.A(net304),
    .B(curr_PC[0]),
    .Y(_02284_));
 sky130_fd_sc_hd__or2_1 _09132_ (.A(net304),
    .B(curr_PC[0]),
    .X(_02285_));
 sky130_fd_sc_hd__a21oi_1 _09133_ (.A1(_02284_),
    .A2(_02285_),
    .B1(net241),
    .Y(_02286_));
 sky130_fd_sc_hd__a211o_1 _09134_ (.A1(net241),
    .A2(_02283_),
    .B1(_02286_),
    .C1(net214),
    .X(_02287_));
 sky130_fd_sc_hd__nor2_2 _09135_ (.A(net305),
    .B(_06417_),
    .Y(_02288_));
 sky130_fd_sc_hd__nand2_1 _09136_ (.A(net299),
    .B(_06416_),
    .Y(_02289_));
 sky130_fd_sc_hd__nor2_2 _09137_ (.A(_06415_),
    .B(_06423_),
    .Y(_02290_));
 sky130_fd_sc_hd__or2_4 _09138_ (.A(_06415_),
    .B(_06423_),
    .X(_02291_));
 sky130_fd_sc_hd__nor2_1 _09139_ (.A(_06370_),
    .B(_06414_),
    .Y(_02292_));
 sky130_fd_sc_hd__or2_4 _09140_ (.A(_06370_),
    .B(_06414_),
    .X(_02293_));
 sky130_fd_sc_hd__nor2_8 _09141_ (.A(_06386_),
    .B(_06423_),
    .Y(_02294_));
 sky130_fd_sc_hd__or2_4 _09142_ (.A(_06386_),
    .B(_06423_),
    .X(_02295_));
 sky130_fd_sc_hd__o21a_1 _09143_ (.A1(net251),
    .A2(_02294_),
    .B1(_06371_),
    .X(_02296_));
 sky130_fd_sc_hd__o21a_1 _09144_ (.A1(net205),
    .A2(_02296_),
    .B1(_06372_),
    .X(_02297_));
 sky130_fd_sc_hd__nor2_8 _09145_ (.A(_06370_),
    .B(_06395_),
    .Y(_02298_));
 sky130_fd_sc_hd__or2_2 _09146_ (.A(_06370_),
    .B(_06395_),
    .X(_02299_));
 sky130_fd_sc_hd__and4bb_4 _09147_ (.A_N(instruction[4]),
    .B_N(instruction[6]),
    .C(instruction[5]),
    .D(instruction[3]),
    .X(_02300_));
 sky130_fd_sc_hd__or3b_4 _09148_ (.A(_06388_),
    .B(instruction[6]),
    .C_N(instruction[5]),
    .X(_02301_));
 sky130_fd_sc_hd__a21oi_1 _09149_ (.A1(net250),
    .A2(_02301_),
    .B1(_06371_),
    .Y(_02302_));
 sky130_fd_sc_hd__nor2_2 _09150_ (.A(_06386_),
    .B(_06395_),
    .Y(_02303_));
 sky130_fd_sc_hd__or2_1 _09151_ (.A(_06386_),
    .B(_06395_),
    .X(_02304_));
 sky130_fd_sc_hd__nor2_2 _09152_ (.A(_06395_),
    .B(_06415_),
    .Y(_02305_));
 sky130_fd_sc_hd__or2_1 _09153_ (.A(_06395_),
    .B(_06415_),
    .X(_02306_));
 sky130_fd_sc_hd__a221o_1 _09154_ (.A1(\div_shifter[32] ),
    .A2(_02303_),
    .B1(_02305_),
    .B2(\div_res[0] ),
    .C1(_02302_),
    .X(_02307_));
 sky130_fd_sc_hd__nor2_1 _09155_ (.A(_02297_),
    .B(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__nand2_4 _09156_ (.A(reg1_val[31]),
    .B(net215),
    .Y(_02309_));
 sky130_fd_sc_hd__inv_2 _09157_ (.A(_02309_),
    .Y(_02310_));
 sky130_fd_sc_hd__nor2_1 _09158_ (.A(net237),
    .B(_02310_),
    .Y(_02311_));
 sky130_fd_sc_hd__nand2_8 _09159_ (.A(net238),
    .B(_02309_),
    .Y(_02312_));
 sky130_fd_sc_hd__mux2_1 _09160_ (.A0(_02266_),
    .A1(_02309_),
    .S(net227),
    .X(_02313_));
 sky130_fd_sc_hd__inv_2 _09161_ (.A(_02313_),
    .Y(_02314_));
 sky130_fd_sc_hd__a21o_1 _09162_ (.A1(net230),
    .A2(_02309_),
    .B1(_02313_),
    .X(_02315_));
 sky130_fd_sc_hd__nand2_1 _09163_ (.A(net232),
    .B(_02309_),
    .Y(_02316_));
 sky130_fd_sc_hd__and2b_1 _09164_ (.A_N(_02315_),
    .B(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__nand2_2 _09165_ (.A(net234),
    .B(_02309_),
    .Y(_02318_));
 sky130_fd_sc_hd__nand2_1 _09166_ (.A(_02317_),
    .B(_02318_),
    .Y(_02319_));
 sky130_fd_sc_hd__inv_2 _09167_ (.A(_02319_),
    .Y(_02320_));
 sky130_fd_sc_hd__or2_2 _09168_ (.A(_02311_),
    .B(_02319_),
    .X(_02321_));
 sky130_fd_sc_hd__o221a_1 _09169_ (.A1(_02283_),
    .A2(net182),
    .B1(_02321_),
    .B2(net186),
    .C1(_02308_),
    .X(_02322_));
 sky130_fd_sc_hd__o311a_1 _09170_ (.A1(instruction[5]),
    .A2(_06357_),
    .A3(_06386_),
    .B1(_02287_),
    .C1(_02322_),
    .X(_02323_));
 sky130_fd_sc_hd__o21a_1 _09171_ (.A1(_02215_),
    .A2(_02216_),
    .B1(_02323_),
    .X(_02324_));
 sky130_fd_sc_hd__a21bo_1 _09172_ (.A1(_06368_),
    .A2(_06424_),
    .B1_N(_02324_),
    .X(_02325_));
 sky130_fd_sc_hd__a22o_1 _09173_ (.A1(net227),
    .A2(net212),
    .B1(_06427_),
    .B2(_02325_),
    .X(_02326_));
 sky130_fd_sc_hd__mux2_8 _09174_ (.A0(_04514_),
    .A1(_02326_),
    .S(net258),
    .X(dest_val[0]));
 sky130_fd_sc_hd__a21oi_4 _09175_ (.A1(_02036_),
    .A2(_02130_),
    .B1(_02129_),
    .Y(_02327_));
 sky130_fd_sc_hd__o21ai_4 _09176_ (.A1(_02124_),
    .A2(_02125_),
    .B1(_02127_),
    .Y(_02328_));
 sky130_fd_sc_hd__a32o_2 _09177_ (.A1(_02076_),
    .A2(_02077_),
    .A3(_02086_),
    .B1(_02087_),
    .B2(_02067_),
    .X(_02329_));
 sky130_fd_sc_hd__o22a_1 _09178_ (.A1(net149),
    .A2(net12),
    .B1(net45),
    .B2(net143),
    .X(_02330_));
 sky130_fd_sc_hd__xnor2_1 _09179_ (.A(net97),
    .B(_02330_),
    .Y(_02331_));
 sky130_fd_sc_hd__o22ai_1 _09180_ (.A1(net144),
    .A2(_00306_),
    .B1(net47),
    .B2(net132),
    .Y(_02332_));
 sky130_fd_sc_hd__xor2_1 _09181_ (.A(net109),
    .B(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__and2b_1 _09182_ (.A_N(_02331_),
    .B(_02333_),
    .X(_02334_));
 sky130_fd_sc_hd__and2b_1 _09183_ (.A_N(_02333_),
    .B(_02331_),
    .X(_02335_));
 sky130_fd_sc_hd__or2_1 _09184_ (.A(_02334_),
    .B(_02335_),
    .X(_02336_));
 sky130_fd_sc_hd__o22a_1 _09185_ (.A1(net53),
    .A2(net147),
    .B1(net141),
    .B2(net14),
    .X(_02337_));
 sky130_fd_sc_hd__xnor2_1 _09186_ (.A(net112),
    .B(_02337_),
    .Y(_02338_));
 sky130_fd_sc_hd__and2b_1 _09187_ (.A_N(_02336_),
    .B(_02338_),
    .X(_02339_));
 sky130_fd_sc_hd__and2b_1 _09188_ (.A_N(_02338_),
    .B(_02336_),
    .X(_02340_));
 sky130_fd_sc_hd__or2_2 _09189_ (.A(_02339_),
    .B(_02340_),
    .X(_02341_));
 sky130_fd_sc_hd__a21oi_2 _09190_ (.A1(_00785_),
    .A2(_02053_),
    .B1(_02055_),
    .Y(_02342_));
 sky130_fd_sc_hd__xnor2_2 _09191_ (.A(_02341_),
    .B(_02342_),
    .Y(_02343_));
 sky130_fd_sc_hd__and2b_1 _09192_ (.A_N(_02343_),
    .B(_02329_),
    .X(_02344_));
 sky130_fd_sc_hd__xor2_4 _09193_ (.A(_02329_),
    .B(_02343_),
    .X(_02345_));
 sky130_fd_sc_hd__nand2_1 _09194_ (.A(_02072_),
    .B(_02076_),
    .Y(_02346_));
 sky130_fd_sc_hd__a21oi_1 _09195_ (.A1(_02106_),
    .A2(_02108_),
    .B1(_02104_),
    .Y(_02347_));
 sky130_fd_sc_hd__o21ba_1 _09196_ (.A1(_02059_),
    .A2(_02065_),
    .B1_N(_02064_),
    .X(_02348_));
 sky130_fd_sc_hd__or2_1 _09197_ (.A(_02347_),
    .B(_02348_),
    .X(_02349_));
 sky130_fd_sc_hd__xnor2_1 _09198_ (.A(_02347_),
    .B(_02348_),
    .Y(_02350_));
 sky130_fd_sc_hd__nand2b_1 _09199_ (.A_N(_02350_),
    .B(_02346_),
    .Y(_02351_));
 sky130_fd_sc_hd__xnor2_1 _09200_ (.A(_02346_),
    .B(_02350_),
    .Y(_02352_));
 sky130_fd_sc_hd__o22a_1 _09201_ (.A1(net152),
    .A2(net58),
    .B1(net55),
    .B2(net150),
    .X(_02353_));
 sky130_fd_sc_hd__xnor2_1 _09202_ (.A(net191),
    .B(_02353_),
    .Y(_02354_));
 sky130_fd_sc_hd__o22a_1 _09203_ (.A1(net116),
    .A2(net68),
    .B1(net65),
    .B2(net114),
    .X(_02355_));
 sky130_fd_sc_hd__xnor2_1 _09204_ (.A(net179),
    .B(_02355_),
    .Y(_02356_));
 sky130_fd_sc_hd__o22a_1 _09205_ (.A1(net177),
    .A2(net63),
    .B1(net60),
    .B2(net175),
    .X(_02357_));
 sky130_fd_sc_hd__xnor2_1 _09206_ (.A(net189),
    .B(_02357_),
    .Y(_02358_));
 sky130_fd_sc_hd__or2_1 _09207_ (.A(_02356_),
    .B(_02358_),
    .X(_02359_));
 sky130_fd_sc_hd__and2_1 _09208_ (.A(_02356_),
    .B(_02358_),
    .X(_02360_));
 sky130_fd_sc_hd__nand2_1 _09209_ (.A(_02356_),
    .B(_02358_),
    .Y(_02361_));
 sky130_fd_sc_hd__nand2_1 _09210_ (.A(_02359_),
    .B(_02361_),
    .Y(_02362_));
 sky130_fd_sc_hd__xnor2_1 _09211_ (.A(_02354_),
    .B(_02362_),
    .Y(_02363_));
 sky130_fd_sc_hd__o22a_1 _09212_ (.A1(net128),
    .A2(net42),
    .B1(net94),
    .B2(net100),
    .X(_02364_));
 sky130_fd_sc_hd__xnor2_1 _09213_ (.A(net138),
    .B(_02364_),
    .Y(_02365_));
 sky130_fd_sc_hd__o22a_1 _09214_ (.A1(net82),
    .A2(net76),
    .B1(net74),
    .B2(net130),
    .X(_02366_));
 sky130_fd_sc_hd__xnor2_1 _09215_ (.A(net157),
    .B(_02366_),
    .Y(_02367_));
 sky130_fd_sc_hd__inv_2 _09216_ (.A(_02367_),
    .Y(_02368_));
 sky130_fd_sc_hd__xnor2_1 _09217_ (.A(_02365_),
    .B(_02367_),
    .Y(_02369_));
 sky130_fd_sc_hd__o22a_1 _09218_ (.A1(net78),
    .A2(net119),
    .B1(net71),
    .B2(net123),
    .X(_02370_));
 sky130_fd_sc_hd__xnor2_1 _09219_ (.A(net154),
    .B(_02370_),
    .Y(_02371_));
 sky130_fd_sc_hd__and2_1 _09220_ (.A(_02369_),
    .B(_02371_),
    .X(_02372_));
 sky130_fd_sc_hd__xor2_1 _09221_ (.A(_02369_),
    .B(_02371_),
    .X(_02373_));
 sky130_fd_sc_hd__o22a_1 _09222_ (.A1(net173),
    .A2(net9),
    .B1(net4),
    .B2(net171),
    .X(_02374_));
 sky130_fd_sc_hd__xnor2_1 _09223_ (.A(_00180_),
    .B(_02374_),
    .Y(_02375_));
 sky130_fd_sc_hd__nand3_1 _09224_ (.A(_00208_),
    .B(_00219_),
    .C(_00221_),
    .Y(_02376_));
 sky130_fd_sc_hd__a21o_1 _09225_ (.A1(_00225_),
    .A2(_00226_),
    .B1(net167),
    .X(_02377_));
 sky130_fd_sc_hd__a21o_1 _09226_ (.A1(_02376_),
    .A2(_02377_),
    .B1(net210),
    .X(_02378_));
 sky130_fd_sc_hd__nand3_1 _09227_ (.A(net210),
    .B(_02376_),
    .C(_02377_),
    .Y(_02379_));
 sky130_fd_sc_hd__and3_1 _09228_ (.A(net256),
    .B(_02378_),
    .C(_02379_),
    .X(_02380_));
 sky130_fd_sc_hd__a21oi_1 _09229_ (.A1(_02378_),
    .A2(_02379_),
    .B1(net256),
    .Y(_02381_));
 sky130_fd_sc_hd__nor3b_1 _09230_ (.A(_02380_),
    .B(_02381_),
    .C_N(_02375_),
    .Y(_02382_));
 sky130_fd_sc_hd__or3b_1 _09231_ (.A(_02380_),
    .B(_02381_),
    .C_N(_02375_),
    .X(_02383_));
 sky130_fd_sc_hd__o21bai_1 _09232_ (.A1(_02380_),
    .A2(_02381_),
    .B1_N(_02375_),
    .Y(_02384_));
 sky130_fd_sc_hd__and3_1 _09233_ (.A(_02373_),
    .B(_02383_),
    .C(_02384_),
    .X(_02385_));
 sky130_fd_sc_hd__a21oi_1 _09234_ (.A1(_02383_),
    .A2(_02384_),
    .B1(_02373_),
    .Y(_02386_));
 sky130_fd_sc_hd__nor3_2 _09235_ (.A(_02363_),
    .B(_02385_),
    .C(_02386_),
    .Y(_02387_));
 sky130_fd_sc_hd__o21a_1 _09236_ (.A1(_02385_),
    .A2(_02386_),
    .B1(_02363_),
    .X(_02388_));
 sky130_fd_sc_hd__nor2_1 _09237_ (.A(net163),
    .B(net32),
    .Y(_02389_));
 sky130_fd_sc_hd__a21oi_2 _09238_ (.A1(_02080_),
    .A2(_02085_),
    .B1(_02084_),
    .Y(_02390_));
 sky130_fd_sc_hd__o22a_1 _09239_ (.A1(net165),
    .A2(net8),
    .B1(net161),
    .B2(net6),
    .X(_02391_));
 sky130_fd_sc_hd__xnor2_1 _09240_ (.A(net31),
    .B(_02391_),
    .Y(_02392_));
 sky130_fd_sc_hd__nor2_1 _09241_ (.A(_02390_),
    .B(_02392_),
    .Y(_02393_));
 sky130_fd_sc_hd__xor2_1 _09242_ (.A(_02390_),
    .B(_02392_),
    .X(_02394_));
 sky130_fd_sc_hd__xnor2_1 _09243_ (.A(_02389_),
    .B(_02394_),
    .Y(_02395_));
 sky130_fd_sc_hd__or3_2 _09244_ (.A(_02387_),
    .B(_02388_),
    .C(_02395_),
    .X(_02396_));
 sky130_fd_sc_hd__o21ai_1 _09245_ (.A1(_02387_),
    .A2(_02388_),
    .B1(_02395_),
    .Y(_02397_));
 sky130_fd_sc_hd__nand3_1 _09246_ (.A(_02352_),
    .B(_02396_),
    .C(_02397_),
    .Y(_02398_));
 sky130_fd_sc_hd__a21o_1 _09247_ (.A1(_02396_),
    .A2(_02397_),
    .B1(_02352_),
    .X(_02399_));
 sky130_fd_sc_hd__and2_1 _09248_ (.A(_02398_),
    .B(_02399_),
    .X(_02400_));
 sky130_fd_sc_hd__a21o_1 _09249_ (.A1(_02040_),
    .A2(_02042_),
    .B1(_02046_),
    .X(_02401_));
 sky130_fd_sc_hd__o22a_1 _09250_ (.A1(net121),
    .A2(net36),
    .B1(net34),
    .B2(net80),
    .X(_02402_));
 sky130_fd_sc_hd__xnor2_1 _09251_ (.A(net135),
    .B(_02402_),
    .Y(_02403_));
 sky130_fd_sc_hd__o22a_1 _09252_ (.A1(net51),
    .A2(net90),
    .B1(net87),
    .B2(net49),
    .X(_02404_));
 sky130_fd_sc_hd__xnor2_1 _09253_ (.A(net106),
    .B(_02404_),
    .Y(_02405_));
 sky130_fd_sc_hd__nand2_1 _09254_ (.A(_02403_),
    .B(_02405_),
    .Y(_02406_));
 sky130_fd_sc_hd__xor2_1 _09255_ (.A(_02403_),
    .B(_02405_),
    .X(_02407_));
 sky130_fd_sc_hd__o22a_1 _09256_ (.A1(net92),
    .A2(net40),
    .B1(net38),
    .B2(net125),
    .X(_02408_));
 sky130_fd_sc_hd__xnor2_1 _09257_ (.A(net102),
    .B(_02408_),
    .Y(_02409_));
 sky130_fd_sc_hd__nand2_1 _09258_ (.A(_02407_),
    .B(_02409_),
    .Y(_02410_));
 sky130_fd_sc_hd__or2_1 _09259_ (.A(_02407_),
    .B(_02409_),
    .X(_02411_));
 sky130_fd_sc_hd__nand2_2 _09260_ (.A(_02410_),
    .B(_02411_),
    .Y(_02412_));
 sky130_fd_sc_hd__a21boi_2 _09261_ (.A1(_02089_),
    .A2(_02094_),
    .B1_N(_02093_),
    .Y(_02413_));
 sky130_fd_sc_hd__nor2_1 _09262_ (.A(_02412_),
    .B(_02413_),
    .Y(_02414_));
 sky130_fd_sc_hd__xor2_2 _09263_ (.A(_02412_),
    .B(_02413_),
    .X(_02415_));
 sky130_fd_sc_hd__xor2_1 _09264_ (.A(_02401_),
    .B(_02415_),
    .X(_02416_));
 sky130_fd_sc_hd__nand2_1 _09265_ (.A(_02400_),
    .B(_02416_),
    .Y(_02417_));
 sky130_fd_sc_hd__or2_1 _09266_ (.A(_02400_),
    .B(_02416_),
    .X(_02418_));
 sky130_fd_sc_hd__nand2_2 _09267_ (.A(_02417_),
    .B(_02418_),
    .Y(_02419_));
 sky130_fd_sc_hd__xor2_4 _09268_ (.A(_02345_),
    .B(_02419_),
    .X(_02420_));
 sky130_fd_sc_hd__a21o_1 _09269_ (.A1(_02052_),
    .A2(_02115_),
    .B1(_02114_),
    .X(_02421_));
 sky130_fd_sc_hd__a21o_2 _09270_ (.A1(_02037_),
    .A2(_02051_),
    .B1(_02049_),
    .X(_02422_));
 sky130_fd_sc_hd__a21o_2 _09271_ (.A1(_02057_),
    .A2(_02097_),
    .B1(_02096_),
    .X(_02423_));
 sky130_fd_sc_hd__a21o_1 _09272_ (.A1(_02099_),
    .A2(_02112_),
    .B1(_02111_),
    .X(_02424_));
 sky130_fd_sc_hd__nand2_1 _09273_ (.A(_02423_),
    .B(_02424_),
    .Y(_02425_));
 sky130_fd_sc_hd__xor2_4 _09274_ (.A(_02423_),
    .B(_02424_),
    .X(_02426_));
 sky130_fd_sc_hd__xnor2_4 _09275_ (.A(_02422_),
    .B(_02426_),
    .Y(_02427_));
 sky130_fd_sc_hd__a21oi_4 _09276_ (.A1(_02119_),
    .A2(_02123_),
    .B1(_02122_),
    .Y(_02428_));
 sky130_fd_sc_hd__xnor2_2 _09277_ (.A(_02427_),
    .B(_02428_),
    .Y(_02429_));
 sky130_fd_sc_hd__nand2b_1 _09278_ (.A_N(_02429_),
    .B(_02421_),
    .Y(_02430_));
 sky130_fd_sc_hd__xnor2_2 _09279_ (.A(_02421_),
    .B(_02429_),
    .Y(_02431_));
 sky130_fd_sc_hd__and2_1 _09280_ (.A(_02420_),
    .B(_02431_),
    .X(_02432_));
 sky130_fd_sc_hd__xor2_4 _09281_ (.A(_02420_),
    .B(_02431_),
    .X(_02433_));
 sky130_fd_sc_hd__xnor2_4 _09282_ (.A(_02328_),
    .B(_02433_),
    .Y(_02434_));
 sky130_fd_sc_hd__xor2_4 _09283_ (.A(_02327_),
    .B(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__a21o_1 _09284_ (.A1(_02035_),
    .A2(_02134_),
    .B1(_02133_),
    .X(_02436_));
 sky130_fd_sc_hd__xnor2_4 _09285_ (.A(_02435_),
    .B(_02436_),
    .Y(_02437_));
 sky130_fd_sc_hd__o21ai_1 _09286_ (.A1(_02135_),
    .A2(_02212_),
    .B1(net22),
    .Y(_02438_));
 sky130_fd_sc_hd__a21oi_1 _09287_ (.A1(_02437_),
    .A2(_02438_),
    .B1(_02214_),
    .Y(_02439_));
 sky130_fd_sc_hd__o21a_1 _09288_ (.A1(_02437_),
    .A2(_02438_),
    .B1(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__mux2_1 _09289_ (.A0(_02268_),
    .A1(_02310_),
    .S(net230),
    .X(_02441_));
 sky130_fd_sc_hd__o21a_1 _09290_ (.A1(net232),
    .A2(_02441_),
    .B1(_02316_),
    .X(_02442_));
 sky130_fd_sc_hd__o21a_1 _09291_ (.A1(net235),
    .A2(_02442_),
    .B1(_02318_),
    .X(_02443_));
 sky130_fd_sc_hd__o21ai_2 _09292_ (.A1(net238),
    .A2(_02443_),
    .B1(_02312_),
    .Y(_02444_));
 sky130_fd_sc_hd__nor2_1 _09293_ (.A(net186),
    .B(_02444_),
    .Y(_02445_));
 sky130_fd_sc_hd__mux2_1 _09294_ (.A0(_02220_),
    .A1(_02223_),
    .S(net227),
    .X(_02446_));
 sky130_fd_sc_hd__mux2_1 _09295_ (.A0(_02222_),
    .A1(_02230_),
    .S(net227),
    .X(_02447_));
 sky130_fd_sc_hd__mux2_1 _09296_ (.A0(_02446_),
    .A1(_02447_),
    .S(net230),
    .X(_02448_));
 sky130_fd_sc_hd__mux2_1 _09297_ (.A0(_02226_),
    .A1(_02245_),
    .S(net227),
    .X(_02449_));
 sky130_fd_sc_hd__mux2_1 _09298_ (.A0(_02227_),
    .A1(_02229_),
    .S(net224),
    .X(_02450_));
 sky130_fd_sc_hd__mux2_1 _09299_ (.A0(_02449_),
    .A1(_02450_),
    .S(net228),
    .X(_02451_));
 sky130_fd_sc_hd__mux2_1 _09300_ (.A0(_02448_),
    .A1(_02451_),
    .S(net231),
    .X(_02452_));
 sky130_fd_sc_hd__mux2_1 _09301_ (.A0(_02234_),
    .A1(_02261_),
    .S(net227),
    .X(_02453_));
 sky130_fd_sc_hd__mux2_1 _09302_ (.A0(_02235_),
    .A1(_02237_),
    .S(net225),
    .X(_02454_));
 sky130_fd_sc_hd__mux2_1 _09303_ (.A0(_02453_),
    .A1(_02454_),
    .S(net228),
    .X(_02455_));
 sky130_fd_sc_hd__mux2_1 _09304_ (.A0(_02238_),
    .A1(_02241_),
    .S(net225),
    .X(_02456_));
 sky130_fd_sc_hd__mux2_1 _09305_ (.A0(_02242_),
    .A1(_02244_),
    .S(net224),
    .X(_02457_));
 sky130_fd_sc_hd__mux2_1 _09306_ (.A0(_02456_),
    .A1(_02457_),
    .S(net228),
    .X(_02458_));
 sky130_fd_sc_hd__mux2_1 _09307_ (.A0(_02458_),
    .A1(_02455_),
    .S(net231),
    .X(_02459_));
 sky130_fd_sc_hd__mux2_1 _09308_ (.A0(_02452_),
    .A1(_02459_),
    .S(net236),
    .X(_02460_));
 sky130_fd_sc_hd__mux2_1 _09309_ (.A0(_02250_),
    .A1(_02277_),
    .S(net227),
    .X(_02461_));
 sky130_fd_sc_hd__mux2_1 _09310_ (.A0(_02251_),
    .A1(_02253_),
    .S(net224),
    .X(_02462_));
 sky130_fd_sc_hd__mux2_1 _09311_ (.A0(_02461_),
    .A1(_02462_),
    .S(net228),
    .X(_02463_));
 sky130_fd_sc_hd__mux2_1 _09312_ (.A0(_02254_),
    .A1(_02257_),
    .S(net225),
    .X(_02464_));
 sky130_fd_sc_hd__mux2_1 _09313_ (.A0(_02258_),
    .A1(_02260_),
    .S(net225),
    .X(_02465_));
 sky130_fd_sc_hd__mux2_1 _09314_ (.A0(_02464_),
    .A1(_02465_),
    .S(net228),
    .X(_02466_));
 sky130_fd_sc_hd__mux2_1 _09315_ (.A0(_02466_),
    .A1(_02463_),
    .S(net231),
    .X(_02467_));
 sky130_fd_sc_hd__mux2_1 _09316_ (.A0(_02267_),
    .A1(_02269_),
    .S(net224),
    .X(_02468_));
 sky130_fd_sc_hd__mux2_1 _09317_ (.A0(_02314_),
    .A1(_02468_),
    .S(net228),
    .X(_02469_));
 sky130_fd_sc_hd__mux2_1 _09318_ (.A0(_02270_),
    .A1(_02273_),
    .S(net224),
    .X(_02470_));
 sky130_fd_sc_hd__mux2_1 _09319_ (.A0(_02274_),
    .A1(_02276_),
    .S(net224),
    .X(_02471_));
 sky130_fd_sc_hd__mux2_1 _09320_ (.A0(_02470_),
    .A1(_02471_),
    .S(net228),
    .X(_02472_));
 sky130_fd_sc_hd__mux2_1 _09321_ (.A0(_02472_),
    .A1(_02469_),
    .S(net233),
    .X(_02473_));
 sky130_fd_sc_hd__mux2_1 _09322_ (.A0(_02467_),
    .A1(_02473_),
    .S(net236),
    .X(_02474_));
 sky130_fd_sc_hd__mux2_1 _09323_ (.A0(_02460_),
    .A1(_02474_),
    .S(net238),
    .X(_02475_));
 sky130_fd_sc_hd__inv_2 _09324_ (.A(_02475_),
    .Y(_02476_));
 sky130_fd_sc_hd__nand2_1 _09325_ (.A(reg1_val[1]),
    .B(curr_PC[1]),
    .Y(_02477_));
 sky130_fd_sc_hd__or2_1 _09326_ (.A(reg1_val[1]),
    .B(curr_PC[1]),
    .X(_02478_));
 sky130_fd_sc_hd__nand2_1 _09327_ (.A(_02477_),
    .B(_02478_),
    .Y(_02479_));
 sky130_fd_sc_hd__xnor2_1 _09328_ (.A(_02284_),
    .B(_02479_),
    .Y(_02480_));
 sky130_fd_sc_hd__a21o_1 _09329_ (.A1(net263),
    .A2(_02480_),
    .B1(net214),
    .X(_02481_));
 sky130_fd_sc_hd__nand2_1 _09330_ (.A(net182),
    .B(_02481_),
    .Y(_02482_));
 sky130_fd_sc_hd__a31o_1 _09331_ (.A1(net306),
    .A2(_04785_),
    .A3(_00187_),
    .B1(_06371_),
    .X(_02483_));
 sky130_fd_sc_hd__a21o_1 _09332_ (.A1(net254),
    .A2(net85),
    .B1(_02483_),
    .X(_02484_));
 sky130_fd_sc_hd__xnor2_1 _09333_ (.A(_01975_),
    .B(_02484_),
    .Y(_02485_));
 sky130_fd_sc_hd__a21oi_1 _09334_ (.A1(\div_res[0] ),
    .A2(net26),
    .B1(\div_res[1] ),
    .Y(_02486_));
 sky130_fd_sc_hd__a31o_1 _09335_ (.A1(\div_res[1] ),
    .A2(\div_res[0] ),
    .A3(net26),
    .B1(net203),
    .X(_02487_));
 sky130_fd_sc_hd__or3_1 _09336_ (.A(net304),
    .B(_06305_),
    .C(net226),
    .X(_02488_));
 sky130_fd_sc_hd__nand2_1 _09337_ (.A(_06310_),
    .B(_02488_),
    .Y(_02489_));
 sky130_fd_sc_hd__o21ai_1 _09338_ (.A1(net305),
    .A2(net226),
    .B1(_02489_),
    .Y(_02490_));
 sky130_fd_sc_hd__o31a_1 _09339_ (.A1(net306),
    .A2(net226),
    .A3(_02489_),
    .B1(net251),
    .X(_02491_));
 sky130_fd_sc_hd__nand2_1 _09340_ (.A(_02490_),
    .B(_02491_),
    .Y(_02492_));
 sky130_fd_sc_hd__o22a_1 _09341_ (.A1(_06303_),
    .A2(_02291_),
    .B1(net204),
    .B2(_06302_),
    .X(_02493_));
 sky130_fd_sc_hd__and2_1 _09342_ (.A(divi1_sign),
    .B(net307),
    .X(_02494_));
 sky130_fd_sc_hd__and3_1 _09343_ (.A(\div_shifter[33] ),
    .B(\div_shifter[32] ),
    .C(net246),
    .X(_02495_));
 sky130_fd_sc_hd__a21oi_1 _09344_ (.A1(\div_shifter[32] ),
    .A2(net247),
    .B1(\div_shifter[33] ),
    .Y(_02496_));
 sky130_fd_sc_hd__o32a_1 _09345_ (.A1(net248),
    .A2(_02495_),
    .A3(_02496_),
    .B1(_06426_),
    .B2(net229),
    .X(_02497_));
 sky130_fd_sc_hd__o211a_1 _09346_ (.A1(net242),
    .A2(_02481_),
    .B1(_02493_),
    .C1(_02497_),
    .X(_02498_));
 sky130_fd_sc_hd__o211a_1 _09347_ (.A1(_06305_),
    .A2(_02295_),
    .B1(_02492_),
    .C1(_02498_),
    .X(_02499_));
 sky130_fd_sc_hd__o21ai_1 _09348_ (.A1(_02486_),
    .A2(_02487_),
    .B1(_02499_),
    .Y(_02500_));
 sky130_fd_sc_hd__a221o_1 _09349_ (.A1(_02475_),
    .A2(_02482_),
    .B1(_02485_),
    .B2(_02298_),
    .C1(_02500_),
    .X(_02501_));
 sky130_fd_sc_hd__o31a_1 _09350_ (.A1(_02440_),
    .A2(_02445_),
    .A3(_02501_),
    .B1(net261),
    .X(_02502_));
 sky130_fd_sc_hd__or2_1 _09351_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .X(_02503_));
 sky130_fd_sc_hd__nand2_1 _09352_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .Y(_02504_));
 sky130_fd_sc_hd__a31o_4 _09353_ (.A1(net262),
    .A2(_02503_),
    .A3(_02504_),
    .B1(_02502_),
    .X(dest_val[1]));
 sky130_fd_sc_hd__a21o_2 _09354_ (.A1(_02328_),
    .A2(_02433_),
    .B1(_02432_),
    .X(_02505_));
 sky130_fd_sc_hd__o21ai_4 _09355_ (.A1(_02427_),
    .A2(_02428_),
    .B1(_02430_),
    .Y(_02506_));
 sky130_fd_sc_hd__nor2_2 _09356_ (.A(_02385_),
    .B(_02387_),
    .Y(_02507_));
 sky130_fd_sc_hd__o22a_1 _09357_ (.A1(net143),
    .A2(net12),
    .B1(net45),
    .B2(net141),
    .X(_02508_));
 sky130_fd_sc_hd__xnor2_1 _09358_ (.A(net97),
    .B(_02508_),
    .Y(_02509_));
 sky130_fd_sc_hd__o22ai_1 _09359_ (.A1(net13),
    .A2(net133),
    .B1(net90),
    .B2(net47),
    .Y(_02510_));
 sky130_fd_sc_hd__xor2_1 _09360_ (.A(net109),
    .B(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__and2b_1 _09361_ (.A_N(_02509_),
    .B(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__and2b_1 _09362_ (.A_N(_02511_),
    .B(_02509_),
    .X(_02513_));
 sky130_fd_sc_hd__or2_1 _09363_ (.A(_02512_),
    .B(_02513_),
    .X(_02514_));
 sky130_fd_sc_hd__o22a_1 _09364_ (.A1(net15),
    .A2(net147),
    .B1(net144),
    .B2(net53),
    .X(_02515_));
 sky130_fd_sc_hd__xnor2_1 _09365_ (.A(net112),
    .B(_02515_),
    .Y(_02516_));
 sky130_fd_sc_hd__and2b_1 _09366_ (.A_N(_02514_),
    .B(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__and2b_1 _09367_ (.A_N(_02516_),
    .B(_02514_),
    .X(_02518_));
 sky130_fd_sc_hd__or2_1 _09368_ (.A(_02517_),
    .B(_02518_),
    .X(_02519_));
 sky130_fd_sc_hd__a21o_1 _09369_ (.A1(_02349_),
    .A2(_02351_),
    .B1(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__nand3_1 _09370_ (.A(_02349_),
    .B(_02351_),
    .C(_02519_),
    .Y(_02521_));
 sky130_fd_sc_hd__nand2_2 _09371_ (.A(_02520_),
    .B(_02521_),
    .Y(_02522_));
 sky130_fd_sc_hd__xor2_4 _09372_ (.A(_02507_),
    .B(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__or2_1 _09373_ (.A(_02334_),
    .B(_02339_),
    .X(_02524_));
 sky130_fd_sc_hd__o22a_1 _09374_ (.A1(net49),
    .A2(net92),
    .B1(net88),
    .B2(net51),
    .X(_02525_));
 sky130_fd_sc_hd__xnor2_1 _09375_ (.A(net106),
    .B(_02525_),
    .Y(_02526_));
 sky130_fd_sc_hd__o22a_1 _09376_ (.A1(net80),
    .A2(net36),
    .B1(net34),
    .B2(net128),
    .X(_02527_));
 sky130_fd_sc_hd__xnor2_1 _09377_ (.A(net135),
    .B(_02527_),
    .Y(_02528_));
 sky130_fd_sc_hd__nand2_1 _09378_ (.A(_02526_),
    .B(_02528_),
    .Y(_02529_));
 sky130_fd_sc_hd__xor2_1 _09379_ (.A(_02526_),
    .B(_02528_),
    .X(_02530_));
 sky130_fd_sc_hd__o22a_1 _09380_ (.A1(net126),
    .A2(net40),
    .B1(net38),
    .B2(net121),
    .X(_02531_));
 sky130_fd_sc_hd__xnor2_1 _09381_ (.A(net102),
    .B(_02531_),
    .Y(_02532_));
 sky130_fd_sc_hd__nand2_1 _09382_ (.A(_02530_),
    .B(_02532_),
    .Y(_02533_));
 sky130_fd_sc_hd__or2_1 _09383_ (.A(_02530_),
    .B(_02532_),
    .X(_02534_));
 sky130_fd_sc_hd__nand2_1 _09384_ (.A(_02533_),
    .B(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__a21oi_1 _09385_ (.A1(_02389_),
    .A2(_02394_),
    .B1(_02393_),
    .Y(_02536_));
 sky130_fd_sc_hd__or2_1 _09386_ (.A(_02535_),
    .B(_02536_),
    .X(_02537_));
 sky130_fd_sc_hd__xor2_1 _09387_ (.A(_02535_),
    .B(_02536_),
    .X(_02538_));
 sky130_fd_sc_hd__nand2_1 _09388_ (.A(_02524_),
    .B(_02538_),
    .Y(_02539_));
 sky130_fd_sc_hd__or2_1 _09389_ (.A(_02524_),
    .B(_02538_),
    .X(_02540_));
 sky130_fd_sc_hd__nand2_1 _09390_ (.A(_02539_),
    .B(_02540_),
    .Y(_02541_));
 sky130_fd_sc_hd__a21o_1 _09391_ (.A1(_02365_),
    .A2(_02368_),
    .B1(_02372_),
    .X(_02542_));
 sky130_fd_sc_hd__o21a_1 _09392_ (.A1(_02354_),
    .A2(_02360_),
    .B1(_02359_),
    .X(_02543_));
 sky130_fd_sc_hd__a21oi_1 _09393_ (.A1(_02406_),
    .A2(_02410_),
    .B1(_02543_),
    .Y(_02544_));
 sky130_fd_sc_hd__and3_1 _09394_ (.A(_02406_),
    .B(_02410_),
    .C(_02543_),
    .X(_02545_));
 sky130_fd_sc_hd__nor2_1 _09395_ (.A(_02544_),
    .B(_02545_),
    .Y(_02546_));
 sky130_fd_sc_hd__xor2_1 _09396_ (.A(_02542_),
    .B(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__o22a_1 _09397_ (.A1(net150),
    .A2(net63),
    .B1(net55),
    .B2(net152),
    .X(_02548_));
 sky130_fd_sc_hd__xnor2_1 _09398_ (.A(net191),
    .B(_02548_),
    .Y(_02549_));
 sky130_fd_sc_hd__inv_2 _09399_ (.A(_02549_),
    .Y(_02550_));
 sky130_fd_sc_hd__o22ai_2 _09400_ (.A1(net177),
    .A2(net60),
    .B1(_00223_),
    .B2(net175),
    .Y(_02551_));
 sky130_fd_sc_hd__xor2_2 _09401_ (.A(net189),
    .B(_02551_),
    .X(_02552_));
 sky130_fd_sc_hd__o22a_1 _09402_ (.A1(net116),
    .A2(net64),
    .B1(net58),
    .B2(net114),
    .X(_02553_));
 sky130_fd_sc_hd__xnor2_2 _09403_ (.A(net179),
    .B(_02553_),
    .Y(_02554_));
 sky130_fd_sc_hd__nor2_1 _09404_ (.A(_02552_),
    .B(_02554_),
    .Y(_02555_));
 sky130_fd_sc_hd__xor2_2 _09405_ (.A(_02552_),
    .B(_02554_),
    .X(_02556_));
 sky130_fd_sc_hd__xnor2_2 _09406_ (.A(_02550_),
    .B(_02556_),
    .Y(_02557_));
 sky130_fd_sc_hd__o22a_1 _09407_ (.A1(net99),
    .A2(net42),
    .B1(net94),
    .B2(net118),
    .X(_02558_));
 sky130_fd_sc_hd__xnor2_1 _09408_ (.A(net138),
    .B(_02558_),
    .Y(_02559_));
 sky130_fd_sc_hd__o22a_1 _09409_ (.A1(net82),
    .A2(net74),
    .B1(net68),
    .B2(net130),
    .X(_02560_));
 sky130_fd_sc_hd__xnor2_2 _09410_ (.A(net157),
    .B(_02560_),
    .Y(_02561_));
 sky130_fd_sc_hd__inv_2 _09411_ (.A(_02561_),
    .Y(_02562_));
 sky130_fd_sc_hd__xnor2_1 _09412_ (.A(_02559_),
    .B(_02561_),
    .Y(_02563_));
 sky130_fd_sc_hd__o22a_1 _09413_ (.A1(net123),
    .A2(net77),
    .B1(net70),
    .B2(net78),
    .X(_02564_));
 sky130_fd_sc_hd__xnor2_1 _09414_ (.A(net154),
    .B(_02564_),
    .Y(_02565_));
 sky130_fd_sc_hd__and2_1 _09415_ (.A(_02563_),
    .B(_02565_),
    .X(_02566_));
 sky130_fd_sc_hd__nor2_1 _09416_ (.A(_02563_),
    .B(_02565_),
    .Y(_02567_));
 sky130_fd_sc_hd__nor2_1 _09417_ (.A(_02566_),
    .B(_02567_),
    .Y(_02568_));
 sky130_fd_sc_hd__o22a_1 _09418_ (.A1(net169),
    .A2(net17),
    .B1(net9),
    .B2(net167),
    .X(_02569_));
 sky130_fd_sc_hd__xnor2_2 _09419_ (.A(net210),
    .B(_02569_),
    .Y(_02570_));
 sky130_fd_sc_hd__nor2_1 _09420_ (.A(net255),
    .B(_02570_),
    .Y(_02571_));
 sky130_fd_sc_hd__xnor2_2 _09421_ (.A(net256),
    .B(_02570_),
    .Y(_02572_));
 sky130_fd_sc_hd__nor2_1 _09422_ (.A(net173),
    .B(net4),
    .Y(_02573_));
 sky130_fd_sc_hd__xnor2_2 _09423_ (.A(net208),
    .B(_02573_),
    .Y(_02574_));
 sky130_fd_sc_hd__xor2_2 _09424_ (.A(_02572_),
    .B(_02574_),
    .X(_02575_));
 sky130_fd_sc_hd__nand2_1 _09425_ (.A(_02568_),
    .B(_02575_),
    .Y(_02576_));
 sky130_fd_sc_hd__xnor2_2 _09426_ (.A(_02568_),
    .B(_02575_),
    .Y(_02577_));
 sky130_fd_sc_hd__xnor2_2 _09427_ (.A(_02557_),
    .B(_02577_),
    .Y(_02578_));
 sky130_fd_sc_hd__nor2_1 _09428_ (.A(net161),
    .B(net31),
    .Y(_02579_));
 sky130_fd_sc_hd__o22a_1 _09429_ (.A1(net149),
    .A2(net8),
    .B1(net6),
    .B2(net165),
    .X(_02580_));
 sky130_fd_sc_hd__xnor2_1 _09430_ (.A(net33),
    .B(_02580_),
    .Y(_02581_));
 sky130_fd_sc_hd__o21ai_1 _09431_ (.A1(_02380_),
    .A2(_02382_),
    .B1(_02581_),
    .Y(_02582_));
 sky130_fd_sc_hd__or3_1 _09432_ (.A(_02380_),
    .B(_02382_),
    .C(_02581_),
    .X(_02583_));
 sky130_fd_sc_hd__and2_1 _09433_ (.A(_02582_),
    .B(_02583_),
    .X(_02584_));
 sky130_fd_sc_hd__xnor2_2 _09434_ (.A(_02579_),
    .B(_02584_),
    .Y(_02585_));
 sky130_fd_sc_hd__nor2_1 _09435_ (.A(_02578_),
    .B(_02585_),
    .Y(_02586_));
 sky130_fd_sc_hd__xor2_2 _09436_ (.A(_02578_),
    .B(_02585_),
    .X(_02587_));
 sky130_fd_sc_hd__xnor2_1 _09437_ (.A(_02547_),
    .B(_02587_),
    .Y(_02588_));
 sky130_fd_sc_hd__nor2_1 _09438_ (.A(_02541_),
    .B(_02588_),
    .Y(_02589_));
 sky130_fd_sc_hd__nand2_1 _09439_ (.A(_02541_),
    .B(_02588_),
    .Y(_02590_));
 sky130_fd_sc_hd__and2b_1 _09440_ (.A_N(_02589_),
    .B(_02590_),
    .X(_02591_));
 sky130_fd_sc_hd__xor2_4 _09441_ (.A(_02523_),
    .B(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__o21ai_4 _09442_ (.A1(_02345_),
    .A2(_02419_),
    .B1(_02417_),
    .Y(_02593_));
 sky130_fd_sc_hd__o21bai_2 _09443_ (.A1(_02341_),
    .A2(_02342_),
    .B1_N(_02344_),
    .Y(_02594_));
 sky130_fd_sc_hd__nand2_1 _09444_ (.A(_02396_),
    .B(_02398_),
    .Y(_02595_));
 sky130_fd_sc_hd__a21oi_2 _09445_ (.A1(_02401_),
    .A2(_02415_),
    .B1(_02414_),
    .Y(_02596_));
 sky130_fd_sc_hd__a21oi_1 _09446_ (.A1(_02396_),
    .A2(_02398_),
    .B1(_02596_),
    .Y(_02597_));
 sky130_fd_sc_hd__xnor2_2 _09447_ (.A(_02595_),
    .B(_02596_),
    .Y(_02598_));
 sky130_fd_sc_hd__xnor2_2 _09448_ (.A(_02594_),
    .B(_02598_),
    .Y(_02599_));
 sky130_fd_sc_hd__a21boi_2 _09449_ (.A1(_02422_),
    .A2(_02426_),
    .B1_N(_02425_),
    .Y(_02600_));
 sky130_fd_sc_hd__xnor2_2 _09450_ (.A(_02599_),
    .B(_02600_),
    .Y(_02601_));
 sky130_fd_sc_hd__nand2b_1 _09451_ (.A_N(_02601_),
    .B(_02593_),
    .Y(_02602_));
 sky130_fd_sc_hd__xnor2_4 _09452_ (.A(_02593_),
    .B(_02601_),
    .Y(_02603_));
 sky130_fd_sc_hd__nand2_1 _09453_ (.A(_02592_),
    .B(_02603_),
    .Y(_02604_));
 sky130_fd_sc_hd__xor2_4 _09454_ (.A(_02592_),
    .B(_02603_),
    .X(_02605_));
 sky130_fd_sc_hd__nand2_1 _09455_ (.A(_02506_),
    .B(_02605_),
    .Y(_02606_));
 sky130_fd_sc_hd__xnor2_4 _09456_ (.A(_02506_),
    .B(_02605_),
    .Y(_02607_));
 sky130_fd_sc_hd__nand2b_1 _09457_ (.A_N(_02607_),
    .B(_02505_),
    .Y(_02608_));
 sky130_fd_sc_hd__xnor2_4 _09458_ (.A(_02505_),
    .B(_02607_),
    .Y(_02609_));
 sky130_fd_sc_hd__o22a_1 _09459_ (.A1(_02131_),
    .A2(_02132_),
    .B1(_02327_),
    .B2(_02434_),
    .X(_02610_));
 sky130_fd_sc_hd__a21oi_1 _09460_ (.A1(_02327_),
    .A2(_02434_),
    .B1(_02610_),
    .Y(_02611_));
 sky130_fd_sc_hd__and2_1 _09461_ (.A(_02134_),
    .B(_02435_),
    .X(_02612_));
 sky130_fd_sc_hd__a21o_2 _09462_ (.A1(_02035_),
    .A2(_02612_),
    .B1(_02611_),
    .X(_02613_));
 sky130_fd_sc_hd__xnor2_4 _09463_ (.A(_02609_),
    .B(_02613_),
    .Y(_02614_));
 sky130_fd_sc_hd__or3b_1 _09464_ (.A(_02135_),
    .B(_02212_),
    .C_N(_02437_),
    .X(_02615_));
 sky130_fd_sc_hd__nand2_1 _09465_ (.A(net22),
    .B(_02615_),
    .Y(_02616_));
 sky130_fd_sc_hd__o21ai_1 _09466_ (.A1(_02614_),
    .A2(_02616_),
    .B1(net206),
    .Y(_02617_));
 sky130_fd_sc_hd__a21o_1 _09467_ (.A1(_02614_),
    .A2(_02616_),
    .B1(_02617_),
    .X(_02618_));
 sky130_fd_sc_hd__a21oi_1 _09468_ (.A1(_01976_),
    .A2(net20),
    .B1(_02167_),
    .Y(_02619_));
 sky130_fd_sc_hd__a311o_1 _09469_ (.A1(_01974_),
    .A2(_01976_),
    .A3(net20),
    .B1(net250),
    .C1(_02619_),
    .X(_02620_));
 sky130_fd_sc_hd__o21ai_1 _09470_ (.A1(net231),
    .A2(_02469_),
    .B1(_02316_),
    .Y(_02621_));
 sky130_fd_sc_hd__inv_2 _09471_ (.A(_02621_),
    .Y(_02622_));
 sky130_fd_sc_hd__o21a_1 _09472_ (.A1(net235),
    .A2(_02622_),
    .B1(_02318_),
    .X(_02623_));
 sky130_fd_sc_hd__inv_2 _09473_ (.A(_02623_),
    .Y(_02624_));
 sky130_fd_sc_hd__o21a_1 _09474_ (.A1(net238),
    .A2(_02623_),
    .B1(_02312_),
    .X(_02625_));
 sky130_fd_sc_hd__mux2_1 _09475_ (.A0(_02224_),
    .A1(_02231_),
    .S(net230),
    .X(_02626_));
 sky130_fd_sc_hd__mux2_1 _09476_ (.A0(_02228_),
    .A1(_02246_),
    .S(net230),
    .X(_02627_));
 sky130_fd_sc_hd__mux2_1 _09477_ (.A0(_02626_),
    .A1(_02627_),
    .S(net232),
    .X(_02628_));
 sky130_fd_sc_hd__mux2_1 _09478_ (.A0(_02236_),
    .A1(_02262_),
    .S(net230),
    .X(_02629_));
 sky130_fd_sc_hd__mux2_1 _09479_ (.A0(_02239_),
    .A1(_02243_),
    .S(net229),
    .X(_02630_));
 sky130_fd_sc_hd__mux2_1 _09480_ (.A0(_02630_),
    .A1(_02629_),
    .S(net232),
    .X(_02631_));
 sky130_fd_sc_hd__mux2_1 _09481_ (.A0(_02628_),
    .A1(_02631_),
    .S(net234),
    .X(_02632_));
 sky130_fd_sc_hd__mux2_1 _09482_ (.A0(_02252_),
    .A1(_02278_),
    .S(net230),
    .X(_02633_));
 sky130_fd_sc_hd__mux2_1 _09483_ (.A0(_02255_),
    .A1(_02259_),
    .S(net228),
    .X(_02634_));
 sky130_fd_sc_hd__mux2_1 _09484_ (.A0(_02634_),
    .A1(_02633_),
    .S(net232),
    .X(_02635_));
 sky130_fd_sc_hd__mux2_1 _09485_ (.A0(_02271_),
    .A1(_02275_),
    .S(net228),
    .X(_02636_));
 sky130_fd_sc_hd__mux2_1 _09486_ (.A0(_02636_),
    .A1(_02441_),
    .S(net233),
    .X(_02637_));
 sky130_fd_sc_hd__mux2_1 _09487_ (.A0(_02635_),
    .A1(_02637_),
    .S(net234),
    .X(_02638_));
 sky130_fd_sc_hd__mux2_2 _09488_ (.A0(_02632_),
    .A1(_02638_),
    .S(net238),
    .X(_02639_));
 sky130_fd_sc_hd__o21a_1 _09489_ (.A1(_02284_),
    .A2(_02479_),
    .B1(_02477_),
    .X(_02640_));
 sky130_fd_sc_hd__nor2_1 _09490_ (.A(reg1_val[2]),
    .B(curr_PC[2]),
    .Y(_02641_));
 sky130_fd_sc_hd__nand2_1 _09491_ (.A(reg1_val[2]),
    .B(curr_PC[2]),
    .Y(_02642_));
 sky130_fd_sc_hd__nand2b_1 _09492_ (.A_N(_02641_),
    .B(_02642_),
    .Y(_02643_));
 sky130_fd_sc_hd__xor2_1 _09493_ (.A(_02640_),
    .B(_02643_),
    .X(_02644_));
 sky130_fd_sc_hd__a21oi_1 _09494_ (.A1(_06302_),
    .A2(_06371_),
    .B1(_06303_),
    .Y(_02645_));
 sky130_fd_sc_hd__and3_1 _09495_ (.A(net307),
    .B(_06301_),
    .C(_06310_),
    .X(_02646_));
 sky130_fd_sc_hd__a21o_1 _09496_ (.A1(net300),
    .A2(_02645_),
    .B1(_02646_),
    .X(_02647_));
 sky130_fd_sc_hd__xor2_1 _09497_ (.A(_06295_),
    .B(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__nor2_1 _09498_ (.A(_02293_),
    .B(_02648_),
    .Y(_02649_));
 sky130_fd_sc_hd__o21ai_1 _09499_ (.A1(\div_res[1] ),
    .A2(\div_res[0] ),
    .B1(net26),
    .Y(_02650_));
 sky130_fd_sc_hd__xnor2_1 _09500_ (.A(\div_res[2] ),
    .B(_02650_),
    .Y(_02651_));
 sky130_fd_sc_hd__nor2_1 _09501_ (.A(_06295_),
    .B(_02295_),
    .Y(_02652_));
 sky130_fd_sc_hd__o21ai_1 _09502_ (.A1(\div_shifter[33] ),
    .A2(\div_shifter[32] ),
    .B1(net246),
    .Y(_02653_));
 sky130_fd_sc_hd__xnor2_1 _09503_ (.A(\div_shifter[34] ),
    .B(_02653_),
    .Y(_02654_));
 sky130_fd_sc_hd__a22o_1 _09504_ (.A1(net233),
    .A2(net213),
    .B1(_02303_),
    .B2(_02654_),
    .X(_02655_));
 sky130_fd_sc_hd__o21a_1 _09505_ (.A1(reg1_val[2]),
    .A2(net233),
    .B1(net205),
    .X(_02656_));
 sky130_fd_sc_hd__mux2_1 _09506_ (.A0(_02625_),
    .A1(_02639_),
    .S(net299),
    .X(_02657_));
 sky130_fd_sc_hd__mux2_1 _09507_ (.A0(_02639_),
    .A1(_02644_),
    .S(net263),
    .X(_02658_));
 sky130_fd_sc_hd__a311o_1 _09508_ (.A1(reg1_val[2]),
    .A2(net233),
    .A3(_02300_),
    .B1(_02655_),
    .C1(_02656_),
    .X(_02659_));
 sky130_fd_sc_hd__a211o_1 _09509_ (.A1(_02305_),
    .A2(_02651_),
    .B1(_02652_),
    .C1(_02659_),
    .X(_02660_));
 sky130_fd_sc_hd__a211o_1 _09510_ (.A1(net215),
    .A2(_02658_),
    .B1(_02660_),
    .C1(_02649_),
    .X(_02661_));
 sky130_fd_sc_hd__a21oi_1 _09511_ (.A1(_06416_),
    .A2(_02657_),
    .B1(_02661_),
    .Y(_02662_));
 sky130_fd_sc_hd__a31o_2 _09512_ (.A1(_02618_),
    .A2(_02620_),
    .A3(_02662_),
    .B1(_06390_),
    .X(_02663_));
 sky130_fd_sc_hd__and3_1 _09513_ (.A(curr_PC[0]),
    .B(curr_PC[1]),
    .C(curr_PC[2]),
    .X(_02664_));
 sky130_fd_sc_hd__a21oi_1 _09514_ (.A1(curr_PC[0]),
    .A2(curr_PC[1]),
    .B1(curr_PC[2]),
    .Y(_02665_));
 sky130_fd_sc_hd__o31ai_4 _09515_ (.A1(net257),
    .A2(_02664_),
    .A3(_02665_),
    .B1(_02663_),
    .Y(dest_val[2]));
 sky130_fd_sc_hd__o21ai_1 _09516_ (.A1(_02599_),
    .A2(_02600_),
    .B1(_02602_),
    .Y(_02666_));
 sky130_fd_sc_hd__o21ai_2 _09517_ (.A1(_02557_),
    .A2(_02577_),
    .B1(_02576_),
    .Y(_02667_));
 sky130_fd_sc_hd__o22a_1 _09518_ (.A1(net141),
    .A2(net12),
    .B1(net45),
    .B2(net147),
    .X(_02668_));
 sky130_fd_sc_hd__xnor2_1 _09519_ (.A(net97),
    .B(_02668_),
    .Y(_02669_));
 sky130_fd_sc_hd__inv_2 _09520_ (.A(_02669_),
    .Y(_02670_));
 sky130_fd_sc_hd__o22ai_2 _09521_ (.A1(net13),
    .A2(net90),
    .B1(net88),
    .B2(_00309_),
    .Y(_02671_));
 sky130_fd_sc_hd__xor2_1 _09522_ (.A(net109),
    .B(_02671_),
    .X(_02672_));
 sky130_fd_sc_hd__xor2_1 _09523_ (.A(_02669_),
    .B(_02672_),
    .X(_02673_));
 sky130_fd_sc_hd__o22a_1 _09524_ (.A1(net15),
    .A2(net144),
    .B1(net133),
    .B2(net52),
    .X(_02674_));
 sky130_fd_sc_hd__xnor2_1 _09525_ (.A(net112),
    .B(_02674_),
    .Y(_02675_));
 sky130_fd_sc_hd__and2b_1 _09526_ (.A_N(_02673_),
    .B(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__and2b_1 _09527_ (.A_N(_02675_),
    .B(_02673_),
    .X(_02677_));
 sky130_fd_sc_hd__or2_2 _09528_ (.A(_02676_),
    .B(_02677_),
    .X(_02678_));
 sky130_fd_sc_hd__a21oi_2 _09529_ (.A1(_02542_),
    .A2(_02546_),
    .B1(_02544_),
    .Y(_02679_));
 sky130_fd_sc_hd__xnor2_1 _09530_ (.A(_02678_),
    .B(_02679_),
    .Y(_02680_));
 sky130_fd_sc_hd__nand2b_1 _09531_ (.A_N(_02680_),
    .B(_02667_),
    .Y(_02681_));
 sky130_fd_sc_hd__xnor2_1 _09532_ (.A(_02667_),
    .B(_02680_),
    .Y(_02682_));
 sky130_fd_sc_hd__a21o_1 _09533_ (.A1(_02559_),
    .A2(_02562_),
    .B1(_02566_),
    .X(_02683_));
 sky130_fd_sc_hd__nand2_1 _09534_ (.A(_02529_),
    .B(_02533_),
    .Y(_02684_));
 sky130_fd_sc_hd__a21oi_2 _09535_ (.A1(_02550_),
    .A2(_02556_),
    .B1(_02555_),
    .Y(_02685_));
 sky130_fd_sc_hd__a21oi_1 _09536_ (.A1(_02529_),
    .A2(_02533_),
    .B1(_02685_),
    .Y(_02686_));
 sky130_fd_sc_hd__xnor2_2 _09537_ (.A(_02684_),
    .B(_02685_),
    .Y(_02687_));
 sky130_fd_sc_hd__xor2_1 _09538_ (.A(_02683_),
    .B(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__o22a_1 _09539_ (.A1(net152),
    .A2(net63),
    .B1(net60),
    .B2(net150),
    .X(_02689_));
 sky130_fd_sc_hd__xnor2_2 _09540_ (.A(net191),
    .B(_02689_),
    .Y(_02690_));
 sky130_fd_sc_hd__o22a_1 _09541_ (.A1(net116),
    .A2(net58),
    .B1(net55),
    .B2(net114),
    .X(_02691_));
 sky130_fd_sc_hd__xor2_1 _09542_ (.A(net179),
    .B(_02691_),
    .X(_02692_));
 sky130_fd_sc_hd__nand3b_1 _09543_ (.A_N(net177),
    .B(_00219_),
    .C(_00221_),
    .Y(_02693_));
 sky130_fd_sc_hd__a21o_1 _09544_ (.A1(_00225_),
    .A2(_00226_),
    .B1(net175),
    .X(_02694_));
 sky130_fd_sc_hd__a21o_1 _09545_ (.A1(_02693_),
    .A2(_02694_),
    .B1(net189),
    .X(_02695_));
 sky130_fd_sc_hd__nand3_1 _09546_ (.A(net189),
    .B(_02693_),
    .C(_02694_),
    .Y(_02696_));
 sky130_fd_sc_hd__and3_1 _09547_ (.A(_02692_),
    .B(_02695_),
    .C(_02696_),
    .X(_02697_));
 sky130_fd_sc_hd__a21oi_1 _09548_ (.A1(_02695_),
    .A2(_02696_),
    .B1(_02692_),
    .Y(_02698_));
 sky130_fd_sc_hd__nor2_1 _09549_ (.A(_02697_),
    .B(_02698_),
    .Y(_02699_));
 sky130_fd_sc_hd__xnor2_2 _09550_ (.A(_02690_),
    .B(_02699_),
    .Y(_02700_));
 sky130_fd_sc_hd__o22a_1 _09551_ (.A1(net82),
    .A2(net68),
    .B1(net65),
    .B2(net130),
    .X(_02701_));
 sky130_fd_sc_hd__xnor2_1 _09552_ (.A(net157),
    .B(_02701_),
    .Y(_02702_));
 sky130_fd_sc_hd__o22a_1 _09553_ (.A1(net119),
    .A2(net42),
    .B1(net94),
    .B2(net71),
    .X(_02703_));
 sky130_fd_sc_hd__xnor2_1 _09554_ (.A(net138),
    .B(_02703_),
    .Y(_02704_));
 sky130_fd_sc_hd__nand2b_1 _09555_ (.A_N(_02702_),
    .B(_02704_),
    .Y(_02705_));
 sky130_fd_sc_hd__xor2_1 _09556_ (.A(_02702_),
    .B(_02704_),
    .X(_02706_));
 sky130_fd_sc_hd__o22a_1 _09557_ (.A1(net78),
    .A2(net77),
    .B1(net74),
    .B2(net123),
    .X(_02707_));
 sky130_fd_sc_hd__xor2_1 _09558_ (.A(net154),
    .B(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__xnor2_1 _09559_ (.A(_02706_),
    .B(_02708_),
    .Y(_02709_));
 sky130_fd_sc_hd__o22a_1 _09560_ (.A1(net169),
    .A2(net9),
    .B1(net4),
    .B2(_00209_),
    .X(_02710_));
 sky130_fd_sc_hd__xnor2_1 _09561_ (.A(net210),
    .B(_02710_),
    .Y(_02711_));
 sky130_fd_sc_hd__or2_1 _09562_ (.A(net256),
    .B(_02711_),
    .X(_02712_));
 sky130_fd_sc_hd__xnor2_2 _09563_ (.A(net256),
    .B(_02711_),
    .Y(_02713_));
 sky130_fd_sc_hd__xnor2_2 _09564_ (.A(_00180_),
    .B(_02713_),
    .Y(_02714_));
 sky130_fd_sc_hd__nor2_1 _09565_ (.A(_02709_),
    .B(_02714_),
    .Y(_02715_));
 sky130_fd_sc_hd__xor2_1 _09566_ (.A(_02709_),
    .B(_02714_),
    .X(_02716_));
 sky130_fd_sc_hd__xnor2_1 _09567_ (.A(_02700_),
    .B(_02716_),
    .Y(_02717_));
 sky130_fd_sc_hd__nor2_1 _09568_ (.A(net165),
    .B(net31),
    .Y(_02718_));
 sky130_fd_sc_hd__a21oi_2 _09569_ (.A1(_02572_),
    .A2(_02574_),
    .B1(_02571_),
    .Y(_02719_));
 sky130_fd_sc_hd__o22a_1 _09570_ (.A1(net143),
    .A2(net8),
    .B1(net6),
    .B2(net149),
    .X(_02720_));
 sky130_fd_sc_hd__xnor2_1 _09571_ (.A(net31),
    .B(_02720_),
    .Y(_02721_));
 sky130_fd_sc_hd__nor2_1 _09572_ (.A(_02719_),
    .B(_02721_),
    .Y(_02722_));
 sky130_fd_sc_hd__xor2_1 _09573_ (.A(_02719_),
    .B(_02721_),
    .X(_02723_));
 sky130_fd_sc_hd__xnor2_1 _09574_ (.A(_02718_),
    .B(_02723_),
    .Y(_02724_));
 sky130_fd_sc_hd__nor2_1 _09575_ (.A(_02717_),
    .B(_02724_),
    .Y(_02725_));
 sky130_fd_sc_hd__xor2_1 _09576_ (.A(_02717_),
    .B(_02724_),
    .X(_02726_));
 sky130_fd_sc_hd__xor2_1 _09577_ (.A(_02688_),
    .B(_02726_),
    .X(_02727_));
 sky130_fd_sc_hd__nor2_1 _09578_ (.A(_02512_),
    .B(_02517_),
    .Y(_02728_));
 sky130_fd_sc_hd__o22a_1 _09579_ (.A1(net128),
    .A2(net36),
    .B1(net34),
    .B2(net99),
    .X(_02729_));
 sky130_fd_sc_hd__xnor2_1 _09580_ (.A(net135),
    .B(_02729_),
    .Y(_02730_));
 sky130_fd_sc_hd__o22a_1 _09581_ (.A1(net126),
    .A2(net49),
    .B1(net92),
    .B2(net50),
    .X(_02731_));
 sky130_fd_sc_hd__xnor2_1 _09582_ (.A(net106),
    .B(_02731_),
    .Y(_02732_));
 sky130_fd_sc_hd__and2_1 _09583_ (.A(_02730_),
    .B(_02732_),
    .X(_02733_));
 sky130_fd_sc_hd__xor2_1 _09584_ (.A(_02730_),
    .B(_02732_),
    .X(_02734_));
 sky130_fd_sc_hd__o22a_1 _09585_ (.A1(net121),
    .A2(net40),
    .B1(net38),
    .B2(net80),
    .X(_02735_));
 sky130_fd_sc_hd__xnor2_1 _09586_ (.A(net102),
    .B(_02735_),
    .Y(_02736_));
 sky130_fd_sc_hd__xnor2_1 _09587_ (.A(_02734_),
    .B(_02736_),
    .Y(_02737_));
 sky130_fd_sc_hd__a21boi_2 _09588_ (.A1(_02579_),
    .A2(_02583_),
    .B1_N(_02582_),
    .Y(_02738_));
 sky130_fd_sc_hd__nor2_1 _09589_ (.A(_02737_),
    .B(_02738_),
    .Y(_02739_));
 sky130_fd_sc_hd__xor2_1 _09590_ (.A(_02737_),
    .B(_02738_),
    .X(_02740_));
 sky130_fd_sc_hd__and2b_1 _09591_ (.A_N(_02728_),
    .B(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__xnor2_1 _09592_ (.A(_02728_),
    .B(_02740_),
    .Y(_02742_));
 sky130_fd_sc_hd__and2_1 _09593_ (.A(_02727_),
    .B(_02742_),
    .X(_02743_));
 sky130_fd_sc_hd__nor2_1 _09594_ (.A(_02727_),
    .B(_02742_),
    .Y(_02744_));
 sky130_fd_sc_hd__nor2_1 _09595_ (.A(_02743_),
    .B(_02744_),
    .Y(_02745_));
 sky130_fd_sc_hd__xor2_1 _09596_ (.A(_02682_),
    .B(_02745_),
    .X(_02746_));
 sky130_fd_sc_hd__a21o_1 _09597_ (.A1(_02523_),
    .A2(_02590_),
    .B1(_02589_),
    .X(_02747_));
 sky130_fd_sc_hd__a21o_1 _09598_ (.A1(_02594_),
    .A2(_02598_),
    .B1(_02597_),
    .X(_02748_));
 sky130_fd_sc_hd__o21ai_2 _09599_ (.A1(_02507_),
    .A2(_02522_),
    .B1(_02520_),
    .Y(_02749_));
 sky130_fd_sc_hd__nand2_1 _09600_ (.A(_02537_),
    .B(_02539_),
    .Y(_02750_));
 sky130_fd_sc_hd__a21oi_2 _09601_ (.A1(_02547_),
    .A2(_02587_),
    .B1(_02586_),
    .Y(_02751_));
 sky130_fd_sc_hd__a21oi_1 _09602_ (.A1(_02537_),
    .A2(_02539_),
    .B1(_02751_),
    .Y(_02752_));
 sky130_fd_sc_hd__xnor2_2 _09603_ (.A(_02750_),
    .B(_02751_),
    .Y(_02753_));
 sky130_fd_sc_hd__xor2_1 _09604_ (.A(_02749_),
    .B(_02753_),
    .X(_02754_));
 sky130_fd_sc_hd__xnor2_1 _09605_ (.A(_02748_),
    .B(_02754_),
    .Y(_02755_));
 sky130_fd_sc_hd__nand2b_1 _09606_ (.A_N(_02755_),
    .B(_02747_),
    .Y(_02756_));
 sky130_fd_sc_hd__xnor2_1 _09607_ (.A(_02747_),
    .B(_02755_),
    .Y(_02757_));
 sky130_fd_sc_hd__and2_1 _09608_ (.A(_02746_),
    .B(_02757_),
    .X(_02758_));
 sky130_fd_sc_hd__xor2_1 _09609_ (.A(_02746_),
    .B(_02757_),
    .X(_02759_));
 sky130_fd_sc_hd__xnor2_1 _09610_ (.A(_02666_),
    .B(_02759_),
    .Y(_02760_));
 sky130_fd_sc_hd__a21oi_1 _09611_ (.A1(_02604_),
    .A2(_02606_),
    .B1(_02760_),
    .Y(_02761_));
 sky130_fd_sc_hd__a21o_1 _09612_ (.A1(_02604_),
    .A2(_02606_),
    .B1(_02760_),
    .X(_02762_));
 sky130_fd_sc_hd__and3_1 _09613_ (.A(_02604_),
    .B(_02606_),
    .C(_02760_),
    .X(_02763_));
 sky130_fd_sc_hd__nor2_2 _09614_ (.A(_02761_),
    .B(_02763_),
    .Y(_02764_));
 sky130_fd_sc_hd__a21boi_2 _09615_ (.A1(_02609_),
    .A2(_02613_),
    .B1_N(_02608_),
    .Y(_02765_));
 sky130_fd_sc_hd__xnor2_4 _09616_ (.A(_02764_),
    .B(_02765_),
    .Y(_02766_));
 sky130_fd_sc_hd__nand3b_1 _09617_ (.A_N(_02135_),
    .B(_02437_),
    .C(_02614_),
    .Y(_02767_));
 sky130_fd_sc_hd__or2_1 _09618_ (.A(_02212_),
    .B(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__a21oi_1 _09619_ (.A1(net21),
    .A2(_02768_),
    .B1(_02766_),
    .Y(_02769_));
 sky130_fd_sc_hd__a311oi_1 _09620_ (.A1(net21),
    .A2(_02766_),
    .A3(_02768_),
    .B1(_02769_),
    .C1(_02214_),
    .Y(_02770_));
 sky130_fd_sc_hd__or3_1 _09621_ (.A(net86),
    .B(_02166_),
    .C(_02168_),
    .X(_02771_));
 sky130_fd_sc_hd__o21ai_1 _09622_ (.A1(net86),
    .A2(_02168_),
    .B1(_02166_),
    .Y(_02772_));
 sky130_fd_sc_hd__mux2_1 _09623_ (.A0(_02447_),
    .A1(_02450_),
    .S(net230),
    .X(_02773_));
 sky130_fd_sc_hd__mux2_1 _09624_ (.A0(_02449_),
    .A1(_02457_),
    .S(net230),
    .X(_02774_));
 sky130_fd_sc_hd__mux2_1 _09625_ (.A0(_02773_),
    .A1(_02774_),
    .S(net231),
    .X(_02775_));
 sky130_fd_sc_hd__mux2_1 _09626_ (.A0(_02453_),
    .A1(_02465_),
    .S(net230),
    .X(_02776_));
 sky130_fd_sc_hd__mux2_1 _09627_ (.A0(_02454_),
    .A1(_02456_),
    .S(net228),
    .X(_02777_));
 sky130_fd_sc_hd__mux2_1 _09628_ (.A0(_02777_),
    .A1(_02776_),
    .S(net231),
    .X(_02778_));
 sky130_fd_sc_hd__mux2_1 _09629_ (.A0(_02775_),
    .A1(_02778_),
    .S(net235),
    .X(_02779_));
 sky130_fd_sc_hd__mux2_1 _09630_ (.A0(_02461_),
    .A1(_02471_),
    .S(net230),
    .X(_02780_));
 sky130_fd_sc_hd__mux2_1 _09631_ (.A0(_02462_),
    .A1(_02464_),
    .S(net228),
    .X(_02781_));
 sky130_fd_sc_hd__mux2_1 _09632_ (.A0(_02781_),
    .A1(_02780_),
    .S(net231),
    .X(_02782_));
 sky130_fd_sc_hd__mux2_1 _09633_ (.A0(_02468_),
    .A1(_02470_),
    .S(net228),
    .X(_02783_));
 sky130_fd_sc_hd__nor2_1 _09634_ (.A(net233),
    .B(_02783_),
    .Y(_02784_));
 sky130_fd_sc_hd__a21oi_1 _09635_ (.A1(net231),
    .A2(_02315_),
    .B1(_02784_),
    .Y(_02785_));
 sky130_fd_sc_hd__mux2_1 _09636_ (.A0(_02782_),
    .A1(_02785_),
    .S(net235),
    .X(_02786_));
 sky130_fd_sc_hd__mux2_2 _09637_ (.A0(_02779_),
    .A1(_02786_),
    .S(net238),
    .X(_02787_));
 sky130_fd_sc_hd__o21a_1 _09638_ (.A1(_02640_),
    .A2(_02641_),
    .B1(_02642_),
    .X(_02788_));
 sky130_fd_sc_hd__nor2_1 _09639_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .Y(_02789_));
 sky130_fd_sc_hd__or2_1 _09640_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .X(_02790_));
 sky130_fd_sc_hd__nand2_1 _09641_ (.A(reg1_val[3]),
    .B(curr_PC[3]),
    .Y(_02791_));
 sky130_fd_sc_hd__a21oi_1 _09642_ (.A1(_02790_),
    .A2(_02791_),
    .B1(_02788_),
    .Y(_02792_));
 sky130_fd_sc_hd__a31o_1 _09643_ (.A1(_02788_),
    .A2(_02790_),
    .A3(_02791_),
    .B1(net241),
    .X(_02793_));
 sky130_fd_sc_hd__o31a_1 _09644_ (.A1(\div_res[2] ),
    .A2(\div_res[1] ),
    .A3(\div_res[0] ),
    .B1(net26),
    .X(_02794_));
 sky130_fd_sc_hd__xor2_1 _09645_ (.A(\div_res[3] ),
    .B(_02794_),
    .X(_02795_));
 sky130_fd_sc_hd__o31a_1 _09646_ (.A1(\div_shifter[34] ),
    .A2(\div_shifter[33] ),
    .A3(\div_shifter[32] ),
    .B1(net246),
    .X(_02796_));
 sky130_fd_sc_hd__nor2_1 _09647_ (.A(\div_shifter[35] ),
    .B(_02796_),
    .Y(_02797_));
 sky130_fd_sc_hd__and2_1 _09648_ (.A(\div_shifter[35] ),
    .B(_02796_),
    .X(_02798_));
 sky130_fd_sc_hd__a21o_1 _09649_ (.A1(reg1_val[2]),
    .A2(_06293_),
    .B1(_02645_),
    .X(_02799_));
 sky130_fd_sc_hd__o21ai_1 _09650_ (.A1(reg1_val[2]),
    .A2(net233),
    .B1(_02799_),
    .Y(_02800_));
 sky130_fd_sc_hd__or3_1 _09651_ (.A(net300),
    .B(_06294_),
    .C(_06311_),
    .X(_02801_));
 sky130_fd_sc_hd__o21a_1 _09652_ (.A1(instruction[7]),
    .A2(_02800_),
    .B1(_02801_),
    .X(_02802_));
 sky130_fd_sc_hd__o21ai_1 _09653_ (.A1(_06291_),
    .A2(_02802_),
    .B1(net251),
    .Y(_02803_));
 sky130_fd_sc_hd__a21oi_1 _09654_ (.A1(_06291_),
    .A2(_02802_),
    .B1(_02803_),
    .Y(_02804_));
 sky130_fd_sc_hd__o21a_1 _09655_ (.A1(net233),
    .A2(_02272_),
    .B1(_02316_),
    .X(_02805_));
 sky130_fd_sc_hd__o21a_1 _09656_ (.A1(net234),
    .A2(_02805_),
    .B1(_02318_),
    .X(_02806_));
 sky130_fd_sc_hd__o21ai_2 _09657_ (.A1(net238),
    .A2(_02806_),
    .B1(_02312_),
    .Y(_02807_));
 sky130_fd_sc_hd__inv_2 _09658_ (.A(_02807_),
    .Y(_02808_));
 sky130_fd_sc_hd__nand2_1 _09659_ (.A(net305),
    .B(_02807_),
    .Y(_02809_));
 sky130_fd_sc_hd__o211a_1 _09660_ (.A1(net305),
    .A2(_02787_),
    .B1(_02809_),
    .C1(_06416_),
    .X(_02810_));
 sky130_fd_sc_hd__o221a_1 _09661_ (.A1(net263),
    .A2(_02787_),
    .B1(_02792_),
    .B2(_02793_),
    .C1(_06412_),
    .X(_02811_));
 sky130_fd_sc_hd__o32a_1 _09662_ (.A1(net249),
    .A2(_02797_),
    .A3(_02798_),
    .B1(net204),
    .B2(_06290_),
    .X(_02812_));
 sky130_fd_sc_hd__o221a_1 _09663_ (.A1(_06289_),
    .A2(_02291_),
    .B1(_02295_),
    .B2(_06291_),
    .C1(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__or3b_1 _09664_ (.A(_02804_),
    .B(_02811_),
    .C_N(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__a211o_1 _09665_ (.A1(_02305_),
    .A2(_02795_),
    .B1(_02810_),
    .C1(_02814_),
    .X(_02815_));
 sky130_fd_sc_hd__a31o_1 _09666_ (.A1(_02298_),
    .A2(_02771_),
    .A3(_02772_),
    .B1(_02815_),
    .X(_02816_));
 sky130_fd_sc_hd__a211o_2 _09667_ (.A1(net236),
    .A2(net212),
    .B1(_02770_),
    .C1(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__or2_1 _09668_ (.A(curr_PC[3]),
    .B(_02664_),
    .X(_02818_));
 sky130_fd_sc_hd__and2_1 _09669_ (.A(curr_PC[3]),
    .B(_02664_),
    .X(_02819_));
 sky130_fd_sc_hd__nor2_1 _09670_ (.A(net257),
    .B(_02819_),
    .Y(_02820_));
 sky130_fd_sc_hd__a22o_4 _09671_ (.A1(net257),
    .A2(_02817_),
    .B1(_02818_),
    .B2(_02820_),
    .X(dest_val[3]));
 sky130_fd_sc_hd__a21o_1 _09672_ (.A1(_02666_),
    .A2(_02759_),
    .B1(_02758_),
    .X(_02821_));
 sky130_fd_sc_hd__a21bo_1 _09673_ (.A1(_02748_),
    .A2(_02754_),
    .B1_N(_02756_),
    .X(_02822_));
 sky130_fd_sc_hd__a21o_1 _09674_ (.A1(_02700_),
    .A2(_02716_),
    .B1(_02715_),
    .X(_02823_));
 sky130_fd_sc_hd__o22a_1 _09675_ (.A1(net147),
    .A2(net12),
    .B1(net45),
    .B2(net144),
    .X(_02824_));
 sky130_fd_sc_hd__xnor2_1 _09676_ (.A(net97),
    .B(_02824_),
    .Y(_02825_));
 sky130_fd_sc_hd__inv_2 _09677_ (.A(_02825_),
    .Y(_02826_));
 sky130_fd_sc_hd__a2bb2o_1 _09678_ (.A1_N(_00306_),
    .A2_N(net88),
    .B1(_00430_),
    .B2(_00308_),
    .X(_02827_));
 sky130_fd_sc_hd__xor2_1 _09679_ (.A(net109),
    .B(_02827_),
    .X(_02828_));
 sky130_fd_sc_hd__xor2_1 _09680_ (.A(_02825_),
    .B(_02828_),
    .X(_02829_));
 sky130_fd_sc_hd__o22a_1 _09681_ (.A1(net14),
    .A2(net133),
    .B1(net90),
    .B2(net52),
    .X(_02830_));
 sky130_fd_sc_hd__xnor2_1 _09682_ (.A(net112),
    .B(_02830_),
    .Y(_02831_));
 sky130_fd_sc_hd__and2b_1 _09683_ (.A_N(_02829_),
    .B(_02831_),
    .X(_02832_));
 sky130_fd_sc_hd__and2b_1 _09684_ (.A_N(_02831_),
    .B(_02829_),
    .X(_02833_));
 sky130_fd_sc_hd__or2_2 _09685_ (.A(_02832_),
    .B(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__a21oi_2 _09686_ (.A1(_02683_),
    .A2(_02687_),
    .B1(_02686_),
    .Y(_02835_));
 sky130_fd_sc_hd__xnor2_1 _09687_ (.A(_02834_),
    .B(_02835_),
    .Y(_02836_));
 sky130_fd_sc_hd__nand2b_1 _09688_ (.A_N(_02836_),
    .B(_02823_),
    .Y(_02837_));
 sky130_fd_sc_hd__xnor2_1 _09689_ (.A(_02823_),
    .B(_02836_),
    .Y(_02838_));
 sky130_fd_sc_hd__o21ai_2 _09690_ (.A1(_02706_),
    .A2(_02708_),
    .B1(_02705_),
    .Y(_02839_));
 sky130_fd_sc_hd__a21oi_1 _09691_ (.A1(_02734_),
    .A2(_02736_),
    .B1(_02733_),
    .Y(_02840_));
 sky130_fd_sc_hd__o21ba_1 _09692_ (.A1(_02690_),
    .A2(_02698_),
    .B1_N(_02697_),
    .X(_02841_));
 sky130_fd_sc_hd__nor2_1 _09693_ (.A(_02840_),
    .B(_02841_),
    .Y(_02842_));
 sky130_fd_sc_hd__and2_1 _09694_ (.A(_02840_),
    .B(_02841_),
    .X(_02843_));
 sky130_fd_sc_hd__or2_1 _09695_ (.A(_02842_),
    .B(_02843_),
    .X(_02844_));
 sky130_fd_sc_hd__and2b_1 _09696_ (.A_N(_02844_),
    .B(_02839_),
    .X(_02845_));
 sky130_fd_sc_hd__xnor2_2 _09697_ (.A(_02839_),
    .B(_02844_),
    .Y(_02846_));
 sky130_fd_sc_hd__nor2_2 _09698_ (.A(net149),
    .B(net31),
    .Y(_02847_));
 sky130_fd_sc_hd__o21a_2 _09699_ (.A1(_00180_),
    .A2(_02713_),
    .B1(_02712_),
    .X(_02848_));
 sky130_fd_sc_hd__o22a_2 _09700_ (.A1(net141),
    .A2(net8),
    .B1(net6),
    .B2(net143),
    .X(_02849_));
 sky130_fd_sc_hd__xnor2_4 _09701_ (.A(net31),
    .B(_02849_),
    .Y(_02850_));
 sky130_fd_sc_hd__nor2_1 _09702_ (.A(_02848_),
    .B(_02850_),
    .Y(_02851_));
 sky130_fd_sc_hd__xor2_4 _09703_ (.A(_02848_),
    .B(_02850_),
    .X(_02852_));
 sky130_fd_sc_hd__xnor2_2 _09704_ (.A(_02847_),
    .B(_02852_),
    .Y(_02853_));
 sky130_fd_sc_hd__o22a_1 _09705_ (.A1(net114),
    .A2(net63),
    .B1(net55),
    .B2(net116),
    .X(_02854_));
 sky130_fd_sc_hd__xnor2_2 _09706_ (.A(net179),
    .B(_02854_),
    .Y(_02855_));
 sky130_fd_sc_hd__a32o_1 _09707_ (.A1(_00138_),
    .A2(_00219_),
    .A3(_00221_),
    .B1(_00197_),
    .B2(_06498_),
    .X(_02856_));
 sky130_fd_sc_hd__xnor2_1 _09708_ (.A(_06490_),
    .B(_02856_),
    .Y(_02857_));
 sky130_fd_sc_hd__o22a_1 _09709_ (.A1(net83),
    .A2(net65),
    .B1(net58),
    .B2(net130),
    .X(_02858_));
 sky130_fd_sc_hd__xnor2_1 _09710_ (.A(net157),
    .B(_02858_),
    .Y(_02859_));
 sky130_fd_sc_hd__or2_1 _09711_ (.A(_02857_),
    .B(_02859_),
    .X(_02860_));
 sky130_fd_sc_hd__nand2_1 _09712_ (.A(_02857_),
    .B(_02859_),
    .Y(_02861_));
 sky130_fd_sc_hd__nand2_1 _09713_ (.A(_02860_),
    .B(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__xor2_2 _09714_ (.A(_02855_),
    .B(_02862_),
    .X(_02863_));
 sky130_fd_sc_hd__o22a_1 _09715_ (.A1(net78),
    .A2(net74),
    .B1(net68),
    .B2(net123),
    .X(_02864_));
 sky130_fd_sc_hd__xnor2_1 _09716_ (.A(net154),
    .B(_02864_),
    .Y(_02865_));
 sky130_fd_sc_hd__o22a_1 _09717_ (.A1(net99),
    .A2(net36),
    .B1(net34),
    .B2(net119),
    .X(_02866_));
 sky130_fd_sc_hd__xnor2_1 _09718_ (.A(net135),
    .B(_02866_),
    .Y(_02867_));
 sky130_fd_sc_hd__nand2_1 _09719_ (.A(_02865_),
    .B(_02867_),
    .Y(_02868_));
 sky130_fd_sc_hd__xor2_1 _09720_ (.A(_02865_),
    .B(_02867_),
    .X(_02869_));
 sky130_fd_sc_hd__o22a_1 _09721_ (.A1(net71),
    .A2(net42),
    .B1(net94),
    .B2(net77),
    .X(_02870_));
 sky130_fd_sc_hd__xnor2_1 _09722_ (.A(net138),
    .B(_02870_),
    .Y(_02871_));
 sky130_fd_sc_hd__nand2_1 _09723_ (.A(_02869_),
    .B(_02871_),
    .Y(_02872_));
 sky130_fd_sc_hd__xor2_1 _09724_ (.A(_02869_),
    .B(_02871_),
    .X(_02873_));
 sky130_fd_sc_hd__o22a_1 _09725_ (.A1(net177),
    .A2(net17),
    .B1(net10),
    .B2(net175),
    .X(_02874_));
 sky130_fd_sc_hd__xor2_1 _09726_ (.A(net189),
    .B(_02874_),
    .X(_02875_));
 sky130_fd_sc_hd__nor2_1 _09727_ (.A(net169),
    .B(net3),
    .Y(_02876_));
 sky130_fd_sc_hd__xnor2_1 _09728_ (.A(net210),
    .B(_02876_),
    .Y(_02877_));
 sky130_fd_sc_hd__nor2_1 _09729_ (.A(_02875_),
    .B(_02877_),
    .Y(_02878_));
 sky130_fd_sc_hd__xnor2_1 _09730_ (.A(_02875_),
    .B(_02877_),
    .Y(_02879_));
 sky130_fd_sc_hd__and2_1 _09731_ (.A(_02873_),
    .B(_02879_),
    .X(_02880_));
 sky130_fd_sc_hd__nor2_1 _09732_ (.A(_02873_),
    .B(_02879_),
    .Y(_02881_));
 sky130_fd_sc_hd__nor2_1 _09733_ (.A(_02880_),
    .B(_02881_),
    .Y(_02882_));
 sky130_fd_sc_hd__xnor2_2 _09734_ (.A(_02863_),
    .B(_02882_),
    .Y(_02883_));
 sky130_fd_sc_hd__nor2_1 _09735_ (.A(_02853_),
    .B(_02883_),
    .Y(_02884_));
 sky130_fd_sc_hd__xor2_2 _09736_ (.A(_02853_),
    .B(_02883_),
    .X(_02885_));
 sky130_fd_sc_hd__xnor2_1 _09737_ (.A(_02846_),
    .B(_02885_),
    .Y(_02886_));
 sky130_fd_sc_hd__a21o_1 _09738_ (.A1(_02670_),
    .A2(_02672_),
    .B1(_02676_),
    .X(_02887_));
 sky130_fd_sc_hd__o22a_1 _09739_ (.A1(net126),
    .A2(net50),
    .B1(net48),
    .B2(net121),
    .X(_02888_));
 sky130_fd_sc_hd__xnor2_1 _09740_ (.A(net106),
    .B(_02888_),
    .Y(_02889_));
 sky130_fd_sc_hd__o22a_1 _09741_ (.A1(net80),
    .A2(net40),
    .B1(net38),
    .B2(net128),
    .X(_02890_));
 sky130_fd_sc_hd__xnor2_1 _09742_ (.A(net102),
    .B(_02890_),
    .Y(_02891_));
 sky130_fd_sc_hd__nand2_1 _09743_ (.A(_02889_),
    .B(_02891_),
    .Y(_02892_));
 sky130_fd_sc_hd__or2_1 _09744_ (.A(_02889_),
    .B(_02891_),
    .X(_02893_));
 sky130_fd_sc_hd__nand2_1 _09745_ (.A(_02892_),
    .B(_02893_),
    .Y(_02894_));
 sky130_fd_sc_hd__a21oi_2 _09746_ (.A1(_02718_),
    .A2(_02723_),
    .B1(_02722_),
    .Y(_02895_));
 sky130_fd_sc_hd__nor2_1 _09747_ (.A(_02894_),
    .B(_02895_),
    .Y(_02896_));
 sky130_fd_sc_hd__xor2_2 _09748_ (.A(_02894_),
    .B(_02895_),
    .X(_02897_));
 sky130_fd_sc_hd__xnor2_1 _09749_ (.A(_02887_),
    .B(_02897_),
    .Y(_02898_));
 sky130_fd_sc_hd__nor2_1 _09750_ (.A(_02886_),
    .B(_02898_),
    .Y(_02899_));
 sky130_fd_sc_hd__nand2_1 _09751_ (.A(_02886_),
    .B(_02898_),
    .Y(_02900_));
 sky130_fd_sc_hd__and2b_1 _09752_ (.A_N(_02899_),
    .B(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__xor2_1 _09753_ (.A(_02838_),
    .B(_02901_),
    .X(_02902_));
 sky130_fd_sc_hd__a21o_1 _09754_ (.A1(_02682_),
    .A2(_02745_),
    .B1(_02743_),
    .X(_02903_));
 sky130_fd_sc_hd__o21ai_4 _09755_ (.A1(_02678_),
    .A2(_02679_),
    .B1(_02681_),
    .Y(_02904_));
 sky130_fd_sc_hd__a21o_2 _09756_ (.A1(_02688_),
    .A2(_02726_),
    .B1(_02725_),
    .X(_02905_));
 sky130_fd_sc_hd__nor2_2 _09757_ (.A(_02739_),
    .B(_02741_),
    .Y(_02906_));
 sky130_fd_sc_hd__o21ai_1 _09758_ (.A1(_02739_),
    .A2(_02741_),
    .B1(_02905_),
    .Y(_02907_));
 sky130_fd_sc_hd__xnor2_4 _09759_ (.A(_02905_),
    .B(_02906_),
    .Y(_02908_));
 sky130_fd_sc_hd__xnor2_2 _09760_ (.A(_02904_),
    .B(_02908_),
    .Y(_02909_));
 sky130_fd_sc_hd__a21oi_2 _09761_ (.A1(_02749_),
    .A2(_02753_),
    .B1(_02752_),
    .Y(_02910_));
 sky130_fd_sc_hd__xnor2_1 _09762_ (.A(_02909_),
    .B(_02910_),
    .Y(_02911_));
 sky130_fd_sc_hd__nand2b_1 _09763_ (.A_N(_02911_),
    .B(_02903_),
    .Y(_02912_));
 sky130_fd_sc_hd__xnor2_1 _09764_ (.A(_02903_),
    .B(_02911_),
    .Y(_02913_));
 sky130_fd_sc_hd__and2_1 _09765_ (.A(_02902_),
    .B(_02913_),
    .X(_02914_));
 sky130_fd_sc_hd__xor2_1 _09766_ (.A(_02902_),
    .B(_02913_),
    .X(_02915_));
 sky130_fd_sc_hd__xor2_1 _09767_ (.A(_02822_),
    .B(_02915_),
    .X(_02916_));
 sky130_fd_sc_hd__and2_1 _09768_ (.A(_02821_),
    .B(_02916_),
    .X(_02917_));
 sky130_fd_sc_hd__nor2_1 _09769_ (.A(_02821_),
    .B(_02916_),
    .Y(_02918_));
 sky130_fd_sc_hd__nor2_2 _09770_ (.A(_02917_),
    .B(_02918_),
    .Y(_02919_));
 sky130_fd_sc_hd__and3b_1 _09771_ (.A_N(_02763_),
    .B(_02609_),
    .C(_02762_),
    .X(_02920_));
 sky130_fd_sc_hd__a21oi_1 _09772_ (.A1(_02608_),
    .A2(_02762_),
    .B1(_02763_),
    .Y(_02921_));
 sky130_fd_sc_hd__a21oi_1 _09773_ (.A1(_02611_),
    .A2(_02920_),
    .B1(_02921_),
    .Y(_02922_));
 sky130_fd_sc_hd__nand2_2 _09774_ (.A(_02612_),
    .B(_02920_),
    .Y(_02923_));
 sky130_fd_sc_hd__inv_2 _09775_ (.A(_02923_),
    .Y(_02924_));
 sky130_fd_sc_hd__a21bo_2 _09776_ (.A1(_02035_),
    .A2(_02924_),
    .B1_N(_02922_),
    .X(_02925_));
 sky130_fd_sc_hd__xor2_4 _09777_ (.A(_02919_),
    .B(_02925_),
    .X(_02926_));
 sky130_fd_sc_hd__o21a_1 _09778_ (.A1(_02766_),
    .A2(_02768_),
    .B1(net21),
    .X(_02927_));
 sky130_fd_sc_hd__o21ai_1 _09779_ (.A1(_02926_),
    .A2(_02927_),
    .B1(net206),
    .Y(_02928_));
 sky130_fd_sc_hd__a21oi_1 _09780_ (.A1(_02926_),
    .A2(_02927_),
    .B1(_02928_),
    .Y(_02929_));
 sky130_fd_sc_hd__and2_1 _09781_ (.A(net21),
    .B(_02169_),
    .X(_02930_));
 sky130_fd_sc_hd__a21oi_1 _09782_ (.A1(_02164_),
    .A2(_02930_),
    .B1(net250),
    .Y(_02931_));
 sky130_fd_sc_hd__o21a_1 _09783_ (.A1(_02164_),
    .A2(_02930_),
    .B1(_02931_),
    .X(_02932_));
 sky130_fd_sc_hd__o21a_1 _09784_ (.A1(_06289_),
    .A2(_02800_),
    .B1(_06290_),
    .X(_02933_));
 sky130_fd_sc_hd__or3_1 _09785_ (.A(net300),
    .B(_06288_),
    .C(_06312_),
    .X(_02934_));
 sky130_fd_sc_hd__o21a_1 _09786_ (.A1(net307),
    .A2(_02933_),
    .B1(_02934_),
    .X(_02935_));
 sky130_fd_sc_hd__a21oi_1 _09787_ (.A1(_06285_),
    .A2(_02935_),
    .B1(_02293_),
    .Y(_02936_));
 sky130_fd_sc_hd__o21a_1 _09788_ (.A1(_06285_),
    .A2(_02935_),
    .B1(_02936_),
    .X(_02937_));
 sky130_fd_sc_hd__mux2_1 _09789_ (.A0(_02232_),
    .A1(_02247_),
    .S(net232),
    .X(_02938_));
 sky130_fd_sc_hd__mux2_1 _09790_ (.A0(_02240_),
    .A1(_02263_),
    .S(net232),
    .X(_02939_));
 sky130_fd_sc_hd__mux2_1 _09791_ (.A0(_02938_),
    .A1(_02939_),
    .S(net234),
    .X(_02940_));
 sky130_fd_sc_hd__mux2_1 _09792_ (.A0(_02256_),
    .A1(_02279_),
    .S(net232),
    .X(_02941_));
 sky130_fd_sc_hd__mux2_1 _09793_ (.A0(_02941_),
    .A1(_02805_),
    .S(net234),
    .X(_02942_));
 sky130_fd_sc_hd__or2_1 _09794_ (.A(net239),
    .B(_02940_),
    .X(_02943_));
 sky130_fd_sc_hd__o21ai_2 _09795_ (.A1(net237),
    .A2(_02942_),
    .B1(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__nand2_1 _09796_ (.A(net241),
    .B(_02944_),
    .Y(_02945_));
 sky130_fd_sc_hd__o21a_1 _09797_ (.A1(_02788_),
    .A2(_02789_),
    .B1(_02791_),
    .X(_02946_));
 sky130_fd_sc_hd__nor2_1 _09798_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .Y(_02947_));
 sky130_fd_sc_hd__or2_1 _09799_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .X(_02948_));
 sky130_fd_sc_hd__nand2_1 _09800_ (.A(reg1_val[4]),
    .B(curr_PC[4]),
    .Y(_02949_));
 sky130_fd_sc_hd__and3_1 _09801_ (.A(_02946_),
    .B(_02948_),
    .C(_02949_),
    .X(_02950_));
 sky130_fd_sc_hd__a21oi_1 _09802_ (.A1(_02948_),
    .A2(_02949_),
    .B1(_02946_),
    .Y(_02951_));
 sky130_fd_sc_hd__o311a_1 _09803_ (.A1(net241),
    .A2(_02950_),
    .A3(_02951_),
    .B1(_06412_),
    .C1(_02945_),
    .X(_02952_));
 sky130_fd_sc_hd__or4_2 _09804_ (.A(\div_res[3] ),
    .B(\div_res[2] ),
    .C(\div_res[1] ),
    .D(\div_res[0] ),
    .X(_02953_));
 sky130_fd_sc_hd__and3_1 _09805_ (.A(\div_res[4] ),
    .B(net25),
    .C(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__a21oi_1 _09806_ (.A1(net25),
    .A2(_02953_),
    .B1(\div_res[4] ),
    .Y(_02955_));
 sky130_fd_sc_hd__or4_2 _09807_ (.A(\div_shifter[35] ),
    .B(\div_shifter[34] ),
    .C(\div_shifter[33] ),
    .D(\div_shifter[32] ),
    .X(_02956_));
 sky130_fd_sc_hd__and3_1 _09808_ (.A(\div_shifter[36] ),
    .B(net246),
    .C(_02956_),
    .X(_02957_));
 sky130_fd_sc_hd__a21oi_1 _09809_ (.A1(net246),
    .A2(_02956_),
    .B1(\div_shifter[36] ),
    .Y(_02958_));
 sky130_fd_sc_hd__or3_1 _09810_ (.A(net249),
    .B(_02957_),
    .C(_02958_),
    .X(_02959_));
 sky130_fd_sc_hd__o221a_1 _09811_ (.A1(_06281_),
    .A2(_06426_),
    .B1(_02301_),
    .B2(_06284_),
    .C1(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__o221a_1 _09812_ (.A1(_06283_),
    .A2(_02291_),
    .B1(_02295_),
    .B2(_06285_),
    .C1(_02960_),
    .X(_02961_));
 sky130_fd_sc_hd__o31a_1 _09813_ (.A1(net202),
    .A2(_02954_),
    .A3(_02955_),
    .B1(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__o21ai_1 _09814_ (.A1(net235),
    .A2(_02785_),
    .B1(_02318_),
    .Y(_02963_));
 sky130_fd_sc_hd__a21o_1 _09815_ (.A1(net237),
    .A2(_02963_),
    .B1(_02311_),
    .X(_02964_));
 sky130_fd_sc_hd__o221a_1 _09816_ (.A1(net182),
    .A2(_02944_),
    .B1(_02964_),
    .B2(net184),
    .C1(_02962_),
    .X(_02965_));
 sky130_fd_sc_hd__or4b_1 _09817_ (.A(_02932_),
    .B(_02937_),
    .C(_02952_),
    .D_N(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__o21a_1 _09818_ (.A1(_02929_),
    .A2(_02966_),
    .B1(net258),
    .X(_02967_));
 sky130_fd_sc_hd__nand2_1 _09819_ (.A(curr_PC[4]),
    .B(_02819_),
    .Y(_02968_));
 sky130_fd_sc_hd__or2_1 _09820_ (.A(curr_PC[4]),
    .B(_02819_),
    .X(_02969_));
 sky130_fd_sc_hd__a31o_4 _09821_ (.A1(net262),
    .A2(_02968_),
    .A3(_02969_),
    .B1(_02967_),
    .X(dest_val[4]));
 sky130_fd_sc_hd__a21o_1 _09822_ (.A1(_02822_),
    .A2(_02915_),
    .B1(_02914_),
    .X(_02970_));
 sky130_fd_sc_hd__o21ai_2 _09823_ (.A1(_02909_),
    .A2(_02910_),
    .B1(_02912_),
    .Y(_02971_));
 sky130_fd_sc_hd__a21o_1 _09824_ (.A1(_02863_),
    .A2(_02882_),
    .B1(_02880_),
    .X(_02972_));
 sky130_fd_sc_hd__o22a_1 _09825_ (.A1(net121),
    .A2(net51),
    .B1(net49),
    .B2(net80),
    .X(_02973_));
 sky130_fd_sc_hd__xnor2_1 _09826_ (.A(net106),
    .B(_02973_),
    .Y(_02974_));
 sky130_fd_sc_hd__o22a_1 _09827_ (.A1(net15),
    .A2(net90),
    .B1(net88),
    .B2(net52),
    .X(_02975_));
 sky130_fd_sc_hd__xnor2_1 _09828_ (.A(net112),
    .B(_02975_),
    .Y(_02976_));
 sky130_fd_sc_hd__and2_1 _09829_ (.A(_02974_),
    .B(_02976_),
    .X(_02977_));
 sky130_fd_sc_hd__nor2_1 _09830_ (.A(_02974_),
    .B(_02976_),
    .Y(_02978_));
 sky130_fd_sc_hd__nor2_1 _09831_ (.A(_02977_),
    .B(_02978_),
    .Y(_02979_));
 sky130_fd_sc_hd__a2bb2o_1 _09832_ (.A1_N(net125),
    .A2_N(net47),
    .B1(_00430_),
    .B2(_00307_),
    .X(_02980_));
 sky130_fd_sc_hd__xnor2_2 _09833_ (.A(net109),
    .B(_02980_),
    .Y(_02981_));
 sky130_fd_sc_hd__xnor2_1 _09834_ (.A(_02979_),
    .B(_02981_),
    .Y(_02982_));
 sky130_fd_sc_hd__o21a_1 _09835_ (.A1(_02842_),
    .A2(_02845_),
    .B1(_02982_),
    .X(_02983_));
 sky130_fd_sc_hd__nor3_1 _09836_ (.A(_02842_),
    .B(_02845_),
    .C(_02982_),
    .Y(_02984_));
 sky130_fd_sc_hd__nor2_1 _09837_ (.A(_02983_),
    .B(_02984_),
    .Y(_02985_));
 sky130_fd_sc_hd__xor2_2 _09838_ (.A(_02972_),
    .B(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__a21o_2 _09839_ (.A1(_02826_),
    .A2(_02828_),
    .B1(_02832_),
    .X(_02987_));
 sky130_fd_sc_hd__o22a_2 _09840_ (.A1(net77),
    .A2(net42),
    .B1(net94),
    .B2(net74),
    .X(_02988_));
 sky130_fd_sc_hd__xnor2_4 _09841_ (.A(net138),
    .B(_02988_),
    .Y(_02989_));
 sky130_fd_sc_hd__o22a_1 _09842_ (.A1(net128),
    .A2(net40),
    .B1(net38),
    .B2(net100),
    .X(_02990_));
 sky130_fd_sc_hd__xnor2_2 _09843_ (.A(net102),
    .B(_02990_),
    .Y(_02991_));
 sky130_fd_sc_hd__and2_1 _09844_ (.A(_02989_),
    .B(_02991_),
    .X(_02992_));
 sky130_fd_sc_hd__xor2_4 _09845_ (.A(_02989_),
    .B(_02991_),
    .X(_02993_));
 sky130_fd_sc_hd__o22a_2 _09846_ (.A1(net119),
    .A2(net36),
    .B1(net34),
    .B2(net71),
    .X(_02994_));
 sky130_fd_sc_hd__xnor2_4 _09847_ (.A(net135),
    .B(_02994_),
    .Y(_02995_));
 sky130_fd_sc_hd__xnor2_4 _09848_ (.A(_02993_),
    .B(_02995_),
    .Y(_02996_));
 sky130_fd_sc_hd__a21oi_4 _09849_ (.A1(_02847_),
    .A2(_02852_),
    .B1(_02851_),
    .Y(_02997_));
 sky130_fd_sc_hd__nor2_1 _09850_ (.A(_02996_),
    .B(_02997_),
    .Y(_02998_));
 sky130_fd_sc_hd__xor2_4 _09851_ (.A(_02996_),
    .B(_02997_),
    .X(_02999_));
 sky130_fd_sc_hd__xor2_2 _09852_ (.A(_02987_),
    .B(_02999_),
    .X(_03000_));
 sky130_fd_sc_hd__o21ai_2 _09853_ (.A1(_02855_),
    .A2(_02862_),
    .B1(_02860_),
    .Y(_03001_));
 sky130_fd_sc_hd__a21oi_1 _09854_ (.A1(_02868_),
    .A2(_02872_),
    .B1(_02878_),
    .Y(_03002_));
 sky130_fd_sc_hd__nand3_1 _09855_ (.A(_02868_),
    .B(_02872_),
    .C(_02878_),
    .Y(_03003_));
 sky130_fd_sc_hd__nand2b_1 _09856_ (.A_N(_03002_),
    .B(_03003_),
    .Y(_03004_));
 sky130_fd_sc_hd__xor2_2 _09857_ (.A(_03001_),
    .B(_03004_),
    .X(_03005_));
 sky130_fd_sc_hd__o22a_2 _09858_ (.A1(net177),
    .A2(net9),
    .B1(net3),
    .B2(_00168_),
    .X(_03006_));
 sky130_fd_sc_hd__xnor2_4 _09859_ (.A(net189),
    .B(_03006_),
    .Y(_03007_));
 sky130_fd_sc_hd__o22a_1 _09860_ (.A1(net152),
    .A2(_00223_),
    .B1(net17),
    .B2(net150),
    .X(_03008_));
 sky130_fd_sc_hd__xnor2_1 _09861_ (.A(net191),
    .B(_03008_),
    .Y(_03009_));
 sky130_fd_sc_hd__nand2b_2 _09862_ (.A_N(_03009_),
    .B(net210),
    .Y(_03010_));
 sky130_fd_sc_hd__nand2b_1 _09863_ (.A_N(net210),
    .B(_03009_),
    .Y(_03011_));
 sky130_fd_sc_hd__nand2_2 _09864_ (.A(_03010_),
    .B(_03011_),
    .Y(_03012_));
 sky130_fd_sc_hd__xor2_2 _09865_ (.A(_03007_),
    .B(_03012_),
    .X(_03013_));
 sky130_fd_sc_hd__o22a_1 _09866_ (.A1(net116),
    .A2(net63),
    .B1(net60),
    .B2(net114),
    .X(_03014_));
 sky130_fd_sc_hd__xnor2_1 _09867_ (.A(net179),
    .B(_03014_),
    .Y(_03015_));
 sky130_fd_sc_hd__o22a_1 _09868_ (.A1(net78),
    .A2(net68),
    .B1(net65),
    .B2(net123),
    .X(_03016_));
 sky130_fd_sc_hd__xor2_1 _09869_ (.A(net155),
    .B(_03016_),
    .X(_03017_));
 sky130_fd_sc_hd__nor2_1 _09870_ (.A(_03015_),
    .B(_03017_),
    .Y(_03018_));
 sky130_fd_sc_hd__xnor2_1 _09871_ (.A(_03015_),
    .B(_03017_),
    .Y(_03019_));
 sky130_fd_sc_hd__o22a_1 _09872_ (.A1(net83),
    .A2(net58),
    .B1(net55),
    .B2(net130),
    .X(_03020_));
 sky130_fd_sc_hd__xnor2_1 _09873_ (.A(net157),
    .B(_03020_),
    .Y(_03021_));
 sky130_fd_sc_hd__nor2_1 _09874_ (.A(_03019_),
    .B(_03021_),
    .Y(_03022_));
 sky130_fd_sc_hd__xnor2_1 _09875_ (.A(_03019_),
    .B(_03021_),
    .Y(_03023_));
 sky130_fd_sc_hd__nor2_1 _09876_ (.A(_02892_),
    .B(_03023_),
    .Y(_03024_));
 sky130_fd_sc_hd__nand2_1 _09877_ (.A(_02892_),
    .B(_03023_),
    .Y(_03025_));
 sky130_fd_sc_hd__and2b_1 _09878_ (.A_N(_03024_),
    .B(_03025_),
    .X(_03026_));
 sky130_fd_sc_hd__xnor2_1 _09879_ (.A(_03013_),
    .B(_03026_),
    .Y(_03027_));
 sky130_fd_sc_hd__o22a_1 _09880_ (.A1(net147),
    .A2(net8),
    .B1(net6),
    .B2(net141),
    .X(_03028_));
 sky130_fd_sc_hd__xnor2_1 _09881_ (.A(net31),
    .B(_03028_),
    .Y(_03029_));
 sky130_fd_sc_hd__o32a_1 _09882_ (.A1(net144),
    .A2(_00334_),
    .A3(_00335_),
    .B1(net45),
    .B2(net133),
    .X(_03030_));
 sky130_fd_sc_hd__xnor2_2 _09883_ (.A(net97),
    .B(_03030_),
    .Y(_03031_));
 sky130_fd_sc_hd__nor2_1 _09884_ (.A(net143),
    .B(net31),
    .Y(_03032_));
 sky130_fd_sc_hd__or3_1 _09885_ (.A(net143),
    .B(net31),
    .C(_03031_),
    .X(_03033_));
 sky130_fd_sc_hd__xnor2_1 _09886_ (.A(_03031_),
    .B(_03032_),
    .Y(_03034_));
 sky130_fd_sc_hd__nand2b_1 _09887_ (.A_N(_03029_),
    .B(_03034_),
    .Y(_03035_));
 sky130_fd_sc_hd__xor2_1 _09888_ (.A(_03029_),
    .B(_03034_),
    .X(_03036_));
 sky130_fd_sc_hd__or2_1 _09889_ (.A(_03027_),
    .B(_03036_),
    .X(_03037_));
 sky130_fd_sc_hd__and2_1 _09890_ (.A(_03027_),
    .B(_03036_),
    .X(_03038_));
 sky130_fd_sc_hd__nand2_1 _09891_ (.A(_03027_),
    .B(_03036_),
    .Y(_03039_));
 sky130_fd_sc_hd__nand2_1 _09892_ (.A(_03037_),
    .B(_03039_),
    .Y(_03040_));
 sky130_fd_sc_hd__xor2_2 _09893_ (.A(_03005_),
    .B(_03040_),
    .X(_03041_));
 sky130_fd_sc_hd__and2_1 _09894_ (.A(_03000_),
    .B(_03041_),
    .X(_03042_));
 sky130_fd_sc_hd__xor2_2 _09895_ (.A(_03000_),
    .B(_03041_),
    .X(_03043_));
 sky130_fd_sc_hd__xor2_2 _09896_ (.A(_02986_),
    .B(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__a21o_1 _09897_ (.A1(_02838_),
    .A2(_02900_),
    .B1(_02899_),
    .X(_03045_));
 sky130_fd_sc_hd__o21ai_4 _09898_ (.A1(_02834_),
    .A2(_02835_),
    .B1(_02837_),
    .Y(_03046_));
 sky130_fd_sc_hd__a21oi_4 _09899_ (.A1(_02846_),
    .A2(_02885_),
    .B1(_02884_),
    .Y(_03047_));
 sky130_fd_sc_hd__a21oi_4 _09900_ (.A1(_02887_),
    .A2(_02897_),
    .B1(_02896_),
    .Y(_03048_));
 sky130_fd_sc_hd__nor2_1 _09901_ (.A(_03047_),
    .B(_03048_),
    .Y(_03049_));
 sky130_fd_sc_hd__xor2_4 _09902_ (.A(_03047_),
    .B(_03048_),
    .X(_03050_));
 sky130_fd_sc_hd__xnor2_4 _09903_ (.A(_03046_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__a21boi_4 _09904_ (.A1(_02904_),
    .A2(_02908_),
    .B1_N(_02907_),
    .Y(_03052_));
 sky130_fd_sc_hd__xnor2_2 _09905_ (.A(_03051_),
    .B(_03052_),
    .Y(_03053_));
 sky130_fd_sc_hd__nand2b_1 _09906_ (.A_N(_03053_),
    .B(_03045_),
    .Y(_03054_));
 sky130_fd_sc_hd__xnor2_2 _09907_ (.A(_03045_),
    .B(_03053_),
    .Y(_03055_));
 sky130_fd_sc_hd__and2_1 _09908_ (.A(_03044_),
    .B(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__xor2_2 _09909_ (.A(_03044_),
    .B(_03055_),
    .X(_03057_));
 sky130_fd_sc_hd__xor2_1 _09910_ (.A(_02971_),
    .B(_03057_),
    .X(_03058_));
 sky130_fd_sc_hd__and2_1 _09911_ (.A(_02970_),
    .B(_03058_),
    .X(_03059_));
 sky130_fd_sc_hd__nor2_1 _09912_ (.A(_02970_),
    .B(_03058_),
    .Y(_03060_));
 sky130_fd_sc_hd__inv_2 _09913_ (.A(_03060_),
    .Y(_03061_));
 sky130_fd_sc_hd__nor2_2 _09914_ (.A(_03059_),
    .B(_03060_),
    .Y(_03062_));
 sky130_fd_sc_hd__a21oi_2 _09915_ (.A1(_02919_),
    .A2(_02925_),
    .B1(_02917_),
    .Y(_03063_));
 sky130_fd_sc_hd__xnor2_4 _09916_ (.A(_03062_),
    .B(_03063_),
    .Y(_03064_));
 sky130_fd_sc_hd__or3_1 _09917_ (.A(_02766_),
    .B(_02768_),
    .C(_02926_),
    .X(_03065_));
 sky130_fd_sc_hd__a21oi_1 _09918_ (.A1(net21),
    .A2(_03065_),
    .B1(_03064_),
    .Y(_03066_));
 sky130_fd_sc_hd__and3_1 _09919_ (.A(net21),
    .B(_03064_),
    .C(_03065_),
    .X(_03067_));
 sky130_fd_sc_hd__a21oi_1 _09920_ (.A1(net21),
    .A2(_02170_),
    .B1(_02162_),
    .Y(_03068_));
 sky130_fd_sc_hd__a31o_1 _09921_ (.A1(net21),
    .A2(_02162_),
    .A3(_02170_),
    .B1(net250),
    .X(_03069_));
 sky130_fd_sc_hd__or2_1 _09922_ (.A(_03068_),
    .B(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__o21ai_1 _09923_ (.A1(_06283_),
    .A2(_02933_),
    .B1(_06284_),
    .Y(_03071_));
 sky130_fd_sc_hd__or3_1 _09924_ (.A(net300),
    .B(_06282_),
    .C(_06313_),
    .X(_03072_));
 sky130_fd_sc_hd__a21bo_1 _09925_ (.A1(net300),
    .A2(_03071_),
    .B1_N(_03072_),
    .X(_03073_));
 sky130_fd_sc_hd__xnor2_1 _09926_ (.A(_06278_),
    .B(_03073_),
    .Y(_03074_));
 sky130_fd_sc_hd__o21a_1 _09927_ (.A1(_02946_),
    .A2(_02947_),
    .B1(_02949_),
    .X(_03075_));
 sky130_fd_sc_hd__nor2_1 _09928_ (.A(reg1_val[5]),
    .B(curr_PC[5]),
    .Y(_03076_));
 sky130_fd_sc_hd__nand2_1 _09929_ (.A(reg1_val[5]),
    .B(curr_PC[5]),
    .Y(_03077_));
 sky130_fd_sc_hd__and2b_1 _09930_ (.A_N(_03076_),
    .B(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__xnor2_1 _09931_ (.A(_03075_),
    .B(_03078_),
    .Y(_03079_));
 sky130_fd_sc_hd__mux2_1 _09932_ (.A0(_02451_),
    .A1(_02458_),
    .S(net231),
    .X(_03080_));
 sky130_fd_sc_hd__nand2b_1 _09933_ (.A_N(_02466_),
    .B(net231),
    .Y(_03081_));
 sky130_fd_sc_hd__o21ai_1 _09934_ (.A1(net231),
    .A2(_02455_),
    .B1(_03081_),
    .Y(_03082_));
 sky130_fd_sc_hd__nor2_1 _09935_ (.A(net236),
    .B(_03080_),
    .Y(_03083_));
 sky130_fd_sc_hd__a211o_1 _09936_ (.A1(net236),
    .A2(_03082_),
    .B1(_03083_),
    .C1(net238),
    .X(_03084_));
 sky130_fd_sc_hd__nand2b_1 _09937_ (.A_N(_02472_),
    .B(net231),
    .Y(_03085_));
 sky130_fd_sc_hd__o21ai_1 _09938_ (.A1(net231),
    .A2(_02463_),
    .B1(_03085_),
    .Y(_03086_));
 sky130_fd_sc_hd__mux2_1 _09939_ (.A0(_03086_),
    .A1(_02621_),
    .S(net235),
    .X(_03087_));
 sky130_fd_sc_hd__o21a_1 _09940_ (.A1(net237),
    .A2(_03087_),
    .B1(_03084_),
    .X(_03088_));
 sky130_fd_sc_hd__nor2_1 _09941_ (.A(net241),
    .B(_03079_),
    .Y(_03089_));
 sky130_fd_sc_hd__a211o_1 _09942_ (.A1(net242),
    .A2(_03088_),
    .B1(_03089_),
    .C1(net214),
    .X(_03090_));
 sky130_fd_sc_hd__o21ai_1 _09943_ (.A1(\div_res[4] ),
    .A2(_02953_),
    .B1(net25),
    .Y(_03091_));
 sky130_fd_sc_hd__xnor2_1 _09944_ (.A(\div_res[5] ),
    .B(_03091_),
    .Y(_03092_));
 sky130_fd_sc_hd__o21a_1 _09945_ (.A1(\div_shifter[36] ),
    .A2(_02956_),
    .B1(net246),
    .X(_03093_));
 sky130_fd_sc_hd__o21ai_1 _09946_ (.A1(\div_shifter[37] ),
    .A2(_03093_),
    .B1(_02303_),
    .Y(_03094_));
 sky130_fd_sc_hd__a21oi_1 _09947_ (.A1(\div_shifter[37] ),
    .A2(_03093_),
    .B1(_03094_),
    .Y(_03095_));
 sky130_fd_sc_hd__a221o_1 _09948_ (.A1(_06273_),
    .A2(net213),
    .B1(_02300_),
    .B2(_06277_),
    .C1(_03095_),
    .X(_03096_));
 sky130_fd_sc_hd__a221o_1 _09949_ (.A1(_06276_),
    .A2(net205),
    .B1(_02294_),
    .B2(_06278_),
    .C1(_03096_),
    .X(_03097_));
 sky130_fd_sc_hd__a21oi_1 _09950_ (.A1(_02305_),
    .A2(_03092_),
    .B1(_03097_),
    .Y(_03098_));
 sky130_fd_sc_hd__o21ai_1 _09951_ (.A1(net234),
    .A2(_02637_),
    .B1(_02318_),
    .Y(_03099_));
 sky130_fd_sc_hd__a21o_1 _09952_ (.A1(net237),
    .A2(_03099_),
    .B1(_02311_),
    .X(_03100_));
 sky130_fd_sc_hd__o221a_1 _09953_ (.A1(net183),
    .A2(_03088_),
    .B1(_03100_),
    .B2(net186),
    .C1(_03098_),
    .X(_03101_));
 sky130_fd_sc_hd__o211a_1 _09954_ (.A1(_02293_),
    .A2(_03074_),
    .B1(_03090_),
    .C1(_03101_),
    .X(_03102_));
 sky130_fd_sc_hd__o311a_2 _09955_ (.A1(_02214_),
    .A2(_03066_),
    .A3(_03067_),
    .B1(_03070_),
    .C1(_03102_),
    .X(_03103_));
 sky130_fd_sc_hd__a21oi_1 _09956_ (.A1(curr_PC[4]),
    .A2(_02819_),
    .B1(curr_PC[5]),
    .Y(_03104_));
 sky130_fd_sc_hd__and3_1 _09957_ (.A(curr_PC[4]),
    .B(curr_PC[5]),
    .C(_02819_),
    .X(_03105_));
 sky130_fd_sc_hd__or3_1 _09958_ (.A(net257),
    .B(_03104_),
    .C(_03105_),
    .X(_03106_));
 sky130_fd_sc_hd__o21ai_4 _09959_ (.A1(net262),
    .A2(_03103_),
    .B1(_03106_),
    .Y(dest_val[5]));
 sky130_fd_sc_hd__a21oi_4 _09960_ (.A1(_02971_),
    .A2(_03057_),
    .B1(_03056_),
    .Y(_03107_));
 sky130_fd_sc_hd__o21ai_4 _09961_ (.A1(_03051_),
    .A2(_03052_),
    .B1(_03054_),
    .Y(_03108_));
 sky130_fd_sc_hd__a21oi_2 _09962_ (.A1(_03013_),
    .A2(_03025_),
    .B1(_03024_),
    .Y(_03109_));
 sky130_fd_sc_hd__o22a_1 _09963_ (.A1(net126),
    .A2(net13),
    .B1(_00309_),
    .B2(net121),
    .X(_03110_));
 sky130_fd_sc_hd__xnor2_1 _09964_ (.A(net109),
    .B(_03110_),
    .Y(_03111_));
 sky130_fd_sc_hd__o22a_1 _09965_ (.A1(net100),
    .A2(net40),
    .B1(net38),
    .B2(net119),
    .X(_03112_));
 sky130_fd_sc_hd__xnor2_1 _09966_ (.A(net102),
    .B(_03112_),
    .Y(_03113_));
 sky130_fd_sc_hd__and2_1 _09967_ (.A(_03111_),
    .B(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__nor2_1 _09968_ (.A(_03111_),
    .B(_03113_),
    .Y(_03115_));
 sky130_fd_sc_hd__nor2_2 _09969_ (.A(_03114_),
    .B(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__o22a_1 _09970_ (.A1(net80),
    .A2(net50),
    .B1(net49),
    .B2(net128),
    .X(_03117_));
 sky130_fd_sc_hd__xnor2_2 _09971_ (.A(net106),
    .B(_03117_),
    .Y(_03118_));
 sky130_fd_sc_hd__xor2_4 _09972_ (.A(_03116_),
    .B(_03118_),
    .X(_03119_));
 sky130_fd_sc_hd__a21o_2 _09973_ (.A1(_03001_),
    .A2(_03003_),
    .B1(_03002_),
    .X(_03120_));
 sky130_fd_sc_hd__xor2_4 _09974_ (.A(_03119_),
    .B(_03120_),
    .X(_03121_));
 sky130_fd_sc_hd__nand2b_1 _09975_ (.A_N(_03109_),
    .B(_03121_),
    .Y(_03122_));
 sky130_fd_sc_hd__xnor2_4 _09976_ (.A(_03109_),
    .B(_03121_),
    .Y(_03123_));
 sky130_fd_sc_hd__o21bai_2 _09977_ (.A1(_02978_),
    .A2(_02981_),
    .B1_N(_02977_),
    .Y(_03124_));
 sky130_fd_sc_hd__o22a_1 _09978_ (.A1(net74),
    .A2(net42),
    .B1(net94),
    .B2(net68),
    .X(_03125_));
 sky130_fd_sc_hd__xnor2_1 _09979_ (.A(net138),
    .B(_03125_),
    .Y(_03126_));
 sky130_fd_sc_hd__o22a_1 _09980_ (.A1(net71),
    .A2(net36),
    .B1(net34),
    .B2(net76),
    .X(_03127_));
 sky130_fd_sc_hd__xnor2_1 _09981_ (.A(net135),
    .B(_03127_),
    .Y(_03128_));
 sky130_fd_sc_hd__and2_1 _09982_ (.A(_03126_),
    .B(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__nor2_1 _09983_ (.A(_03126_),
    .B(_03128_),
    .Y(_03130_));
 sky130_fd_sc_hd__or2_1 _09984_ (.A(_03129_),
    .B(_03130_),
    .X(_03131_));
 sky130_fd_sc_hd__a21o_1 _09985_ (.A1(_03033_),
    .A2(_03035_),
    .B1(_03131_),
    .X(_03132_));
 sky130_fd_sc_hd__nand3_1 _09986_ (.A(_03033_),
    .B(_03035_),
    .C(_03131_),
    .Y(_03133_));
 sky130_fd_sc_hd__and2_1 _09987_ (.A(_03132_),
    .B(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__nand2_1 _09988_ (.A(_03124_),
    .B(_03134_),
    .Y(_03135_));
 sky130_fd_sc_hd__xnor2_1 _09989_ (.A(_03124_),
    .B(_03134_),
    .Y(_03136_));
 sky130_fd_sc_hd__o21ai_4 _09990_ (.A1(_03007_),
    .A2(_03012_),
    .B1(_03010_),
    .Y(_03137_));
 sky130_fd_sc_hd__o211a_1 _09991_ (.A1(_03018_),
    .A2(_03022_),
    .B1(_00310_),
    .C1(net33),
    .X(_03138_));
 sky130_fd_sc_hd__a211o_1 _09992_ (.A1(_00310_),
    .A2(net33),
    .B1(_03018_),
    .C1(_03022_),
    .X(_03139_));
 sky130_fd_sc_hd__and2b_1 _09993_ (.A_N(_03138_),
    .B(_03139_),
    .X(_03140_));
 sky130_fd_sc_hd__xor2_2 _09994_ (.A(_03137_),
    .B(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__a32o_1 _09995_ (.A1(_00153_),
    .A2(_00219_),
    .A3(_00221_),
    .B1(_00197_),
    .B2(_00151_),
    .X(_03142_));
 sky130_fd_sc_hd__xor2_4 _09996_ (.A(net179),
    .B(_03142_),
    .X(_03143_));
 sky130_fd_sc_hd__o22a_2 _09997_ (.A1(net78),
    .A2(net64),
    .B1(net58),
    .B2(net123),
    .X(_03144_));
 sky130_fd_sc_hd__xor2_4 _09998_ (.A(net155),
    .B(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__nor2_1 _09999_ (.A(_03143_),
    .B(_03145_),
    .Y(_03146_));
 sky130_fd_sc_hd__xor2_4 _10000_ (.A(_03143_),
    .B(_03145_),
    .X(_03147_));
 sky130_fd_sc_hd__o22a_2 _10001_ (.A1(net130),
    .A2(net63),
    .B1(net55),
    .B2(net83),
    .X(_03148_));
 sky130_fd_sc_hd__xnor2_4 _10002_ (.A(_06435_),
    .B(_03148_),
    .Y(_03149_));
 sky130_fd_sc_hd__xnor2_4 _10003_ (.A(_03147_),
    .B(_03149_),
    .Y(_03150_));
 sky130_fd_sc_hd__a21oi_4 _10004_ (.A1(_02993_),
    .A2(_02995_),
    .B1(_02992_),
    .Y(_03151_));
 sky130_fd_sc_hd__nor2_1 _10005_ (.A(_03150_),
    .B(_03151_),
    .Y(_03152_));
 sky130_fd_sc_hd__xnor2_4 _10006_ (.A(_03150_),
    .B(_03151_),
    .Y(_03153_));
 sky130_fd_sc_hd__o22a_1 _10007_ (.A1(net152),
    .A2(net17),
    .B1(net9),
    .B2(net150),
    .X(_03154_));
 sky130_fd_sc_hd__xnor2_1 _10008_ (.A(net191),
    .B(_03154_),
    .Y(_03155_));
 sky130_fd_sc_hd__nor2_1 _10009_ (.A(net177),
    .B(net4),
    .Y(_03156_));
 sky130_fd_sc_hd__xnor2_1 _10010_ (.A(net189),
    .B(_03156_),
    .Y(_03157_));
 sky130_fd_sc_hd__and2b_1 _10011_ (.A_N(_03157_),
    .B(_03155_),
    .X(_03158_));
 sky130_fd_sc_hd__and2b_1 _10012_ (.A_N(_03155_),
    .B(_03157_),
    .X(_03159_));
 sky130_fd_sc_hd__nor2_2 _10013_ (.A(_03158_),
    .B(_03159_),
    .Y(_03160_));
 sky130_fd_sc_hd__xnor2_2 _10014_ (.A(_03153_),
    .B(_03160_),
    .Y(_03161_));
 sky130_fd_sc_hd__o22a_1 _10015_ (.A1(net12),
    .A2(net133),
    .B1(net90),
    .B2(net45),
    .X(_03162_));
 sky130_fd_sc_hd__xnor2_1 _10016_ (.A(net97),
    .B(_03162_),
    .Y(_03163_));
 sky130_fd_sc_hd__o22a_1 _10017_ (.A1(net144),
    .A2(net8),
    .B1(net6),
    .B2(net147),
    .X(_03164_));
 sky130_fd_sc_hd__xnor2_1 _10018_ (.A(net33),
    .B(_03164_),
    .Y(_03165_));
 sky130_fd_sc_hd__o22a_1 _10019_ (.A1(net53),
    .A2(net92),
    .B1(net88),
    .B2(net14),
    .X(_03166_));
 sky130_fd_sc_hd__xnor2_1 _10020_ (.A(net112),
    .B(_03166_),
    .Y(_03167_));
 sky130_fd_sc_hd__and2_1 _10021_ (.A(_03165_),
    .B(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__xnor2_1 _10022_ (.A(_03165_),
    .B(_03167_),
    .Y(_03169_));
 sky130_fd_sc_hd__nor2_1 _10023_ (.A(_03163_),
    .B(_03169_),
    .Y(_03170_));
 sky130_fd_sc_hd__and2_1 _10024_ (.A(_03163_),
    .B(_03169_),
    .X(_03171_));
 sky130_fd_sc_hd__or2_1 _10025_ (.A(_03170_),
    .B(_03171_),
    .X(_03172_));
 sky130_fd_sc_hd__nor2_1 _10026_ (.A(_03161_),
    .B(_03172_),
    .Y(_03173_));
 sky130_fd_sc_hd__xor2_2 _10027_ (.A(_03161_),
    .B(_03172_),
    .X(_03174_));
 sky130_fd_sc_hd__xnor2_1 _10028_ (.A(_03141_),
    .B(_03174_),
    .Y(_03175_));
 sky130_fd_sc_hd__nor2_1 _10029_ (.A(_03136_),
    .B(_03175_),
    .Y(_03176_));
 sky130_fd_sc_hd__nand2_1 _10030_ (.A(_03136_),
    .B(_03175_),
    .Y(_03177_));
 sky130_fd_sc_hd__and2b_1 _10031_ (.A_N(_03176_),
    .B(_03177_),
    .X(_03178_));
 sky130_fd_sc_hd__xor2_4 _10032_ (.A(_03123_),
    .B(_03178_),
    .X(_03179_));
 sky130_fd_sc_hd__a21o_1 _10033_ (.A1(_02986_),
    .A2(_03043_),
    .B1(_03042_),
    .X(_03180_));
 sky130_fd_sc_hd__a21o_2 _10034_ (.A1(_02972_),
    .A2(_02985_),
    .B1(_02983_),
    .X(_03181_));
 sky130_fd_sc_hd__a21oi_4 _10035_ (.A1(_02987_),
    .A2(_02999_),
    .B1(_02998_),
    .Y(_03182_));
 sky130_fd_sc_hd__o21a_2 _10036_ (.A1(_03005_),
    .A2(_03038_),
    .B1(_03037_),
    .X(_03183_));
 sky130_fd_sc_hd__nor2_1 _10037_ (.A(_03182_),
    .B(_03183_),
    .Y(_03184_));
 sky130_fd_sc_hd__xor2_4 _10038_ (.A(_03182_),
    .B(_03183_),
    .X(_03185_));
 sky130_fd_sc_hd__xnor2_4 _10039_ (.A(_03181_),
    .B(_03185_),
    .Y(_03186_));
 sky130_fd_sc_hd__a21oi_4 _10040_ (.A1(_03046_),
    .A2(_03050_),
    .B1(_03049_),
    .Y(_03187_));
 sky130_fd_sc_hd__xnor2_2 _10041_ (.A(_03186_),
    .B(_03187_),
    .Y(_03188_));
 sky130_fd_sc_hd__and2b_1 _10042_ (.A_N(_03188_),
    .B(_03180_),
    .X(_03189_));
 sky130_fd_sc_hd__xnor2_2 _10043_ (.A(_03180_),
    .B(_03188_),
    .Y(_03190_));
 sky130_fd_sc_hd__and2_1 _10044_ (.A(_03179_),
    .B(_03190_),
    .X(_03191_));
 sky130_fd_sc_hd__xor2_4 _10045_ (.A(_03179_),
    .B(_03190_),
    .X(_03192_));
 sky130_fd_sc_hd__xnor2_4 _10046_ (.A(_03108_),
    .B(_03192_),
    .Y(_03193_));
 sky130_fd_sc_hd__nor2_1 _10047_ (.A(_03107_),
    .B(_03193_),
    .Y(_03194_));
 sky130_fd_sc_hd__xor2_4 _10048_ (.A(_03107_),
    .B(_03193_),
    .X(_03195_));
 sky130_fd_sc_hd__or2_1 _10049_ (.A(_02917_),
    .B(_03059_),
    .X(_03196_));
 sky130_fd_sc_hd__a21o_1 _10050_ (.A1(_02919_),
    .A2(_02925_),
    .B1(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__nand2_2 _10051_ (.A(_03061_),
    .B(_03197_),
    .Y(_03198_));
 sky130_fd_sc_hd__xnor2_4 _10052_ (.A(_03195_),
    .B(_03198_),
    .Y(_03199_));
 sky130_fd_sc_hd__or2_2 _10053_ (.A(_03064_),
    .B(_03065_),
    .X(_03200_));
 sky130_fd_sc_hd__a21oi_1 _10054_ (.A1(net19),
    .A2(_03200_),
    .B1(_03199_),
    .Y(_03201_));
 sky130_fd_sc_hd__a311oi_2 _10055_ (.A1(net19),
    .A2(_03199_),
    .A3(_03200_),
    .B1(_03201_),
    .C1(_02214_),
    .Y(_03202_));
 sky130_fd_sc_hd__o21ai_1 _10056_ (.A1(net86),
    .A2(_02171_),
    .B1(_02161_),
    .Y(_03203_));
 sky130_fd_sc_hd__o311a_1 _10057_ (.A1(net86),
    .A2(_02161_),
    .A3(_02171_),
    .B1(_02298_),
    .C1(_03203_),
    .X(_03204_));
 sky130_fd_sc_hd__a21oi_1 _10058_ (.A1(_06276_),
    .A2(_03071_),
    .B1(_06277_),
    .Y(_03205_));
 sky130_fd_sc_hd__nor2_1 _10059_ (.A(instruction[7]),
    .B(_03205_),
    .Y(_03206_));
 sky130_fd_sc_hd__a31o_1 _10060_ (.A1(instruction[7]),
    .A2(_06274_),
    .A3(_06314_),
    .B1(_03206_),
    .X(_03207_));
 sky130_fd_sc_hd__o21ai_1 _10061_ (.A1(_06269_),
    .A2(_03207_),
    .B1(net251),
    .Y(_03208_));
 sky130_fd_sc_hd__a21oi_2 _10062_ (.A1(_06269_),
    .A2(_03207_),
    .B1(_03208_),
    .Y(_03209_));
 sky130_fd_sc_hd__o21a_1 _10063_ (.A1(_03075_),
    .A2(_03076_),
    .B1(_03077_),
    .X(_03210_));
 sky130_fd_sc_hd__nor2_1 _10064_ (.A(reg1_val[6]),
    .B(curr_PC[6]),
    .Y(_03211_));
 sky130_fd_sc_hd__nand2_1 _10065_ (.A(reg1_val[6]),
    .B(curr_PC[6]),
    .Y(_03212_));
 sky130_fd_sc_hd__nand2b_1 _10066_ (.A_N(_03211_),
    .B(_03212_),
    .Y(_03213_));
 sky130_fd_sc_hd__xnor2_1 _10067_ (.A(_03210_),
    .B(_03213_),
    .Y(_03214_));
 sky130_fd_sc_hd__mux2_1 _10068_ (.A0(_02627_),
    .A1(_02630_),
    .S(net232),
    .X(_03215_));
 sky130_fd_sc_hd__nand2b_1 _10069_ (.A_N(_02634_),
    .B(net232),
    .Y(_03216_));
 sky130_fd_sc_hd__o21ai_1 _10070_ (.A1(net232),
    .A2(_02629_),
    .B1(_03216_),
    .Y(_03217_));
 sky130_fd_sc_hd__nand2_1 _10071_ (.A(net234),
    .B(_03217_),
    .Y(_03218_));
 sky130_fd_sc_hd__o211a_1 _10072_ (.A1(net234),
    .A2(_03215_),
    .B1(_03218_),
    .C1(net237),
    .X(_03219_));
 sky130_fd_sc_hd__mux2_1 _10073_ (.A0(_02633_),
    .A1(_02636_),
    .S(net232),
    .X(_03220_));
 sky130_fd_sc_hd__mux2_1 _10074_ (.A0(_03220_),
    .A1(_02442_),
    .S(net235),
    .X(_03221_));
 sky130_fd_sc_hd__a21oi_2 _10075_ (.A1(net239),
    .A2(_03221_),
    .B1(_03219_),
    .Y(_03222_));
 sky130_fd_sc_hd__mux2_1 _10076_ (.A0(_03214_),
    .A1(_03222_),
    .S(net241),
    .X(_03223_));
 sky130_fd_sc_hd__or3_1 _10077_ (.A(\div_res[5] ),
    .B(\div_res[4] ),
    .C(_02953_),
    .X(_03224_));
 sky130_fd_sc_hd__a21oi_1 _10078_ (.A1(net25),
    .A2(_03224_),
    .B1(\div_res[6] ),
    .Y(_03225_));
 sky130_fd_sc_hd__a31o_1 _10079_ (.A1(\div_res[6] ),
    .A2(net25),
    .A3(_03224_),
    .B1(net202),
    .X(_03226_));
 sky130_fd_sc_hd__or3_1 _10080_ (.A(\div_shifter[37] ),
    .B(\div_shifter[36] ),
    .C(_02956_),
    .X(_03227_));
 sky130_fd_sc_hd__a21oi_1 _10081_ (.A1(net246),
    .A2(_03227_),
    .B1(\div_shifter[38] ),
    .Y(_03228_));
 sky130_fd_sc_hd__a31o_1 _10082_ (.A1(\div_shifter[38] ),
    .A2(net246),
    .A3(_03227_),
    .B1(net249),
    .X(_03229_));
 sky130_fd_sc_hd__o2bb2a_1 _10083_ (.A1_N(_06265_),
    .A2_N(net213),
    .B1(_03228_),
    .B2(_03229_),
    .X(_03230_));
 sky130_fd_sc_hd__o221a_1 _10084_ (.A1(_06267_),
    .A2(_02291_),
    .B1(net204),
    .B2(_06268_),
    .C1(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__a21boi_1 _10085_ (.A1(_06269_),
    .A2(_02294_),
    .B1_N(_03231_),
    .Y(_03232_));
 sky130_fd_sc_hd__o21a_1 _10086_ (.A1(_03225_),
    .A2(_03226_),
    .B1(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__o21a_1 _10087_ (.A1(net235),
    .A2(_02473_),
    .B1(_02318_),
    .X(_03234_));
 sky130_fd_sc_hd__o21ai_2 _10088_ (.A1(net239),
    .A2(_03234_),
    .B1(_02312_),
    .Y(_03235_));
 sky130_fd_sc_hd__o221a_1 _10089_ (.A1(net182),
    .A2(_03222_),
    .B1(_03235_),
    .B2(net185),
    .C1(_03233_),
    .X(_03236_));
 sky130_fd_sc_hd__o21ai_2 _10090_ (.A1(net214),
    .A2(_03223_),
    .B1(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__or4_2 _10091_ (.A(_03202_),
    .B(_03204_),
    .C(_03209_),
    .D(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__and2_1 _10092_ (.A(curr_PC[6]),
    .B(_03105_),
    .X(_03239_));
 sky130_fd_sc_hd__o21ai_1 _10093_ (.A1(curr_PC[6]),
    .A2(_03105_),
    .B1(net262),
    .Y(_03240_));
 sky130_fd_sc_hd__a2bb2o_4 _10094_ (.A1_N(_03239_),
    .A2_N(_03240_),
    .B1(net257),
    .B2(_03238_),
    .X(dest_val[6]));
 sky130_fd_sc_hd__a21oi_4 _10095_ (.A1(_03108_),
    .A2(_03192_),
    .B1(_03191_),
    .Y(_03241_));
 sky130_fd_sc_hd__o21bai_4 _10096_ (.A1(_03186_),
    .A2(_03187_),
    .B1_N(_03189_),
    .Y(_03242_));
 sky130_fd_sc_hd__o21bai_4 _10097_ (.A1(_03153_),
    .A2(_03160_),
    .B1_N(_03152_),
    .Y(_03243_));
 sky130_fd_sc_hd__a21oi_4 _10098_ (.A1(_03137_),
    .A2(_03139_),
    .B1(_03138_),
    .Y(_03244_));
 sky130_fd_sc_hd__o22a_1 _10099_ (.A1(net128),
    .A2(net51),
    .B1(net48),
    .B2(net100),
    .X(_03245_));
 sky130_fd_sc_hd__xnor2_1 _10100_ (.A(net105),
    .B(_03245_),
    .Y(_03246_));
 sky130_fd_sc_hd__o22a_1 _10101_ (.A1(net77),
    .A2(net36),
    .B1(net34),
    .B2(net74),
    .X(_03247_));
 sky130_fd_sc_hd__xnor2_1 _10102_ (.A(net135),
    .B(_03247_),
    .Y(_03248_));
 sky130_fd_sc_hd__and2_1 _10103_ (.A(_03246_),
    .B(_03248_),
    .X(_03249_));
 sky130_fd_sc_hd__nor2_1 _10104_ (.A(_03246_),
    .B(_03248_),
    .Y(_03250_));
 sky130_fd_sc_hd__nor2_2 _10105_ (.A(_03249_),
    .B(_03250_),
    .Y(_03251_));
 sky130_fd_sc_hd__o22a_2 _10106_ (.A1(net119),
    .A2(net40),
    .B1(net38),
    .B2(net71),
    .X(_03252_));
 sky130_fd_sc_hd__xnor2_4 _10107_ (.A(net102),
    .B(_03252_),
    .Y(_03253_));
 sky130_fd_sc_hd__xnor2_4 _10108_ (.A(_03251_),
    .B(_03253_),
    .Y(_03254_));
 sky130_fd_sc_hd__nor2_1 _10109_ (.A(_03244_),
    .B(_03254_),
    .Y(_03255_));
 sky130_fd_sc_hd__xor2_4 _10110_ (.A(_03244_),
    .B(_03254_),
    .X(_03256_));
 sky130_fd_sc_hd__xnor2_4 _10111_ (.A(_03243_),
    .B(_03256_),
    .Y(_03257_));
 sky130_fd_sc_hd__o22a_1 _10112_ (.A1(net8),
    .A2(net133),
    .B1(net6),
    .B2(net144),
    .X(_03258_));
 sky130_fd_sc_hd__xnor2_1 _10113_ (.A(net31),
    .B(_03258_),
    .Y(_03259_));
 sky130_fd_sc_hd__nor2_1 _10114_ (.A(_03158_),
    .B(_03259_),
    .Y(_03260_));
 sky130_fd_sc_hd__and2_1 _10115_ (.A(_03158_),
    .B(_03259_),
    .X(_03261_));
 sky130_fd_sc_hd__nor2_1 _10116_ (.A(_03260_),
    .B(_03261_),
    .Y(_03262_));
 sky130_fd_sc_hd__nor2_1 _10117_ (.A(net147),
    .B(net31),
    .Y(_03263_));
 sky130_fd_sc_hd__xnor2_1 _10118_ (.A(_03262_),
    .B(_03263_),
    .Y(_03264_));
 sky130_fd_sc_hd__a21o_1 _10119_ (.A1(_03147_),
    .A2(_03149_),
    .B1(_03146_),
    .X(_03265_));
 sky130_fd_sc_hd__o22a_1 _10120_ (.A1(net152),
    .A2(net9),
    .B1(net3),
    .B2(net150),
    .X(_03266_));
 sky130_fd_sc_hd__xnor2_1 _10121_ (.A(_06490_),
    .B(_03266_),
    .Y(_03267_));
 sky130_fd_sc_hd__nand3_1 _10122_ (.A(_00151_),
    .B(_00219_),
    .C(_00221_),
    .Y(_03268_));
 sky130_fd_sc_hd__a21o_1 _10123_ (.A1(_00225_),
    .A2(_00226_),
    .B1(net114),
    .X(_03269_));
 sky130_fd_sc_hd__a21o_1 _10124_ (.A1(_03268_),
    .A2(_03269_),
    .B1(net179),
    .X(_03270_));
 sky130_fd_sc_hd__nand3_1 _10125_ (.A(net179),
    .B(_03268_),
    .C(_03269_),
    .Y(_03271_));
 sky130_fd_sc_hd__nand3_1 _10126_ (.A(net189),
    .B(_03270_),
    .C(_03271_),
    .Y(_03272_));
 sky130_fd_sc_hd__a21o_1 _10127_ (.A1(_03270_),
    .A2(_03271_),
    .B1(net189),
    .X(_03273_));
 sky130_fd_sc_hd__nand3_1 _10128_ (.A(_03267_),
    .B(_03272_),
    .C(_03273_),
    .Y(_03274_));
 sky130_fd_sc_hd__a21o_1 _10129_ (.A1(_03272_),
    .A2(_03273_),
    .B1(_03267_),
    .X(_03275_));
 sky130_fd_sc_hd__nand3_1 _10130_ (.A(_03265_),
    .B(_03274_),
    .C(_03275_),
    .Y(_03276_));
 sky130_fd_sc_hd__a21o_1 _10131_ (.A1(_03274_),
    .A2(_03275_),
    .B1(_03265_),
    .X(_03277_));
 sky130_fd_sc_hd__nand3_1 _10132_ (.A(_03129_),
    .B(_03276_),
    .C(_03277_),
    .Y(_03278_));
 sky130_fd_sc_hd__a21o_1 _10133_ (.A1(_03276_),
    .A2(_03277_),
    .B1(_03129_),
    .X(_03279_));
 sky130_fd_sc_hd__o32a_1 _10134_ (.A1(_00334_),
    .A2(_00335_),
    .A3(net90),
    .B1(net87),
    .B2(net45),
    .X(_03280_));
 sky130_fd_sc_hd__xnor2_1 _10135_ (.A(net97),
    .B(_03280_),
    .Y(_03281_));
 sky130_fd_sc_hd__a22o_1 _10136_ (.A1(_06483_),
    .A2(_00307_),
    .B1(_00308_),
    .B2(_06459_),
    .X(_03282_));
 sky130_fd_sc_hd__xor2_1 _10137_ (.A(net108),
    .B(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__nand2b_1 _10138_ (.A_N(_03281_),
    .B(_03283_),
    .Y(_03284_));
 sky130_fd_sc_hd__xor2_1 _10139_ (.A(_03281_),
    .B(_03283_),
    .X(_03285_));
 sky130_fd_sc_hd__o22a_1 _10140_ (.A1(net126),
    .A2(net53),
    .B1(net92),
    .B2(net15),
    .X(_03286_));
 sky130_fd_sc_hd__xnor2_1 _10141_ (.A(net112),
    .B(_03286_),
    .Y(_03287_));
 sky130_fd_sc_hd__nand2b_1 _10142_ (.A_N(_03285_),
    .B(_03287_),
    .Y(_03288_));
 sky130_fd_sc_hd__xnor2_1 _10143_ (.A(_03285_),
    .B(_03287_),
    .Y(_03289_));
 sky130_fd_sc_hd__and3_1 _10144_ (.A(_03278_),
    .B(_03279_),
    .C(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__a21oi_1 _10145_ (.A1(_03278_),
    .A2(_03279_),
    .B1(_03289_),
    .Y(_03291_));
 sky130_fd_sc_hd__or3_1 _10146_ (.A(_03264_),
    .B(_03290_),
    .C(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__o21ai_1 _10147_ (.A1(_03290_),
    .A2(_03291_),
    .B1(_03264_),
    .Y(_03293_));
 sky130_fd_sc_hd__a21o_1 _10148_ (.A1(_03116_),
    .A2(_03118_),
    .B1(_03114_),
    .X(_03294_));
 sky130_fd_sc_hd__o22a_1 _10149_ (.A1(net82),
    .A2(net63),
    .B1(net60),
    .B2(net130),
    .X(_03295_));
 sky130_fd_sc_hd__xnor2_1 _10150_ (.A(net157),
    .B(_03295_),
    .Y(_03296_));
 sky130_fd_sc_hd__o22a_1 _10151_ (.A1(net67),
    .A2(net42),
    .B1(net94),
    .B2(net64),
    .X(_03297_));
 sky130_fd_sc_hd__xnor2_1 _10152_ (.A(net137),
    .B(_03297_),
    .Y(_03298_));
 sky130_fd_sc_hd__nand2b_1 _10153_ (.A_N(_03296_),
    .B(_03298_),
    .Y(_03299_));
 sky130_fd_sc_hd__xor2_1 _10154_ (.A(_03296_),
    .B(_03298_),
    .X(_03300_));
 sky130_fd_sc_hd__o22a_1 _10155_ (.A1(net78),
    .A2(net58),
    .B1(net55),
    .B2(net123),
    .X(_03301_));
 sky130_fd_sc_hd__xor2_1 _10156_ (.A(net155),
    .B(_03301_),
    .X(_03302_));
 sky130_fd_sc_hd__xnor2_1 _10157_ (.A(_03300_),
    .B(_03302_),
    .Y(_03303_));
 sky130_fd_sc_hd__o21ba_1 _10158_ (.A1(_03168_),
    .A2(_03170_),
    .B1_N(_03303_),
    .X(_03304_));
 sky130_fd_sc_hd__or3b_1 _10159_ (.A(_03168_),
    .B(_03170_),
    .C_N(_03303_),
    .X(_03305_));
 sky130_fd_sc_hd__nand2b_1 _10160_ (.A_N(_03304_),
    .B(_03305_),
    .Y(_03306_));
 sky130_fd_sc_hd__xnor2_1 _10161_ (.A(_03294_),
    .B(_03306_),
    .Y(_03307_));
 sky130_fd_sc_hd__and3_1 _10162_ (.A(_03292_),
    .B(_03293_),
    .C(_03307_),
    .X(_03308_));
 sky130_fd_sc_hd__a21oi_1 _10163_ (.A1(_03292_),
    .A2(_03293_),
    .B1(_03307_),
    .Y(_03309_));
 sky130_fd_sc_hd__nor2_2 _10164_ (.A(_03308_),
    .B(_03309_),
    .Y(_03310_));
 sky130_fd_sc_hd__xnor2_4 _10165_ (.A(_03257_),
    .B(_03310_),
    .Y(_03311_));
 sky130_fd_sc_hd__a21o_1 _10166_ (.A1(_03123_),
    .A2(_03177_),
    .B1(_03176_),
    .X(_03312_));
 sky130_fd_sc_hd__a21bo_1 _10167_ (.A1(_03119_),
    .A2(_03120_),
    .B1_N(_03122_),
    .X(_03313_));
 sky130_fd_sc_hd__nand2_1 _10168_ (.A(_03132_),
    .B(_03135_),
    .Y(_03314_));
 sky130_fd_sc_hd__a21oi_2 _10169_ (.A1(_03141_),
    .A2(_03174_),
    .B1(_03173_),
    .Y(_03315_));
 sky130_fd_sc_hd__a21o_1 _10170_ (.A1(_03132_),
    .A2(_03135_),
    .B1(_03315_),
    .X(_03316_));
 sky130_fd_sc_hd__xnor2_2 _10171_ (.A(_03314_),
    .B(_03315_),
    .Y(_03317_));
 sky130_fd_sc_hd__xnor2_2 _10172_ (.A(_03313_),
    .B(_03317_),
    .Y(_03318_));
 sky130_fd_sc_hd__a21oi_2 _10173_ (.A1(_03181_),
    .A2(_03185_),
    .B1(_03184_),
    .Y(_03319_));
 sky130_fd_sc_hd__nor2_1 _10174_ (.A(_03318_),
    .B(_03319_),
    .Y(_03320_));
 sky130_fd_sc_hd__xnor2_2 _10175_ (.A(_03318_),
    .B(_03319_),
    .Y(_03321_));
 sky130_fd_sc_hd__and2b_1 _10176_ (.A_N(_03321_),
    .B(_03312_),
    .X(_03322_));
 sky130_fd_sc_hd__xnor2_2 _10177_ (.A(_03312_),
    .B(_03321_),
    .Y(_03323_));
 sky130_fd_sc_hd__and2_1 _10178_ (.A(_03311_),
    .B(_03323_),
    .X(_03324_));
 sky130_fd_sc_hd__xor2_4 _10179_ (.A(_03311_),
    .B(_03323_),
    .X(_03325_));
 sky130_fd_sc_hd__xnor2_4 _10180_ (.A(_03242_),
    .B(_03325_),
    .Y(_03326_));
 sky130_fd_sc_hd__xor2_4 _10181_ (.A(_03241_),
    .B(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__a31o_1 _10182_ (.A1(_03061_),
    .A2(_03195_),
    .A3(_03197_),
    .B1(_03194_),
    .X(_03328_));
 sky130_fd_sc_hd__xor2_4 _10183_ (.A(_03327_),
    .B(_03328_),
    .X(_03329_));
 sky130_fd_sc_hd__o21a_1 _10184_ (.A1(_03199_),
    .A2(_03200_),
    .B1(net19),
    .X(_03330_));
 sky130_fd_sc_hd__o21ai_1 _10185_ (.A1(_03329_),
    .A2(_03330_),
    .B1(net206),
    .Y(_03331_));
 sky130_fd_sc_hd__a21oi_1 _10186_ (.A1(_03329_),
    .A2(_03330_),
    .B1(_03331_),
    .Y(_03332_));
 sky130_fd_sc_hd__nand3_1 _10187_ (.A(net19),
    .B(_02160_),
    .C(_02172_),
    .Y(_03333_));
 sky130_fd_sc_hd__a21o_1 _10188_ (.A1(net19),
    .A2(_02172_),
    .B1(_02160_),
    .X(_03334_));
 sky130_fd_sc_hd__o21a_1 _10189_ (.A1(_06267_),
    .A2(_03205_),
    .B1(_06268_),
    .X(_03335_));
 sky130_fd_sc_hd__mux2_1 _10190_ (.A0(_06316_),
    .A1(_03335_),
    .S(net300),
    .X(_03336_));
 sky130_fd_sc_hd__a21oi_1 _10191_ (.A1(_06263_),
    .A2(_03336_),
    .B1(_02293_),
    .Y(_03337_));
 sky130_fd_sc_hd__o21a_1 _10192_ (.A1(_06263_),
    .A2(_03336_),
    .B1(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__o21a_1 _10193_ (.A1(_03210_),
    .A2(_03211_),
    .B1(_03212_),
    .X(_03339_));
 sky130_fd_sc_hd__nor2_1 _10194_ (.A(reg1_val[7]),
    .B(curr_PC[7]),
    .Y(_03340_));
 sky130_fd_sc_hd__nand2_1 _10195_ (.A(reg1_val[7]),
    .B(curr_PC[7]),
    .Y(_03341_));
 sky130_fd_sc_hd__and2b_1 _10196_ (.A_N(_03340_),
    .B(_03341_),
    .X(_03342_));
 sky130_fd_sc_hd__xnor2_1 _10197_ (.A(_03339_),
    .B(_03342_),
    .Y(_03343_));
 sky130_fd_sc_hd__mux2_1 _10198_ (.A0(_02774_),
    .A1(_02777_),
    .S(net231),
    .X(_03344_));
 sky130_fd_sc_hd__mux2_1 _10199_ (.A0(_02776_),
    .A1(_02781_),
    .S(net231),
    .X(_03345_));
 sky130_fd_sc_hd__mux2_1 _10200_ (.A0(_03344_),
    .A1(_03345_),
    .S(net235),
    .X(_03346_));
 sky130_fd_sc_hd__mux2_1 _10201_ (.A0(_02780_),
    .A1(_02783_),
    .S(net231),
    .X(_03347_));
 sky130_fd_sc_hd__mux2_1 _10202_ (.A0(_03347_),
    .A1(_02317_),
    .S(net235),
    .X(_03348_));
 sky130_fd_sc_hd__mux2_1 _10203_ (.A0(_03346_),
    .A1(_03348_),
    .S(net239),
    .X(_03349_));
 sky130_fd_sc_hd__inv_2 _10204_ (.A(_03349_),
    .Y(_03350_));
 sky130_fd_sc_hd__or2_1 _10205_ (.A(net242),
    .B(_03343_),
    .X(_03351_));
 sky130_fd_sc_hd__o211a_1 _10206_ (.A1(net263),
    .A2(_03349_),
    .B1(_03351_),
    .C1(net215),
    .X(_03352_));
 sky130_fd_sc_hd__or2_1 _10207_ (.A(\div_res[6] ),
    .B(_03224_),
    .X(_03353_));
 sky130_fd_sc_hd__and3_1 _10208_ (.A(\div_res[7] ),
    .B(net25),
    .C(_03353_),
    .X(_03354_));
 sky130_fd_sc_hd__a21oi_1 _10209_ (.A1(net25),
    .A2(_03353_),
    .B1(\div_res[7] ),
    .Y(_03355_));
 sky130_fd_sc_hd__or2_1 _10210_ (.A(\div_shifter[38] ),
    .B(_03227_),
    .X(_03356_));
 sky130_fd_sc_hd__a21oi_1 _10211_ (.A1(net246),
    .A2(_03356_),
    .B1(\div_shifter[39] ),
    .Y(_03357_));
 sky130_fd_sc_hd__a31o_1 _10212_ (.A1(\div_shifter[39] ),
    .A2(net246),
    .A3(_03356_),
    .B1(net249),
    .X(_03358_));
 sky130_fd_sc_hd__a2bb2o_1 _10213_ (.A1_N(_03357_),
    .A2_N(_03358_),
    .B1(_06258_),
    .B2(net213),
    .X(_03359_));
 sky130_fd_sc_hd__a21oi_1 _10214_ (.A1(_06261_),
    .A2(net205),
    .B1(_03359_),
    .Y(_03360_));
 sky130_fd_sc_hd__o221a_1 _10215_ (.A1(_06263_),
    .A2(_02295_),
    .B1(_02301_),
    .B2(_06262_),
    .C1(_03360_),
    .X(_03361_));
 sky130_fd_sc_hd__o31a_1 _10216_ (.A1(net202),
    .A2(_03354_),
    .A3(_03355_),
    .B1(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__o21a_1 _10217_ (.A1(net234),
    .A2(_02280_),
    .B1(_02318_),
    .X(_03363_));
 sky130_fd_sc_hd__o21ai_2 _10218_ (.A1(net239),
    .A2(_03363_),
    .B1(_02312_),
    .Y(_03364_));
 sky130_fd_sc_hd__o221a_1 _10219_ (.A1(net183),
    .A2(_03350_),
    .B1(_03364_),
    .B2(net185),
    .C1(_03362_),
    .X(_03365_));
 sky130_fd_sc_hd__or3b_2 _10220_ (.A(_03338_),
    .B(_03352_),
    .C_N(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__a311o_1 _10221_ (.A1(_02298_),
    .A2(_03333_),
    .A3(_03334_),
    .B1(_03366_),
    .C1(_03332_),
    .X(_03367_));
 sky130_fd_sc_hd__or2_1 _10222_ (.A(curr_PC[7]),
    .B(_03239_),
    .X(_03368_));
 sky130_fd_sc_hd__a21oi_1 _10223_ (.A1(curr_PC[7]),
    .A2(_03239_),
    .B1(net257),
    .Y(_03369_));
 sky130_fd_sc_hd__a22o_4 _10224_ (.A1(net257),
    .A2(_03367_),
    .B1(_03368_),
    .B2(_03369_),
    .X(dest_val[7]));
 sky130_fd_sc_hd__a21o_1 _10225_ (.A1(_03242_),
    .A2(_03325_),
    .B1(_03324_),
    .X(_03370_));
 sky130_fd_sc_hd__a32o_1 _10226_ (.A1(_06461_),
    .A2(_00219_),
    .A3(_00221_),
    .B1(_00197_),
    .B2(_06445_),
    .X(_03371_));
 sky130_fd_sc_hd__xnor2_1 _10227_ (.A(net157),
    .B(_03371_),
    .Y(_03372_));
 sky130_fd_sc_hd__o22a_1 _10228_ (.A1(net123),
    .A2(net63),
    .B1(net55),
    .B2(net78),
    .X(_03373_));
 sky130_fd_sc_hd__xnor2_1 _10229_ (.A(net154),
    .B(_03373_),
    .Y(_03374_));
 sky130_fd_sc_hd__xnor2_1 _10230_ (.A(_03372_),
    .B(_03374_),
    .Y(_03375_));
 sky130_fd_sc_hd__a21oi_1 _10231_ (.A1(_03284_),
    .A2(_03288_),
    .B1(_03375_),
    .Y(_03376_));
 sky130_fd_sc_hd__and3_1 _10232_ (.A(_03284_),
    .B(_03288_),
    .C(_03375_),
    .X(_03377_));
 sky130_fd_sc_hd__or2_1 _10233_ (.A(_03376_),
    .B(_03377_),
    .X(_03378_));
 sky130_fd_sc_hd__a21o_1 _10234_ (.A1(_03251_),
    .A2(_03253_),
    .B1(_03249_),
    .X(_03379_));
 sky130_fd_sc_hd__and2b_1 _10235_ (.A_N(_03378_),
    .B(_03379_),
    .X(_03380_));
 sky130_fd_sc_hd__xor2_1 _10236_ (.A(_03378_),
    .B(_03379_),
    .X(_03381_));
 sky130_fd_sc_hd__o22a_1 _10237_ (.A1(_00421_),
    .A2(net90),
    .B1(net6),
    .B2(net133),
    .X(_03382_));
 sky130_fd_sc_hd__xnor2_1 _10238_ (.A(net29),
    .B(_03382_),
    .Y(_03383_));
 sky130_fd_sc_hd__nor2_1 _10239_ (.A(net144),
    .B(net29),
    .Y(_03384_));
 sky130_fd_sc_hd__o22a_1 _10240_ (.A1(net44),
    .A2(net92),
    .B1(net88),
    .B2(net11),
    .X(_03385_));
 sky130_fd_sc_hd__xor2_1 _10241_ (.A(net96),
    .B(_03385_),
    .X(_03386_));
 sky130_fd_sc_hd__and2_1 _10242_ (.A(_03384_),
    .B(_03386_),
    .X(_03387_));
 sky130_fd_sc_hd__xnor2_1 _10243_ (.A(_03384_),
    .B(_03386_),
    .Y(_03388_));
 sky130_fd_sc_hd__nor2_1 _10244_ (.A(_03383_),
    .B(_03388_),
    .Y(_03389_));
 sky130_fd_sc_hd__and2_1 _10245_ (.A(_03383_),
    .B(_03388_),
    .X(_03390_));
 sky130_fd_sc_hd__nor2_1 _10246_ (.A(_03389_),
    .B(_03390_),
    .Y(_03391_));
 sky130_fd_sc_hd__o21ai_1 _10247_ (.A1(_03300_),
    .A2(_03302_),
    .B1(_03299_),
    .Y(_03392_));
 sky130_fd_sc_hd__a21boi_1 _10248_ (.A1(_03267_),
    .A2(_03273_),
    .B1_N(_03272_),
    .Y(_03393_));
 sky130_fd_sc_hd__o22a_1 _10249_ (.A1(net116),
    .A2(net16),
    .B1(net9),
    .B2(net114),
    .X(_03394_));
 sky130_fd_sc_hd__xnor2_1 _10250_ (.A(net179),
    .B(_03394_),
    .Y(_03395_));
 sky130_fd_sc_hd__nand2_1 _10251_ (.A(_06498_),
    .B(_00756_),
    .Y(_03396_));
 sky130_fd_sc_hd__xnor2_1 _10252_ (.A(net191),
    .B(_03396_),
    .Y(_03397_));
 sky130_fd_sc_hd__nand2_1 _10253_ (.A(_03395_),
    .B(_03397_),
    .Y(_03398_));
 sky130_fd_sc_hd__xnor2_1 _10254_ (.A(_03395_),
    .B(_03397_),
    .Y(_03399_));
 sky130_fd_sc_hd__and2b_1 _10255_ (.A_N(_03393_),
    .B(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__xnor2_1 _10256_ (.A(_03393_),
    .B(_03399_),
    .Y(_03401_));
 sky130_fd_sc_hd__xor2_1 _10257_ (.A(_03392_),
    .B(_03401_),
    .X(_03402_));
 sky130_fd_sc_hd__o22a_1 _10258_ (.A1(net126),
    .A2(net14),
    .B1(net52),
    .B2(net121),
    .X(_03403_));
 sky130_fd_sc_hd__xor2_1 _10259_ (.A(net111),
    .B(_03403_),
    .X(_03404_));
 sky130_fd_sc_hd__o22a_1 _10260_ (.A1(net118),
    .A2(net48),
    .B1(net100),
    .B2(net50),
    .X(_03405_));
 sky130_fd_sc_hd__xor2_1 _10261_ (.A(net105),
    .B(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__nor2_1 _10262_ (.A(_03404_),
    .B(_03406_),
    .Y(_03407_));
 sky130_fd_sc_hd__xor2_1 _10263_ (.A(_03404_),
    .B(_03406_),
    .X(_03408_));
 sky130_fd_sc_hd__a22o_1 _10264_ (.A1(_06459_),
    .A2(_00307_),
    .B1(_00308_),
    .B2(_06467_),
    .X(_03409_));
 sky130_fd_sc_hd__xor2_1 _10265_ (.A(net108),
    .B(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__and2_1 _10266_ (.A(_03408_),
    .B(_03410_),
    .X(_03411_));
 sky130_fd_sc_hd__nor2_1 _10267_ (.A(_03408_),
    .B(_03410_),
    .Y(_03412_));
 sky130_fd_sc_hd__nor2_1 _10268_ (.A(_03411_),
    .B(_03412_),
    .Y(_03413_));
 sky130_fd_sc_hd__and2_1 _10269_ (.A(_03402_),
    .B(_03413_),
    .X(_03414_));
 sky130_fd_sc_hd__xor2_1 _10270_ (.A(_03402_),
    .B(_03413_),
    .X(_03415_));
 sky130_fd_sc_hd__xnor2_1 _10271_ (.A(_03391_),
    .B(_03415_),
    .Y(_03416_));
 sky130_fd_sc_hd__nor2_1 _10272_ (.A(_03381_),
    .B(_03416_),
    .Y(_03417_));
 sky130_fd_sc_hd__nand2_1 _10273_ (.A(_03381_),
    .B(_03416_),
    .Y(_03418_));
 sky130_fd_sc_hd__and2b_1 _10274_ (.A_N(_03417_),
    .B(_03418_),
    .X(_03419_));
 sky130_fd_sc_hd__nand2_1 _10275_ (.A(_03276_),
    .B(_03278_),
    .Y(_03420_));
 sky130_fd_sc_hd__o22a_1 _10276_ (.A1(net65),
    .A2(net42),
    .B1(net94),
    .B2(net58),
    .X(_03421_));
 sky130_fd_sc_hd__xnor2_1 _10277_ (.A(net137),
    .B(_03421_),
    .Y(_03422_));
 sky130_fd_sc_hd__o22a_1 _10278_ (.A1(net71),
    .A2(net40),
    .B1(net38),
    .B2(net77),
    .X(_03423_));
 sky130_fd_sc_hd__xnor2_1 _10279_ (.A(net102),
    .B(_03423_),
    .Y(_03424_));
 sky130_fd_sc_hd__and2_1 _10280_ (.A(_03422_),
    .B(_03424_),
    .X(_03425_));
 sky130_fd_sc_hd__nor2_1 _10281_ (.A(_03422_),
    .B(_03424_),
    .Y(_03426_));
 sky130_fd_sc_hd__nor2_1 _10282_ (.A(_03425_),
    .B(_03426_),
    .Y(_03427_));
 sky130_fd_sc_hd__o22a_1 _10283_ (.A1(net73),
    .A2(net36),
    .B1(net34),
    .B2(net67),
    .X(_03428_));
 sky130_fd_sc_hd__xnor2_1 _10284_ (.A(net135),
    .B(_03428_),
    .Y(_03429_));
 sky130_fd_sc_hd__xor2_1 _10285_ (.A(_03427_),
    .B(_03429_),
    .X(_03430_));
 sky130_fd_sc_hd__a21o_1 _10286_ (.A1(_03262_),
    .A2(_03263_),
    .B1(_03260_),
    .X(_03431_));
 sky130_fd_sc_hd__nand2_1 _10287_ (.A(_03430_),
    .B(_03431_),
    .Y(_03432_));
 sky130_fd_sc_hd__xor2_1 _10288_ (.A(_03430_),
    .B(_03431_),
    .X(_03433_));
 sky130_fd_sc_hd__xor2_1 _10289_ (.A(_03420_),
    .B(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__xnor2_1 _10290_ (.A(_03419_),
    .B(_03434_),
    .Y(_03435_));
 sky130_fd_sc_hd__o21bai_1 _10291_ (.A1(_03257_),
    .A2(_03309_),
    .B1_N(_03308_),
    .Y(_03436_));
 sky130_fd_sc_hd__a21bo_1 _10292_ (.A1(_03313_),
    .A2(_03317_),
    .B1_N(_03316_),
    .X(_03437_));
 sky130_fd_sc_hd__a21o_1 _10293_ (.A1(_03243_),
    .A2(_03256_),
    .B1(_03255_),
    .X(_03438_));
 sky130_fd_sc_hd__o21ba_1 _10294_ (.A1(_03264_),
    .A2(_03291_),
    .B1_N(_03290_),
    .X(_03439_));
 sky130_fd_sc_hd__a21oi_1 _10295_ (.A1(_03294_),
    .A2(_03305_),
    .B1(_03304_),
    .Y(_03440_));
 sky130_fd_sc_hd__nor2_1 _10296_ (.A(_03439_),
    .B(_03440_),
    .Y(_03441_));
 sky130_fd_sc_hd__xor2_1 _10297_ (.A(_03439_),
    .B(_03440_),
    .X(_03442_));
 sky130_fd_sc_hd__xnor2_1 _10298_ (.A(_03438_),
    .B(_03442_),
    .Y(_03443_));
 sky130_fd_sc_hd__nand2b_1 _10299_ (.A_N(_03443_),
    .B(_03437_),
    .Y(_03444_));
 sky130_fd_sc_hd__xnor2_1 _10300_ (.A(_03437_),
    .B(_03443_),
    .Y(_03445_));
 sky130_fd_sc_hd__xnor2_1 _10301_ (.A(_03436_),
    .B(_03445_),
    .Y(_03446_));
 sky130_fd_sc_hd__or2_1 _10302_ (.A(_03435_),
    .B(_03446_),
    .X(_03447_));
 sky130_fd_sc_hd__xor2_1 _10303_ (.A(_03435_),
    .B(_03446_),
    .X(_03448_));
 sky130_fd_sc_hd__o21ai_2 _10304_ (.A1(_03320_),
    .A2(_03322_),
    .B1(_03448_),
    .Y(_03449_));
 sky130_fd_sc_hd__or3_1 _10305_ (.A(_03320_),
    .B(_03322_),
    .C(_03448_),
    .X(_03450_));
 sky130_fd_sc_hd__and2_1 _10306_ (.A(_03449_),
    .B(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__nand2_1 _10307_ (.A(_03370_),
    .B(_03451_),
    .Y(_03452_));
 sky130_fd_sc_hd__xnor2_2 _10308_ (.A(_03370_),
    .B(_03451_),
    .Y(_03453_));
 sky130_fd_sc_hd__nand2_1 _10309_ (.A(_03195_),
    .B(_03327_),
    .Y(_03454_));
 sky130_fd_sc_hd__or4b_2 _10310_ (.A(_03059_),
    .B(_03060_),
    .C(_03454_),
    .D_N(_02919_),
    .X(_03455_));
 sky130_fd_sc_hd__or3b_1 _10311_ (.A(_03060_),
    .B(_03454_),
    .C_N(_03196_),
    .X(_03456_));
 sky130_fd_sc_hd__o22a_1 _10312_ (.A1(_03107_),
    .A2(_03193_),
    .B1(_03241_),
    .B2(_03326_),
    .X(_03457_));
 sky130_fd_sc_hd__a21oi_1 _10313_ (.A1(_03241_),
    .A2(_03326_),
    .B1(_03457_),
    .Y(_03458_));
 sky130_fd_sc_hd__inv_2 _10314_ (.A(_03458_),
    .Y(_03459_));
 sky130_fd_sc_hd__o211a_1 _10315_ (.A1(_02922_),
    .A2(_03455_),
    .B1(_03456_),
    .C1(_03459_),
    .X(_03460_));
 sky130_fd_sc_hd__nor2_1 _10316_ (.A(_02923_),
    .B(_03455_),
    .Y(_03461_));
 sky130_fd_sc_hd__a21bo_2 _10317_ (.A1(_02035_),
    .A2(_03461_),
    .B1_N(_03460_),
    .X(_03462_));
 sky130_fd_sc_hd__nand2b_1 _10318_ (.A_N(_03453_),
    .B(_03462_),
    .Y(_03463_));
 sky130_fd_sc_hd__xor2_2 _10319_ (.A(_03453_),
    .B(_03462_),
    .X(_03464_));
 sky130_fd_sc_hd__or2_1 _10320_ (.A(_02212_),
    .B(_02926_),
    .X(_03465_));
 sky130_fd_sc_hd__or4_2 _10321_ (.A(_02766_),
    .B(_02767_),
    .C(_03064_),
    .D(_03465_),
    .X(_03466_));
 sky130_fd_sc_hd__o31ai_1 _10322_ (.A1(_03199_),
    .A2(_03329_),
    .A3(_03466_),
    .B1(net27),
    .Y(_03467_));
 sky130_fd_sc_hd__o21ai_1 _10323_ (.A1(_03464_),
    .A2(_03467_),
    .B1(net206),
    .Y(_03468_));
 sky130_fd_sc_hd__a21o_1 _10324_ (.A1(_03464_),
    .A2(_03467_),
    .B1(_03468_),
    .X(_03469_));
 sky130_fd_sc_hd__a21oi_1 _10325_ (.A1(net19),
    .A2(_02173_),
    .B1(_02159_),
    .Y(_03470_));
 sky130_fd_sc_hd__a31o_1 _10326_ (.A1(net19),
    .A2(_02159_),
    .A3(_02173_),
    .B1(net250),
    .X(_03471_));
 sky130_fd_sc_hd__or2_1 _10327_ (.A(_03470_),
    .B(_03471_),
    .X(_03472_));
 sky130_fd_sc_hd__or3_1 _10328_ (.A(net300),
    .B(_06259_),
    .C(_06317_),
    .X(_03473_));
 sky130_fd_sc_hd__o21a_1 _10329_ (.A1(_06260_),
    .A2(_03335_),
    .B1(_06262_),
    .X(_03474_));
 sky130_fd_sc_hd__o21a_1 _10330_ (.A1(instruction[7]),
    .A2(_03474_),
    .B1(_03473_),
    .X(_03475_));
 sky130_fd_sc_hd__nor2_1 _10331_ (.A(_06256_),
    .B(_03475_),
    .Y(_03476_));
 sky130_fd_sc_hd__a211o_2 _10332_ (.A1(_06256_),
    .A2(_03475_),
    .B1(_03476_),
    .C1(_02293_),
    .X(_03477_));
 sky130_fd_sc_hd__o21a_1 _10333_ (.A1(_03339_),
    .A2(_03340_),
    .B1(_03341_),
    .X(_03478_));
 sky130_fd_sc_hd__nor2_1 _10334_ (.A(reg1_val[8]),
    .B(curr_PC[8]),
    .Y(_03479_));
 sky130_fd_sc_hd__nand2_1 _10335_ (.A(reg1_val[8]),
    .B(curr_PC[8]),
    .Y(_03480_));
 sky130_fd_sc_hd__nand2b_1 _10336_ (.A_N(_03479_),
    .B(_03480_),
    .Y(_03481_));
 sky130_fd_sc_hd__xnor2_1 _10337_ (.A(_03478_),
    .B(_03481_),
    .Y(_03482_));
 sky130_fd_sc_hd__mux2_1 _10338_ (.A0(_02248_),
    .A1(_02264_),
    .S(net234),
    .X(_03483_));
 sky130_fd_sc_hd__or2_1 _10339_ (.A(net238),
    .B(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__o21ai_2 _10340_ (.A1(net237),
    .A2(_03363_),
    .B1(_03484_),
    .Y(_03485_));
 sky130_fd_sc_hd__mux2_1 _10341_ (.A0(_03482_),
    .A1(_03485_),
    .S(net242),
    .X(_03486_));
 sky130_fd_sc_hd__o21a_1 _10342_ (.A1(\div_res[7] ),
    .A2(_03353_),
    .B1(net25),
    .X(_03487_));
 sky130_fd_sc_hd__xnor2_1 _10343_ (.A(\div_res[8] ),
    .B(_03487_),
    .Y(_03488_));
 sky130_fd_sc_hd__a21oi_1 _10344_ (.A1(_06255_),
    .A2(_02294_),
    .B1(_02290_),
    .Y(_03489_));
 sky130_fd_sc_hd__or2_1 _10345_ (.A(\div_shifter[39] ),
    .B(_03356_),
    .X(_03490_));
 sky130_fd_sc_hd__a21oi_1 _10346_ (.A1(net247),
    .A2(_03490_),
    .B1(\div_shifter[40] ),
    .Y(_03491_));
 sky130_fd_sc_hd__a31o_1 _10347_ (.A1(\div_shifter[40] ),
    .A2(net247),
    .A3(_03490_),
    .B1(net249),
    .X(_03492_));
 sky130_fd_sc_hd__o2bb2a_1 _10348_ (.A1_N(_06252_),
    .A2_N(net213),
    .B1(_03491_),
    .B2(_03492_),
    .X(_03493_));
 sky130_fd_sc_hd__o221a_1 _10349_ (.A1(_06255_),
    .A2(net204),
    .B1(_03489_),
    .B2(_06254_),
    .C1(_03493_),
    .X(_03494_));
 sky130_fd_sc_hd__o21ai_2 _10350_ (.A1(net239),
    .A2(_03348_),
    .B1(_02312_),
    .Y(_03495_));
 sky130_fd_sc_hd__o221a_1 _10351_ (.A1(net202),
    .A2(_03488_),
    .B1(_03495_),
    .B2(net185),
    .C1(_03494_),
    .X(_03496_));
 sky130_fd_sc_hd__o221a_2 _10352_ (.A1(net183),
    .A2(_03485_),
    .B1(_03486_),
    .B2(_06413_),
    .C1(_03496_),
    .X(_03497_));
 sky130_fd_sc_hd__a41o_1 _10353_ (.A1(_03469_),
    .A2(_03472_),
    .A3(_03477_),
    .A4(_03497_),
    .B1(net262),
    .X(_03498_));
 sky130_fd_sc_hd__and3_2 _10354_ (.A(curr_PC[7]),
    .B(curr_PC[8]),
    .C(_03239_),
    .X(_03499_));
 sky130_fd_sc_hd__a21oi_2 _10355_ (.A1(curr_PC[7]),
    .A2(_03239_),
    .B1(curr_PC[8]),
    .Y(_03500_));
 sky130_fd_sc_hd__o31ai_4 _10356_ (.A1(net257),
    .A2(_03499_),
    .A3(_03500_),
    .B1(_03498_),
    .Y(dest_val[8]));
 sky130_fd_sc_hd__xor2_1 _10357_ (.A(curr_PC[9]),
    .B(_03499_),
    .X(_03501_));
 sky130_fd_sc_hd__a21bo_1 _10358_ (.A1(_03436_),
    .A2(_03445_),
    .B1_N(_03444_),
    .X(_03502_));
 sky130_fd_sc_hd__o2bb2a_1 _10359_ (.A1_N(_06467_),
    .A2_N(_00307_),
    .B1(net47),
    .B2(net100),
    .X(_03503_));
 sky130_fd_sc_hd__xnor2_1 _10360_ (.A(net108),
    .B(_03503_),
    .Y(_03504_));
 sky130_fd_sc_hd__o22a_1 _10361_ (.A1(net76),
    .A2(net41),
    .B1(net39),
    .B2(net73),
    .X(_03505_));
 sky130_fd_sc_hd__xnor2_1 _10362_ (.A(net104),
    .B(_03505_),
    .Y(_03506_));
 sky130_fd_sc_hd__nand2_1 _10363_ (.A(_03504_),
    .B(_03506_),
    .Y(_03507_));
 sky130_fd_sc_hd__xor2_1 _10364_ (.A(_03504_),
    .B(_03506_),
    .X(_03508_));
 sky130_fd_sc_hd__o22a_1 _10365_ (.A1(net118),
    .A2(net50),
    .B1(net48),
    .B2(net70),
    .X(_03509_));
 sky130_fd_sc_hd__xnor2_1 _10366_ (.A(net105),
    .B(_03509_),
    .Y(_03510_));
 sky130_fd_sc_hd__nand2_1 _10367_ (.A(_03508_),
    .B(_03510_),
    .Y(_03511_));
 sky130_fd_sc_hd__or2_1 _10368_ (.A(_03508_),
    .B(_03510_),
    .X(_03512_));
 sky130_fd_sc_hd__and2_1 _10369_ (.A(_03511_),
    .B(_03512_),
    .X(_03513_));
 sky130_fd_sc_hd__nor2_1 _10370_ (.A(net133),
    .B(net31),
    .Y(_03514_));
 sky130_fd_sc_hd__and3_1 _10371_ (.A(_03372_),
    .B(_03374_),
    .C(_03514_),
    .X(_03515_));
 sky130_fd_sc_hd__a21o_1 _10372_ (.A1(_03372_),
    .A2(_03374_),
    .B1(_03514_),
    .X(_03516_));
 sky130_fd_sc_hd__nand2b_1 _10373_ (.A_N(_03515_),
    .B(_03516_),
    .Y(_03517_));
 sky130_fd_sc_hd__xnor2_2 _10374_ (.A(_03398_),
    .B(_03517_),
    .Y(_03518_));
 sky130_fd_sc_hd__nand2_1 _10375_ (.A(_03513_),
    .B(_03518_),
    .Y(_03519_));
 sky130_fd_sc_hd__xor2_1 _10376_ (.A(_03513_),
    .B(_03518_),
    .X(_03520_));
 sky130_fd_sc_hd__o22a_1 _10377_ (.A1(net126),
    .A2(net44),
    .B1(net92),
    .B2(net11),
    .X(_03521_));
 sky130_fd_sc_hd__xnor2_1 _10378_ (.A(net96),
    .B(_03521_),
    .Y(_03522_));
 sky130_fd_sc_hd__o22a_1 _10379_ (.A1(net7),
    .A2(net87),
    .B1(net5),
    .B2(net89),
    .X(_03523_));
 sky130_fd_sc_hd__xnor2_1 _10380_ (.A(net29),
    .B(_03523_),
    .Y(_03524_));
 sky130_fd_sc_hd__o22a_1 _10381_ (.A1(net121),
    .A2(net14),
    .B1(net52),
    .B2(net80),
    .X(_03525_));
 sky130_fd_sc_hd__xor2_1 _10382_ (.A(net111),
    .B(_03525_),
    .X(_03526_));
 sky130_fd_sc_hd__nor2_1 _10383_ (.A(_03524_),
    .B(_03526_),
    .Y(_03527_));
 sky130_fd_sc_hd__xnor2_1 _10384_ (.A(_03524_),
    .B(_03526_),
    .Y(_03528_));
 sky130_fd_sc_hd__nor2_1 _10385_ (.A(_03522_),
    .B(_03528_),
    .Y(_03529_));
 sky130_fd_sc_hd__and2_1 _10386_ (.A(_03522_),
    .B(_03528_),
    .X(_03530_));
 sky130_fd_sc_hd__nor2_1 _10387_ (.A(_03529_),
    .B(_03530_),
    .Y(_03531_));
 sky130_fd_sc_hd__nand2_1 _10388_ (.A(_03520_),
    .B(_03531_),
    .Y(_03532_));
 sky130_fd_sc_hd__or2_1 _10389_ (.A(_03520_),
    .B(_03531_),
    .X(_03533_));
 sky130_fd_sc_hd__a21o_1 _10390_ (.A1(_03427_),
    .A2(_03429_),
    .B1(_03425_),
    .X(_03534_));
 sky130_fd_sc_hd__o22a_1 _10391_ (.A1(net116),
    .A2(net9),
    .B1(net3),
    .B2(net114),
    .X(_03535_));
 sky130_fd_sc_hd__xnor2_1 _10392_ (.A(net179),
    .B(_03535_),
    .Y(_03536_));
 sky130_fd_sc_hd__and3_1 _10393_ (.A(_06445_),
    .B(_00219_),
    .C(_00221_),
    .X(_03537_));
 sky130_fd_sc_hd__a21oi_1 _10394_ (.A1(_00225_),
    .A2(_00226_),
    .B1(net131),
    .Y(_03538_));
 sky130_fd_sc_hd__or3_1 _10395_ (.A(net157),
    .B(_03537_),
    .C(_03538_),
    .X(_03539_));
 sky130_fd_sc_hd__o21ai_1 _10396_ (.A1(_03537_),
    .A2(_03538_),
    .B1(net157),
    .Y(_03540_));
 sky130_fd_sc_hd__a21oi_1 _10397_ (.A1(_03539_),
    .A2(_03540_),
    .B1(_06490_),
    .Y(_03541_));
 sky130_fd_sc_hd__and3_1 _10398_ (.A(_06490_),
    .B(_03539_),
    .C(_03540_),
    .X(_03542_));
 sky130_fd_sc_hd__nor2_1 _10399_ (.A(_03541_),
    .B(_03542_),
    .Y(_03543_));
 sky130_fd_sc_hd__xnor2_1 _10400_ (.A(_03536_),
    .B(_03543_),
    .Y(_03544_));
 sky130_fd_sc_hd__o21ai_1 _10401_ (.A1(_03407_),
    .A2(_03411_),
    .B1(_03544_),
    .Y(_03545_));
 sky130_fd_sc_hd__or3_1 _10402_ (.A(_03407_),
    .B(_03411_),
    .C(_03544_),
    .X(_03546_));
 sky130_fd_sc_hd__and3_1 _10403_ (.A(_03534_),
    .B(_03545_),
    .C(_03546_),
    .X(_03547_));
 sky130_fd_sc_hd__a21oi_1 _10404_ (.A1(_03545_),
    .A2(_03546_),
    .B1(_03534_),
    .Y(_03548_));
 sky130_fd_sc_hd__nor2_1 _10405_ (.A(_03547_),
    .B(_03548_),
    .Y(_03549_));
 sky130_fd_sc_hd__and3_1 _10406_ (.A(_03532_),
    .B(_03533_),
    .C(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__a21o_1 _10407_ (.A1(_03532_),
    .A2(_03533_),
    .B1(_03549_),
    .X(_03551_));
 sky130_fd_sc_hd__nand2b_1 _10408_ (.A_N(_03550_),
    .B(_03551_),
    .Y(_03552_));
 sky130_fd_sc_hd__a21oi_1 _10409_ (.A1(_03392_),
    .A2(_03401_),
    .B1(_03400_),
    .Y(_03553_));
 sky130_fd_sc_hd__o22a_1 _10410_ (.A1(net67),
    .A2(net37),
    .B1(net35),
    .B2(net64),
    .X(_03554_));
 sky130_fd_sc_hd__xnor2_1 _10411_ (.A(net136),
    .B(_03554_),
    .Y(_03555_));
 sky130_fd_sc_hd__o22a_1 _10412_ (.A1(net78),
    .A2(net62),
    .B1(net60),
    .B2(net123),
    .X(_03556_));
 sky130_fd_sc_hd__xnor2_1 _10413_ (.A(net154),
    .B(_03556_),
    .Y(_03557_));
 sky130_fd_sc_hd__and2_1 _10414_ (.A(_03555_),
    .B(_03557_),
    .X(_03558_));
 sky130_fd_sc_hd__nor2_1 _10415_ (.A(_03555_),
    .B(_03557_),
    .Y(_03559_));
 sky130_fd_sc_hd__nor2_1 _10416_ (.A(_03558_),
    .B(_03559_),
    .Y(_03560_));
 sky130_fd_sc_hd__o22a_1 _10417_ (.A1(net57),
    .A2(net42),
    .B1(net94),
    .B2(net54),
    .X(_03561_));
 sky130_fd_sc_hd__xnor2_1 _10418_ (.A(net137),
    .B(_03561_),
    .Y(_03562_));
 sky130_fd_sc_hd__xor2_1 _10419_ (.A(_03560_),
    .B(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__o21ai_1 _10420_ (.A1(_03387_),
    .A2(_03389_),
    .B1(_03563_),
    .Y(_03564_));
 sky130_fd_sc_hd__or3_1 _10421_ (.A(_03387_),
    .B(_03389_),
    .C(_03563_),
    .X(_03565_));
 sky130_fd_sc_hd__and2_1 _10422_ (.A(_03564_),
    .B(_03565_),
    .X(_03566_));
 sky130_fd_sc_hd__nand2b_1 _10423_ (.A_N(_03553_),
    .B(_03566_),
    .Y(_03567_));
 sky130_fd_sc_hd__xnor2_1 _10424_ (.A(_03553_),
    .B(_03566_),
    .Y(_03568_));
 sky130_fd_sc_hd__xnor2_1 _10425_ (.A(_03552_),
    .B(_03568_),
    .Y(_03569_));
 sky130_fd_sc_hd__a21oi_1 _10426_ (.A1(_03418_),
    .A2(_03434_),
    .B1(_03417_),
    .Y(_03570_));
 sky130_fd_sc_hd__a21oi_1 _10427_ (.A1(_03438_),
    .A2(_03442_),
    .B1(_03441_),
    .Y(_03571_));
 sky130_fd_sc_hd__a21bo_1 _10428_ (.A1(_03420_),
    .A2(_03433_),
    .B1_N(_03432_),
    .X(_03572_));
 sky130_fd_sc_hd__or2_1 _10429_ (.A(_03376_),
    .B(_03380_),
    .X(_03573_));
 sky130_fd_sc_hd__a21oi_1 _10430_ (.A1(_03391_),
    .A2(_03415_),
    .B1(_03414_),
    .Y(_03574_));
 sky130_fd_sc_hd__o21bai_1 _10431_ (.A1(_03376_),
    .A2(_03380_),
    .B1_N(_03574_),
    .Y(_03575_));
 sky130_fd_sc_hd__xnor2_1 _10432_ (.A(_03573_),
    .B(_03574_),
    .Y(_03576_));
 sky130_fd_sc_hd__xnor2_1 _10433_ (.A(_03572_),
    .B(_03576_),
    .Y(_03577_));
 sky130_fd_sc_hd__xor2_1 _10434_ (.A(_03571_),
    .B(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__nand2b_1 _10435_ (.A_N(_03570_),
    .B(_03578_),
    .Y(_03579_));
 sky130_fd_sc_hd__xnor2_1 _10436_ (.A(_03570_),
    .B(_03578_),
    .Y(_03580_));
 sky130_fd_sc_hd__and2_1 _10437_ (.A(_03569_),
    .B(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__xnor2_1 _10438_ (.A(_03569_),
    .B(_03580_),
    .Y(_03582_));
 sky130_fd_sc_hd__and2b_1 _10439_ (.A_N(_03582_),
    .B(_03502_),
    .X(_03583_));
 sky130_fd_sc_hd__xor2_1 _10440_ (.A(_03502_),
    .B(_03582_),
    .X(_03584_));
 sky130_fd_sc_hd__a21oi_1 _10441_ (.A1(_03447_),
    .A2(_03449_),
    .B1(_03584_),
    .Y(_03585_));
 sky130_fd_sc_hd__a21o_1 _10442_ (.A1(_03447_),
    .A2(_03449_),
    .B1(_03584_),
    .X(_03586_));
 sky130_fd_sc_hd__and3_1 _10443_ (.A(_03447_),
    .B(_03449_),
    .C(_03584_),
    .X(_03587_));
 sky130_fd_sc_hd__nor2_2 _10444_ (.A(_03585_),
    .B(_03587_),
    .Y(_03588_));
 sky130_fd_sc_hd__and2_1 _10445_ (.A(_03452_),
    .B(_03463_),
    .X(_03589_));
 sky130_fd_sc_hd__xnor2_4 _10446_ (.A(_03588_),
    .B(_03589_),
    .Y(_03590_));
 sky130_fd_sc_hd__or4b_2 _10447_ (.A(_03199_),
    .B(_03329_),
    .C(_03466_),
    .D_N(_03464_),
    .X(_03591_));
 sky130_fd_sc_hd__a21o_1 _10448_ (.A1(net19),
    .A2(_03591_),
    .B1(_03590_),
    .X(_03592_));
 sky130_fd_sc_hd__nand3_1 _10449_ (.A(net19),
    .B(_03590_),
    .C(_03591_),
    .Y(_03593_));
 sky130_fd_sc_hd__and3_1 _10450_ (.A(net206),
    .B(_03592_),
    .C(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__o21ai_1 _10451_ (.A1(net84),
    .A2(_02174_),
    .B1(_02158_),
    .Y(_03595_));
 sky130_fd_sc_hd__o311a_1 _10452_ (.A1(net84),
    .A2(_02158_),
    .A3(_02174_),
    .B1(_02298_),
    .C1(_03595_),
    .X(_03596_));
 sky130_fd_sc_hd__o21a_1 _10453_ (.A1(_06254_),
    .A2(_03474_),
    .B1(_06255_),
    .X(_03597_));
 sky130_fd_sc_hd__mux2_1 _10454_ (.A0(_06319_),
    .A1(_03597_),
    .S(net299),
    .X(_03598_));
 sky130_fd_sc_hd__a21oi_1 _10455_ (.A1(_06250_),
    .A2(_03598_),
    .B1(_02293_),
    .Y(_03599_));
 sky130_fd_sc_hd__o21a_1 _10456_ (.A1(_06250_),
    .A2(_03598_),
    .B1(_03599_),
    .X(_03600_));
 sky130_fd_sc_hd__o21a_1 _10457_ (.A1(_03478_),
    .A2(_03479_),
    .B1(_03480_),
    .X(_03601_));
 sky130_fd_sc_hd__nor2_1 _10458_ (.A(reg1_val[9]),
    .B(curr_PC[9]),
    .Y(_03602_));
 sky130_fd_sc_hd__nand2_1 _10459_ (.A(reg1_val[9]),
    .B(curr_PC[9]),
    .Y(_03603_));
 sky130_fd_sc_hd__and2b_1 _10460_ (.A_N(_03602_),
    .B(_03603_),
    .X(_03604_));
 sky130_fd_sc_hd__xnor2_1 _10461_ (.A(_03601_),
    .B(_03604_),
    .Y(_03605_));
 sky130_fd_sc_hd__mux2_1 _10462_ (.A0(_02459_),
    .A1(_02467_),
    .S(net236),
    .X(_03606_));
 sky130_fd_sc_hd__mux2_1 _10463_ (.A0(_03234_),
    .A1(_03606_),
    .S(net237),
    .X(_03607_));
 sky130_fd_sc_hd__mux2_1 _10464_ (.A0(_03605_),
    .A1(_03607_),
    .S(net241),
    .X(_03608_));
 sky130_fd_sc_hd__or3_1 _10465_ (.A(\div_res[8] ),
    .B(\div_res[7] ),
    .C(_03353_),
    .X(_03609_));
 sky130_fd_sc_hd__a21oi_1 _10466_ (.A1(net25),
    .A2(_03609_),
    .B1(\div_res[9] ),
    .Y(_03610_));
 sky130_fd_sc_hd__a31o_1 _10467_ (.A1(\div_res[9] ),
    .A2(net25),
    .A3(_03609_),
    .B1(net202),
    .X(_03611_));
 sky130_fd_sc_hd__a21oi_1 _10468_ (.A1(_06249_),
    .A2(_02294_),
    .B1(net205),
    .Y(_03612_));
 sky130_fd_sc_hd__or3_2 _10469_ (.A(\div_shifter[40] ),
    .B(\div_shifter[39] ),
    .C(_03356_),
    .X(_03613_));
 sky130_fd_sc_hd__a21oi_2 _10470_ (.A1(net246),
    .A2(_03613_),
    .B1(\div_shifter[41] ),
    .Y(_03614_));
 sky130_fd_sc_hd__a31o_1 _10471_ (.A1(\div_shifter[41] ),
    .A2(net246),
    .A3(_03613_),
    .B1(net249),
    .X(_03615_));
 sky130_fd_sc_hd__o221a_1 _10472_ (.A1(_06246_),
    .A2(_06426_),
    .B1(net204),
    .B2(_06249_),
    .C1(net261),
    .X(_03616_));
 sky130_fd_sc_hd__o221a_1 _10473_ (.A1(_06248_),
    .A2(_03612_),
    .B1(_03614_),
    .B2(_03615_),
    .C1(_03616_),
    .X(_03617_));
 sky130_fd_sc_hd__o21ai_1 _10474_ (.A1(_03610_),
    .A2(_03611_),
    .B1(_03617_),
    .Y(_03618_));
 sky130_fd_sc_hd__o21ai_1 _10475_ (.A1(net238),
    .A2(_03221_),
    .B1(_02312_),
    .Y(_03619_));
 sky130_fd_sc_hd__inv_2 _10476_ (.A(_03619_),
    .Y(_03620_));
 sky130_fd_sc_hd__a221o_1 _10477_ (.A1(_02288_),
    .A2(_03607_),
    .B1(_03620_),
    .B2(_02217_),
    .C1(_03618_),
    .X(_03621_));
 sky130_fd_sc_hd__a211o_2 _10478_ (.A1(net215),
    .A2(_03608_),
    .B1(_03621_),
    .C1(_03600_),
    .X(_03622_));
 sky130_fd_sc_hd__o32a_4 _10479_ (.A1(_03594_),
    .A2(_03596_),
    .A3(_03622_),
    .B1(_03501_),
    .B2(net257),
    .X(dest_val[9]));
 sky130_fd_sc_hd__o21ai_1 _10480_ (.A1(_03571_),
    .A2(_03577_),
    .B1(_03579_),
    .Y(_03623_));
 sky130_fd_sc_hd__nor2_1 _10481_ (.A(net116),
    .B(net3),
    .Y(_03624_));
 sky130_fd_sc_hd__xnor2_2 _10482_ (.A(net179),
    .B(_03624_),
    .Y(_03625_));
 sky130_fd_sc_hd__a21oi_1 _10483_ (.A1(_03507_),
    .A2(_03511_),
    .B1(_03625_),
    .Y(_03626_));
 sky130_fd_sc_hd__and3_1 _10484_ (.A(_03507_),
    .B(_03511_),
    .C(_03625_),
    .X(_03627_));
 sky130_fd_sc_hd__or2_1 _10485_ (.A(_03626_),
    .B(_03627_),
    .X(_03628_));
 sky130_fd_sc_hd__a21oi_1 _10486_ (.A1(_03560_),
    .A2(_03562_),
    .B1(_03558_),
    .Y(_03629_));
 sky130_fd_sc_hd__nor2_1 _10487_ (.A(_03628_),
    .B(_03629_),
    .Y(_03630_));
 sky130_fd_sc_hd__and2_1 _10488_ (.A(_03628_),
    .B(_03629_),
    .X(_03631_));
 sky130_fd_sc_hd__nor2_1 _10489_ (.A(_03630_),
    .B(_03631_),
    .Y(_03632_));
 sky130_fd_sc_hd__o22a_1 _10490_ (.A1(net125),
    .A2(net11),
    .B1(net44),
    .B2(net121),
    .X(_03633_));
 sky130_fd_sc_hd__xnor2_1 _10491_ (.A(net96),
    .B(_03633_),
    .Y(_03634_));
 sky130_fd_sc_hd__o22a_1 _10492_ (.A1(net118),
    .A2(net47),
    .B1(net99),
    .B2(net13),
    .X(_03635_));
 sky130_fd_sc_hd__xnor2_1 _10493_ (.A(net108),
    .B(_03635_),
    .Y(_03636_));
 sky130_fd_sc_hd__nand2b_1 _10494_ (.A_N(_03634_),
    .B(_03636_),
    .Y(_03637_));
 sky130_fd_sc_hd__nand2b_1 _10495_ (.A_N(_03636_),
    .B(_03634_),
    .Y(_03638_));
 sky130_fd_sc_hd__nand2_1 _10496_ (.A(_03637_),
    .B(_03638_),
    .Y(_03639_));
 sky130_fd_sc_hd__o22a_1 _10497_ (.A1(net81),
    .A2(net14),
    .B1(net52),
    .B2(net129),
    .X(_03640_));
 sky130_fd_sc_hd__xnor2_1 _10498_ (.A(net111),
    .B(_03640_),
    .Y(_03641_));
 sky130_fd_sc_hd__inv_2 _10499_ (.A(_03641_),
    .Y(_03642_));
 sky130_fd_sc_hd__xnor2_1 _10500_ (.A(_03639_),
    .B(_03642_),
    .Y(_03643_));
 sky130_fd_sc_hd__o21ba_1 _10501_ (.A1(_03536_),
    .A2(_03542_),
    .B1_N(_03541_),
    .X(_03644_));
 sky130_fd_sc_hd__o22a_1 _10502_ (.A1(net7),
    .A2(net93),
    .B1(net87),
    .B2(net5),
    .X(_03645_));
 sky130_fd_sc_hd__xnor2_1 _10503_ (.A(net28),
    .B(_03645_),
    .Y(_03646_));
 sky130_fd_sc_hd__xnor2_1 _10504_ (.A(_03644_),
    .B(_03646_),
    .Y(_03647_));
 sky130_fd_sc_hd__nor2_1 _10505_ (.A(net89),
    .B(net28),
    .Y(_03648_));
 sky130_fd_sc_hd__or3_1 _10506_ (.A(net89),
    .B(net28),
    .C(_03647_),
    .X(_03649_));
 sky130_fd_sc_hd__xnor2_1 _10507_ (.A(_03647_),
    .B(_03648_),
    .Y(_03650_));
 sky130_fd_sc_hd__o22a_1 _10508_ (.A1(net70),
    .A2(net50),
    .B1(net48),
    .B2(net76),
    .X(_03651_));
 sky130_fd_sc_hd__xnor2_1 _10509_ (.A(net105),
    .B(_03651_),
    .Y(_03652_));
 sky130_fd_sc_hd__o22a_1 _10510_ (.A1(net64),
    .A2(net37),
    .B1(net35),
    .B2(net57),
    .X(_03653_));
 sky130_fd_sc_hd__xnor2_1 _10511_ (.A(net136),
    .B(_03653_),
    .Y(_03654_));
 sky130_fd_sc_hd__and2_1 _10512_ (.A(_03652_),
    .B(_03654_),
    .X(_03655_));
 sky130_fd_sc_hd__nor2_1 _10513_ (.A(_03652_),
    .B(_03654_),
    .Y(_03656_));
 sky130_fd_sc_hd__nor2_1 _10514_ (.A(_03655_),
    .B(_03656_),
    .Y(_03657_));
 sky130_fd_sc_hd__o22a_1 _10515_ (.A1(net73),
    .A2(net41),
    .B1(net39),
    .B2(net67),
    .X(_03658_));
 sky130_fd_sc_hd__xnor2_1 _10516_ (.A(net104),
    .B(_03658_),
    .Y(_03659_));
 sky130_fd_sc_hd__xor2_1 _10517_ (.A(_03657_),
    .B(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__nand2_1 _10518_ (.A(_03650_),
    .B(_03660_),
    .Y(_03661_));
 sky130_fd_sc_hd__xnor2_1 _10519_ (.A(_03650_),
    .B(_03660_),
    .Y(_03662_));
 sky130_fd_sc_hd__xor2_1 _10520_ (.A(_03643_),
    .B(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__and2_1 _10521_ (.A(_03632_),
    .B(_03663_),
    .X(_03664_));
 sky130_fd_sc_hd__nor2_1 _10522_ (.A(_03632_),
    .B(_03663_),
    .Y(_03665_));
 sky130_fd_sc_hd__nor2_1 _10523_ (.A(_03664_),
    .B(_03665_),
    .Y(_03666_));
 sky130_fd_sc_hd__a21oi_2 _10524_ (.A1(_03398_),
    .A2(_03516_),
    .B1(_03515_),
    .Y(_03667_));
 sky130_fd_sc_hd__o22a_1 _10525_ (.A1(net54),
    .A2(net43),
    .B1(net95),
    .B2(net62),
    .X(_03668_));
 sky130_fd_sc_hd__xnor2_1 _10526_ (.A(net139),
    .B(_03668_),
    .Y(_03669_));
 sky130_fd_sc_hd__inv_2 _10527_ (.A(_03669_),
    .Y(_03670_));
 sky130_fd_sc_hd__o22a_1 _10528_ (.A1(net82),
    .A2(net16),
    .B1(net9),
    .B2(net131),
    .X(_03671_));
 sky130_fd_sc_hd__xnor2_1 _10529_ (.A(net157),
    .B(_03671_),
    .Y(_03672_));
 sky130_fd_sc_hd__nor2_1 _10530_ (.A(_03670_),
    .B(_03672_),
    .Y(_03673_));
 sky130_fd_sc_hd__and2_1 _10531_ (.A(_03670_),
    .B(_03672_),
    .X(_03674_));
 sky130_fd_sc_hd__nor2_1 _10532_ (.A(_03673_),
    .B(_03674_),
    .Y(_03675_));
 sky130_fd_sc_hd__o22a_1 _10533_ (.A1(net78),
    .A2(net60),
    .B1(net18),
    .B2(net123),
    .X(_03676_));
 sky130_fd_sc_hd__xnor2_1 _10534_ (.A(net154),
    .B(_03676_),
    .Y(_03677_));
 sky130_fd_sc_hd__xor2_1 _10535_ (.A(_03675_),
    .B(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__o21a_1 _10536_ (.A1(_03527_),
    .A2(_03529_),
    .B1(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__nor3_1 _10537_ (.A(_03527_),
    .B(_03529_),
    .C(_03678_),
    .Y(_03680_));
 sky130_fd_sc_hd__nor2_1 _10538_ (.A(_03679_),
    .B(_03680_),
    .Y(_03681_));
 sky130_fd_sc_hd__xnor2_1 _10539_ (.A(_03667_),
    .B(_03681_),
    .Y(_03682_));
 sky130_fd_sc_hd__xor2_1 _10540_ (.A(_03666_),
    .B(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__a21oi_1 _10541_ (.A1(_03551_),
    .A2(_03568_),
    .B1(_03550_),
    .Y(_03684_));
 sky130_fd_sc_hd__nand2_1 _10542_ (.A(_03564_),
    .B(_03567_),
    .Y(_03685_));
 sky130_fd_sc_hd__a21boi_1 _10543_ (.A1(_03534_),
    .A2(_03546_),
    .B1_N(_03545_),
    .Y(_03686_));
 sky130_fd_sc_hd__a21oi_1 _10544_ (.A1(_03519_),
    .A2(_03532_),
    .B1(_03686_),
    .Y(_03687_));
 sky130_fd_sc_hd__and3_1 _10545_ (.A(_03519_),
    .B(_03532_),
    .C(_03686_),
    .X(_03688_));
 sky130_fd_sc_hd__nor2_1 _10546_ (.A(_03687_),
    .B(_03688_),
    .Y(_03689_));
 sky130_fd_sc_hd__xnor2_1 _10547_ (.A(_03685_),
    .B(_03689_),
    .Y(_03690_));
 sky130_fd_sc_hd__a21bo_1 _10548_ (.A1(_03572_),
    .A2(_03576_),
    .B1_N(_03575_),
    .X(_03691_));
 sky130_fd_sc_hd__nand2b_1 _10549_ (.A_N(_03690_),
    .B(_03691_),
    .Y(_03692_));
 sky130_fd_sc_hd__xnor2_1 _10550_ (.A(_03690_),
    .B(_03691_),
    .Y(_03693_));
 sky130_fd_sc_hd__nand2b_1 _10551_ (.A_N(_03684_),
    .B(_03693_),
    .Y(_03694_));
 sky130_fd_sc_hd__xnor2_1 _10552_ (.A(_03684_),
    .B(_03693_),
    .Y(_03695_));
 sky130_fd_sc_hd__and2_1 _10553_ (.A(_03683_),
    .B(_03695_),
    .X(_03696_));
 sky130_fd_sc_hd__xor2_1 _10554_ (.A(_03683_),
    .B(_03695_),
    .X(_03697_));
 sky130_fd_sc_hd__xor2_1 _10555_ (.A(_03623_),
    .B(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__o21a_1 _10556_ (.A1(_03581_),
    .A2(_03583_),
    .B1(_03698_),
    .X(_03699_));
 sky130_fd_sc_hd__nor3_1 _10557_ (.A(_03581_),
    .B(_03583_),
    .C(_03698_),
    .Y(_03700_));
 sky130_fd_sc_hd__nor2_2 _10558_ (.A(_03699_),
    .B(_03700_),
    .Y(_03701_));
 sky130_fd_sc_hd__a21oi_1 _10559_ (.A1(_03452_),
    .A2(_03586_),
    .B1(_03587_),
    .Y(_03702_));
 sky130_fd_sc_hd__and2b_1 _10560_ (.A_N(_03453_),
    .B(_03588_),
    .X(_03703_));
 sky130_fd_sc_hd__a21o_2 _10561_ (.A1(_03462_),
    .A2(_03703_),
    .B1(_03702_),
    .X(_03704_));
 sky130_fd_sc_hd__xor2_4 _10562_ (.A(_03701_),
    .B(_03704_),
    .X(_03705_));
 sky130_fd_sc_hd__o21a_1 _10563_ (.A1(_03590_),
    .A2(_03591_),
    .B1(net19),
    .X(_03706_));
 sky130_fd_sc_hd__a21oi_1 _10564_ (.A1(_03705_),
    .A2(_03706_),
    .B1(_02214_),
    .Y(_03707_));
 sky130_fd_sc_hd__o21ai_1 _10565_ (.A1(_03705_),
    .A2(_03706_),
    .B1(_03707_),
    .Y(_03708_));
 sky130_fd_sc_hd__a21oi_1 _10566_ (.A1(net19),
    .A2(_02175_),
    .B1(_02157_),
    .Y(_03709_));
 sky130_fd_sc_hd__a31o_1 _10567_ (.A1(net19),
    .A2(_02157_),
    .A3(_02175_),
    .B1(net250),
    .X(_03710_));
 sky130_fd_sc_hd__o21a_1 _10568_ (.A1(_06248_),
    .A2(_03597_),
    .B1(_06249_),
    .X(_03711_));
 sky130_fd_sc_hd__mux2_1 _10569_ (.A0(_06321_),
    .A1(_03711_),
    .S(net299),
    .X(_03712_));
 sky130_fd_sc_hd__nor2_1 _10570_ (.A(_06243_),
    .B(_03712_),
    .Y(_03713_));
 sky130_fd_sc_hd__a211o_1 _10571_ (.A1(_06243_),
    .A2(_03712_),
    .B1(_03713_),
    .C1(_02293_),
    .X(_03714_));
 sky130_fd_sc_hd__nor2_1 _10572_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .Y(_03715_));
 sky130_fd_sc_hd__and2_1 _10573_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .X(_03716_));
 sky130_fd_sc_hd__nand2_1 _10574_ (.A(reg1_val[10]),
    .B(curr_PC[10]),
    .Y(_03717_));
 sky130_fd_sc_hd__o21a_1 _10575_ (.A1(_03601_),
    .A2(_03602_),
    .B1(_03603_),
    .X(_03718_));
 sky130_fd_sc_hd__o21a_1 _10576_ (.A1(_03715_),
    .A2(_03716_),
    .B1(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__or3_1 _10577_ (.A(_03715_),
    .B(_03716_),
    .C(_03718_),
    .X(_03720_));
 sky130_fd_sc_hd__nand2_1 _10578_ (.A(net263),
    .B(_03720_),
    .Y(_03721_));
 sky130_fd_sc_hd__mux2_1 _10579_ (.A0(_02631_),
    .A1(_02635_),
    .S(net234),
    .X(_03722_));
 sky130_fd_sc_hd__inv_2 _10580_ (.A(_03722_),
    .Y(_03723_));
 sky130_fd_sc_hd__mux2_1 _10581_ (.A0(_03099_),
    .A1(_03723_),
    .S(net237),
    .X(_03724_));
 sky130_fd_sc_hd__o22a_1 _10582_ (.A1(_03719_),
    .A2(_03721_),
    .B1(_03724_),
    .B2(net263),
    .X(_03725_));
 sky130_fd_sc_hd__or2_1 _10583_ (.A(\div_res[9] ),
    .B(_03609_),
    .X(_03726_));
 sky130_fd_sc_hd__a21oi_1 _10584_ (.A1(net23),
    .A2(_03726_),
    .B1(\div_res[10] ),
    .Y(_03727_));
 sky130_fd_sc_hd__a31o_1 _10585_ (.A1(\div_res[10] ),
    .A2(net23),
    .A3(_03726_),
    .B1(net202),
    .X(_03728_));
 sky130_fd_sc_hd__mux2_1 _10586_ (.A0(_02300_),
    .A1(_02294_),
    .S(_06241_),
    .X(_03729_));
 sky130_fd_sc_hd__o21ai_1 _10587_ (.A1(net205),
    .A2(_03729_),
    .B1(_06242_),
    .Y(_03730_));
 sky130_fd_sc_hd__or2_1 _10588_ (.A(\div_shifter[41] ),
    .B(_03613_),
    .X(_03731_));
 sky130_fd_sc_hd__a21oi_1 _10589_ (.A1(net246),
    .A2(_03731_),
    .B1(\div_shifter[42] ),
    .Y(_03732_));
 sky130_fd_sc_hd__a31o_1 _10590_ (.A1(\div_shifter[42] ),
    .A2(net246),
    .A3(_03731_),
    .B1(net249),
    .X(_03733_));
 sky130_fd_sc_hd__o2bb2a_1 _10591_ (.A1_N(_06233_),
    .A2_N(net213),
    .B1(_03732_),
    .B2(_03733_),
    .X(_03734_));
 sky130_fd_sc_hd__o211a_1 _10592_ (.A1(_03727_),
    .A2(_03728_),
    .B1(_03730_),
    .C1(_03734_),
    .X(_03735_));
 sky130_fd_sc_hd__a21o_1 _10593_ (.A1(net237),
    .A2(_03087_),
    .B1(_02311_),
    .X(_03736_));
 sky130_fd_sc_hd__o221a_1 _10594_ (.A1(net183),
    .A2(_03724_),
    .B1(_03736_),
    .B2(net185),
    .C1(_03735_),
    .X(_03737_));
 sky130_fd_sc_hd__o211a_1 _10595_ (.A1(net214),
    .A2(_03725_),
    .B1(_03737_),
    .C1(_03714_),
    .X(_03738_));
 sky130_fd_sc_hd__o211a_1 _10596_ (.A1(_03709_),
    .A2(_03710_),
    .B1(_03738_),
    .C1(_03708_),
    .X(_03739_));
 sky130_fd_sc_hd__and3_1 _10597_ (.A(curr_PC[9]),
    .B(curr_PC[10]),
    .C(_03499_),
    .X(_03740_));
 sky130_fd_sc_hd__a21oi_1 _10598_ (.A1(curr_PC[9]),
    .A2(_03499_),
    .B1(curr_PC[10]),
    .Y(_03741_));
 sky130_fd_sc_hd__or3_1 _10599_ (.A(net257),
    .B(_03740_),
    .C(_03741_),
    .X(_03742_));
 sky130_fd_sc_hd__o21ai_4 _10600_ (.A1(net262),
    .A2(_03739_),
    .B1(_03742_),
    .Y(dest_val[10]));
 sky130_fd_sc_hd__a21oi_1 _10601_ (.A1(_03623_),
    .A2(_03697_),
    .B1(_03696_),
    .Y(_03743_));
 sky130_fd_sc_hd__nand2_1 _10602_ (.A(_03692_),
    .B(_03694_),
    .Y(_03744_));
 sky130_fd_sc_hd__o21ai_2 _10603_ (.A1(_03644_),
    .A2(_03646_),
    .B1(_03649_),
    .Y(_03745_));
 sky130_fd_sc_hd__o22a_1 _10604_ (.A1(net78),
    .A2(net18),
    .B1(net16),
    .B2(net123),
    .X(_03746_));
 sky130_fd_sc_hd__xnor2_1 _10605_ (.A(net154),
    .B(_03746_),
    .Y(_03747_));
 sky130_fd_sc_hd__nand2_1 _10606_ (.A(net179),
    .B(_03747_),
    .Y(_03748_));
 sky130_fd_sc_hd__xor2_1 _10607_ (.A(net179),
    .B(_03747_),
    .X(_03749_));
 sky130_fd_sc_hd__o22a_1 _10608_ (.A1(net82),
    .A2(net9),
    .B1(net3),
    .B2(net131),
    .X(_03750_));
 sky130_fd_sc_hd__xnor2_2 _10609_ (.A(_06435_),
    .B(_03750_),
    .Y(_03751_));
 sky130_fd_sc_hd__nand2_1 _10610_ (.A(_03749_),
    .B(_03751_),
    .Y(_03752_));
 sky130_fd_sc_hd__or2_1 _10611_ (.A(_03749_),
    .B(_03751_),
    .X(_03753_));
 sky130_fd_sc_hd__and2_1 _10612_ (.A(_03752_),
    .B(_03753_),
    .X(_03754_));
 sky130_fd_sc_hd__o21ai_1 _10613_ (.A1(_03639_),
    .A2(_03642_),
    .B1(_03637_),
    .Y(_03755_));
 sky130_fd_sc_hd__and2_1 _10614_ (.A(_03754_),
    .B(_03755_),
    .X(_03756_));
 sky130_fd_sc_hd__nor2_1 _10615_ (.A(_03754_),
    .B(_03755_),
    .Y(_03757_));
 sky130_fd_sc_hd__nor2_1 _10616_ (.A(_03756_),
    .B(_03757_),
    .Y(_03758_));
 sky130_fd_sc_hd__xnor2_2 _10617_ (.A(_03745_),
    .B(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__a21o_1 _10618_ (.A1(_03675_),
    .A2(_03677_),
    .B1(_03673_),
    .X(_03760_));
 sky130_fd_sc_hd__a21o_1 _10619_ (.A1(_03657_),
    .A2(_03659_),
    .B1(_03655_),
    .X(_03761_));
 sky130_fd_sc_hd__and2_1 _10620_ (.A(_03625_),
    .B(_03761_),
    .X(_03762_));
 sky130_fd_sc_hd__xor2_2 _10621_ (.A(_03625_),
    .B(_03761_),
    .X(_03763_));
 sky130_fd_sc_hd__xnor2_2 _10622_ (.A(_03760_),
    .B(_03763_),
    .Y(_03764_));
 sky130_fd_sc_hd__o22a_1 _10623_ (.A1(net129),
    .A2(net14),
    .B1(net52),
    .B2(net99),
    .X(_03765_));
 sky130_fd_sc_hd__xor2_1 _10624_ (.A(net111),
    .B(_03765_),
    .X(_03766_));
 sky130_fd_sc_hd__o22a_1 _10625_ (.A1(net76),
    .A2(net50),
    .B1(net48),
    .B2(net73),
    .X(_03767_));
 sky130_fd_sc_hd__xor2_1 _10626_ (.A(net105),
    .B(_03767_),
    .X(_03768_));
 sky130_fd_sc_hd__nor2_1 _10627_ (.A(_03766_),
    .B(_03768_),
    .Y(_03769_));
 sky130_fd_sc_hd__xor2_1 _10628_ (.A(_03766_),
    .B(_03768_),
    .X(_03770_));
 sky130_fd_sc_hd__o22a_1 _10629_ (.A1(net118),
    .A2(net13),
    .B1(net47),
    .B2(net70),
    .X(_03771_));
 sky130_fd_sc_hd__xnor2_1 _10630_ (.A(net108),
    .B(_03771_),
    .Y(_03772_));
 sky130_fd_sc_hd__and2_1 _10631_ (.A(_03770_),
    .B(_03772_),
    .X(_03773_));
 sky130_fd_sc_hd__nor2_1 _10632_ (.A(_03770_),
    .B(_03772_),
    .Y(_03774_));
 sky130_fd_sc_hd__or2_1 _10633_ (.A(_03773_),
    .B(_03774_),
    .X(_03775_));
 sky130_fd_sc_hd__o22a_1 _10634_ (.A1(net62),
    .A2(net43),
    .B1(net95),
    .B2(net60),
    .X(_03776_));
 sky130_fd_sc_hd__xnor2_1 _10635_ (.A(net139),
    .B(_03776_),
    .Y(_03777_));
 sky130_fd_sc_hd__o22a_1 _10636_ (.A1(net67),
    .A2(net41),
    .B1(net39),
    .B2(net64),
    .X(_03778_));
 sky130_fd_sc_hd__xnor2_1 _10637_ (.A(net104),
    .B(_03778_),
    .Y(_03779_));
 sky130_fd_sc_hd__and2_1 _10638_ (.A(_03777_),
    .B(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__xor2_1 _10639_ (.A(_03777_),
    .B(_03779_),
    .X(_03781_));
 sky130_fd_sc_hd__o22a_1 _10640_ (.A1(net57),
    .A2(net37),
    .B1(net35),
    .B2(net54),
    .X(_03782_));
 sky130_fd_sc_hd__xnor2_1 _10641_ (.A(net136),
    .B(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__and2_1 _10642_ (.A(_03781_),
    .B(_03783_),
    .X(_03784_));
 sky130_fd_sc_hd__nor2_1 _10643_ (.A(_03781_),
    .B(_03783_),
    .Y(_03785_));
 sky130_fd_sc_hd__nor2_1 _10644_ (.A(_03784_),
    .B(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__o22a_1 _10645_ (.A1(net125),
    .A2(net7),
    .B1(net93),
    .B2(net5),
    .X(_03787_));
 sky130_fd_sc_hd__xnor2_1 _10646_ (.A(net28),
    .B(_03787_),
    .Y(_03788_));
 sky130_fd_sc_hd__nor2_1 _10647_ (.A(net87),
    .B(net28),
    .Y(_03789_));
 sky130_fd_sc_hd__o22a_1 _10648_ (.A1(net122),
    .A2(net11),
    .B1(net44),
    .B2(net81),
    .X(_03790_));
 sky130_fd_sc_hd__xor2_1 _10649_ (.A(net96),
    .B(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__nand2_1 _10650_ (.A(_03789_),
    .B(_03791_),
    .Y(_03792_));
 sky130_fd_sc_hd__xnor2_1 _10651_ (.A(_03789_),
    .B(_03791_),
    .Y(_03793_));
 sky130_fd_sc_hd__xor2_1 _10652_ (.A(_03788_),
    .B(_03793_),
    .X(_03794_));
 sky130_fd_sc_hd__and2_1 _10653_ (.A(_03786_),
    .B(_03794_),
    .X(_03795_));
 sky130_fd_sc_hd__xnor2_1 _10654_ (.A(_03786_),
    .B(_03794_),
    .Y(_03796_));
 sky130_fd_sc_hd__nor2_1 _10655_ (.A(_03775_),
    .B(_03796_),
    .Y(_03797_));
 sky130_fd_sc_hd__and2_1 _10656_ (.A(_03775_),
    .B(_03796_),
    .X(_03798_));
 sky130_fd_sc_hd__or2_1 _10657_ (.A(_03797_),
    .B(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__xor2_2 _10658_ (.A(_03764_),
    .B(_03799_),
    .X(_03800_));
 sky130_fd_sc_hd__and2b_1 _10659_ (.A_N(_03759_),
    .B(_03800_),
    .X(_03801_));
 sky130_fd_sc_hd__xnor2_2 _10660_ (.A(_03759_),
    .B(_03800_),
    .Y(_03802_));
 sky130_fd_sc_hd__a21o_1 _10661_ (.A1(_03666_),
    .A2(_03682_),
    .B1(_03664_),
    .X(_03803_));
 sky130_fd_sc_hd__o21bai_2 _10662_ (.A1(_03667_),
    .A2(_03680_),
    .B1_N(_03679_),
    .Y(_03804_));
 sky130_fd_sc_hd__or2_1 _10663_ (.A(_03626_),
    .B(_03630_),
    .X(_03805_));
 sky130_fd_sc_hd__o21a_1 _10664_ (.A1(_03643_),
    .A2(_03662_),
    .B1(_03661_),
    .X(_03806_));
 sky130_fd_sc_hd__o21bai_1 _10665_ (.A1(_03626_),
    .A2(_03630_),
    .B1_N(_03806_),
    .Y(_03807_));
 sky130_fd_sc_hd__xnor2_2 _10666_ (.A(_03805_),
    .B(_03806_),
    .Y(_03808_));
 sky130_fd_sc_hd__xnor2_2 _10667_ (.A(_03804_),
    .B(_03808_),
    .Y(_03809_));
 sky130_fd_sc_hd__a21oi_2 _10668_ (.A1(_03685_),
    .A2(_03689_),
    .B1(_03687_),
    .Y(_03810_));
 sky130_fd_sc_hd__xnor2_2 _10669_ (.A(_03809_),
    .B(_03810_),
    .Y(_03811_));
 sky130_fd_sc_hd__nand2b_1 _10670_ (.A_N(_03811_),
    .B(_03803_),
    .Y(_03812_));
 sky130_fd_sc_hd__xnor2_2 _10671_ (.A(_03803_),
    .B(_03811_),
    .Y(_03813_));
 sky130_fd_sc_hd__and2_1 _10672_ (.A(_03802_),
    .B(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__xor2_2 _10673_ (.A(_03802_),
    .B(_03813_),
    .X(_03815_));
 sky130_fd_sc_hd__xnor2_1 _10674_ (.A(_03744_),
    .B(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hd__and2_1 _10675_ (.A(_03743_),
    .B(_03816_),
    .X(_03817_));
 sky130_fd_sc_hd__nor2_1 _10676_ (.A(_03743_),
    .B(_03816_),
    .Y(_03818_));
 sky130_fd_sc_hd__or2_2 _10677_ (.A(_03817_),
    .B(_03818_),
    .X(_03819_));
 sky130_fd_sc_hd__inv_2 _10678_ (.A(_03819_),
    .Y(_03820_));
 sky130_fd_sc_hd__a21oi_2 _10679_ (.A1(_03701_),
    .A2(_03704_),
    .B1(_03699_),
    .Y(_03821_));
 sky130_fd_sc_hd__xnor2_4 _10680_ (.A(_03819_),
    .B(_03821_),
    .Y(_03822_));
 sky130_fd_sc_hd__nor2_1 _10681_ (.A(_03590_),
    .B(_03705_),
    .Y(_03823_));
 sky130_fd_sc_hd__and2b_1 _10682_ (.A_N(_03591_),
    .B(_03823_),
    .X(_03824_));
 sky130_fd_sc_hd__or2_1 _10683_ (.A(net84),
    .B(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__nor2_1 _10684_ (.A(_03822_),
    .B(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__a21o_1 _10685_ (.A1(_03822_),
    .A2(_03825_),
    .B1(_02214_),
    .X(_03827_));
 sky130_fd_sc_hd__a21oi_1 _10686_ (.A1(net19),
    .A2(_02176_),
    .B1(_02178_),
    .Y(_03828_));
 sky130_fd_sc_hd__a31o_1 _10687_ (.A1(net19),
    .A2(_02176_),
    .A3(_02178_),
    .B1(net250),
    .X(_03829_));
 sky130_fd_sc_hd__or2_1 _10688_ (.A(_03828_),
    .B(_03829_),
    .X(_03830_));
 sky130_fd_sc_hd__and3_1 _10689_ (.A(net305),
    .B(_06240_),
    .C(_06322_),
    .X(_03831_));
 sky130_fd_sc_hd__o21a_1 _10690_ (.A1(_06243_),
    .A2(_03711_),
    .B1(_06241_),
    .X(_03832_));
 sky130_fd_sc_hd__o21ba_1 _10691_ (.A1(net305),
    .A2(_03832_),
    .B1_N(_03831_),
    .X(_03833_));
 sky130_fd_sc_hd__nor2_1 _10692_ (.A(_06216_),
    .B(_03833_),
    .Y(_03834_));
 sky130_fd_sc_hd__a211o_1 _10693_ (.A1(_06216_),
    .A2(_03833_),
    .B1(_03834_),
    .C1(_02293_),
    .X(_03835_));
 sky130_fd_sc_hd__nor2_1 _10694_ (.A(reg1_val[11]),
    .B(curr_PC[11]),
    .Y(_03836_));
 sky130_fd_sc_hd__and2_1 _10695_ (.A(reg1_val[11]),
    .B(curr_PC[11]),
    .X(_03837_));
 sky130_fd_sc_hd__o211a_1 _10696_ (.A1(_03836_),
    .A2(_03837_),
    .B1(_03717_),
    .C1(_03720_),
    .X(_03838_));
 sky130_fd_sc_hd__a211oi_2 _10697_ (.A1(_03717_),
    .A2(_03720_),
    .B1(_03836_),
    .C1(_03837_),
    .Y(_03839_));
 sky130_fd_sc_hd__mux2_1 _10698_ (.A0(_02778_),
    .A1(_02782_),
    .S(net235),
    .X(_03840_));
 sky130_fd_sc_hd__inv_2 _10699_ (.A(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__mux2_1 _10700_ (.A0(_02963_),
    .A1(_03841_),
    .S(net237),
    .X(_03842_));
 sky130_fd_sc_hd__o21a_1 _10701_ (.A1(_03838_),
    .A2(_03839_),
    .B1(net263),
    .X(_03843_));
 sky130_fd_sc_hd__a211o_1 _10702_ (.A1(net241),
    .A2(_03842_),
    .B1(_03843_),
    .C1(net214),
    .X(_03844_));
 sky130_fd_sc_hd__or2_1 _10703_ (.A(\div_res[10] ),
    .B(_03726_),
    .X(_03845_));
 sky130_fd_sc_hd__a21oi_1 _10704_ (.A1(net23),
    .A2(_03845_),
    .B1(\div_res[11] ),
    .Y(_03846_));
 sky130_fd_sc_hd__a31o_1 _10705_ (.A1(\div_res[11] ),
    .A2(net23),
    .A3(_03845_),
    .B1(net202),
    .X(_03847_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(_02300_),
    .A1(_02294_),
    .S(_06198_),
    .X(_03848_));
 sky130_fd_sc_hd__o21a_1 _10707_ (.A1(net205),
    .A2(_03848_),
    .B1(_06207_),
    .X(_03849_));
 sky130_fd_sc_hd__or2_1 _10708_ (.A(\div_shifter[42] ),
    .B(_03731_),
    .X(_03850_));
 sky130_fd_sc_hd__a21oi_1 _10709_ (.A1(net246),
    .A2(_03850_),
    .B1(\div_shifter[43] ),
    .Y(_03851_));
 sky130_fd_sc_hd__a311o_2 _10710_ (.A1(\div_shifter[43] ),
    .A2(net247),
    .A3(_03850_),
    .B1(_03851_),
    .C1(net249),
    .X(_03852_));
 sky130_fd_sc_hd__a21oi_2 _10711_ (.A1(_06181_),
    .A2(net213),
    .B1(_03849_),
    .Y(_03853_));
 sky130_fd_sc_hd__o211a_1 _10712_ (.A1(_03846_),
    .A2(_03847_),
    .B1(_03852_),
    .C1(_03853_),
    .X(_03854_));
 sky130_fd_sc_hd__o21ai_2 _10713_ (.A1(net239),
    .A2(_02942_),
    .B1(_02312_),
    .Y(_03855_));
 sky130_fd_sc_hd__o221a_1 _10714_ (.A1(net182),
    .A2(_03842_),
    .B1(_03855_),
    .B2(net184),
    .C1(_03854_),
    .X(_03856_));
 sky130_fd_sc_hd__and3_1 _10715_ (.A(_03835_),
    .B(_03844_),
    .C(_03856_),
    .X(_03857_));
 sky130_fd_sc_hd__o211a_1 _10716_ (.A1(_03826_),
    .A2(_03827_),
    .B1(_03830_),
    .C1(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__nor2_1 _10717_ (.A(curr_PC[11]),
    .B(_03740_),
    .Y(_03859_));
 sky130_fd_sc_hd__and2_1 _10718_ (.A(curr_PC[11]),
    .B(_03740_),
    .X(_03860_));
 sky130_fd_sc_hd__or3_1 _10719_ (.A(net257),
    .B(_03859_),
    .C(_03860_),
    .X(_03861_));
 sky130_fd_sc_hd__o21ai_4 _10720_ (.A1(net262),
    .A2(_03858_),
    .B1(_03861_),
    .Y(dest_val[11]));
 sky130_fd_sc_hd__o21ai_2 _10721_ (.A1(_03809_),
    .A2(_03810_),
    .B1(_03812_),
    .Y(_03862_));
 sky130_fd_sc_hd__o22a_1 _10722_ (.A1(net81),
    .A2(net11),
    .B1(net44),
    .B2(net129),
    .X(_03863_));
 sky130_fd_sc_hd__xnor2_1 _10723_ (.A(net96),
    .B(_03863_),
    .Y(_03864_));
 sky130_fd_sc_hd__o22a_1 _10724_ (.A1(net122),
    .A2(net7),
    .B1(net5),
    .B2(net125),
    .X(_03865_));
 sky130_fd_sc_hd__xnor2_1 _10725_ (.A(net28),
    .B(_03865_),
    .Y(_03866_));
 sky130_fd_sc_hd__or2_1 _10726_ (.A(_03864_),
    .B(_03866_),
    .X(_03867_));
 sky130_fd_sc_hd__xor2_1 _10727_ (.A(_03864_),
    .B(_03866_),
    .X(_03868_));
 sky130_fd_sc_hd__a32o_1 _10728_ (.A1(_00219_),
    .A2(_00221_),
    .A3(_00392_),
    .B1(_00390_),
    .B2(_00197_),
    .X(_03869_));
 sky130_fd_sc_hd__xor2_2 _10729_ (.A(net137),
    .B(_03869_),
    .X(_03870_));
 sky130_fd_sc_hd__o22a_1 _10730_ (.A1(net64),
    .A2(net41),
    .B1(net39),
    .B2(net57),
    .X(_03871_));
 sky130_fd_sc_hd__xnor2_1 _10731_ (.A(net104),
    .B(_03871_),
    .Y(_03872_));
 sky130_fd_sc_hd__nand2_1 _10732_ (.A(_03870_),
    .B(_03872_),
    .Y(_03873_));
 sky130_fd_sc_hd__xor2_1 _10733_ (.A(_03870_),
    .B(_03872_),
    .X(_03874_));
 sky130_fd_sc_hd__o22a_1 _10734_ (.A1(net54),
    .A2(net37),
    .B1(net35),
    .B2(net62),
    .X(_03875_));
 sky130_fd_sc_hd__xnor2_1 _10735_ (.A(net136),
    .B(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__nand2_1 _10736_ (.A(_03874_),
    .B(_03876_),
    .Y(_03877_));
 sky130_fd_sc_hd__xor2_1 _10737_ (.A(_03874_),
    .B(_03876_),
    .X(_03878_));
 sky130_fd_sc_hd__xnor2_1 _10738_ (.A(_03868_),
    .B(_03878_),
    .Y(_03879_));
 sky130_fd_sc_hd__o22a_1 _10739_ (.A1(net118),
    .A2(net52),
    .B1(net99),
    .B2(net14),
    .X(_03880_));
 sky130_fd_sc_hd__xnor2_2 _10740_ (.A(net111),
    .B(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__o22a_1 _10741_ (.A1(net73),
    .A2(net50),
    .B1(net48),
    .B2(net67),
    .X(_03882_));
 sky130_fd_sc_hd__xnor2_1 _10742_ (.A(net105),
    .B(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__and2_1 _10743_ (.A(_03881_),
    .B(_03883_),
    .X(_03884_));
 sky130_fd_sc_hd__xor2_2 _10744_ (.A(_03881_),
    .B(_03883_),
    .X(_03885_));
 sky130_fd_sc_hd__o22a_1 _10745_ (.A1(net70),
    .A2(net13),
    .B1(net47),
    .B2(net76),
    .X(_03886_));
 sky130_fd_sc_hd__xnor2_2 _10746_ (.A(net108),
    .B(_03886_),
    .Y(_03887_));
 sky130_fd_sc_hd__xor2_1 _10747_ (.A(_03885_),
    .B(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__and2b_1 _10748_ (.A_N(_03879_),
    .B(_03888_),
    .X(_03889_));
 sky130_fd_sc_hd__xnor2_1 _10749_ (.A(_03879_),
    .B(_03888_),
    .Y(_03890_));
 sky130_fd_sc_hd__o211a_1 _10750_ (.A1(_03780_),
    .A2(_03784_),
    .B1(_00430_),
    .C1(net33),
    .X(_03891_));
 sky130_fd_sc_hd__a211oi_2 _10751_ (.A1(_00430_),
    .A2(net33),
    .B1(_03780_),
    .C1(_03784_),
    .Y(_03892_));
 sky130_fd_sc_hd__a211oi_2 _10752_ (.A1(_03748_),
    .A2(_03752_),
    .B1(_03891_),
    .C1(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__o211a_1 _10753_ (.A1(_03891_),
    .A2(_03892_),
    .B1(_03748_),
    .C1(_03752_),
    .X(_03894_));
 sky130_fd_sc_hd__nor2_1 _10754_ (.A(_03893_),
    .B(_03894_),
    .Y(_03895_));
 sky130_fd_sc_hd__nand2_1 _10755_ (.A(_03890_),
    .B(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__or2_1 _10756_ (.A(_03890_),
    .B(_03895_),
    .X(_03897_));
 sky130_fd_sc_hd__nand2_1 _10757_ (.A(_03896_),
    .B(_03897_),
    .Y(_03898_));
 sky130_fd_sc_hd__o21ai_1 _10758_ (.A1(_03788_),
    .A2(_03793_),
    .B1(_03792_),
    .Y(_03899_));
 sky130_fd_sc_hd__o22a_1 _10759_ (.A1(net78),
    .A2(net16),
    .B1(net9),
    .B2(net123),
    .X(_03900_));
 sky130_fd_sc_hd__xnor2_1 _10760_ (.A(net154),
    .B(_03900_),
    .Y(_03901_));
 sky130_fd_sc_hd__nand2_1 _10761_ (.A(_06443_),
    .B(_00756_),
    .Y(_03902_));
 sky130_fd_sc_hd__a22o_1 _10762_ (.A1(_06442_),
    .A2(_00756_),
    .B1(_03902_),
    .B2(_06435_),
    .X(_03903_));
 sky130_fd_sc_hd__nor2_1 _10763_ (.A(_03901_),
    .B(_03903_),
    .Y(_03904_));
 sky130_fd_sc_hd__and2_1 _10764_ (.A(_03901_),
    .B(_03903_),
    .X(_03905_));
 sky130_fd_sc_hd__or2_1 _10765_ (.A(_03904_),
    .B(_03905_),
    .X(_03906_));
 sky130_fd_sc_hd__o21a_1 _10766_ (.A1(_03769_),
    .A2(_03773_),
    .B1(_03906_),
    .X(_03907_));
 sky130_fd_sc_hd__nor3_1 _10767_ (.A(_03769_),
    .B(_03773_),
    .C(_03906_),
    .Y(_03908_));
 sky130_fd_sc_hd__nor2_1 _10768_ (.A(_03907_),
    .B(_03908_),
    .Y(_03909_));
 sky130_fd_sc_hd__and2_1 _10769_ (.A(_03899_),
    .B(_03909_),
    .X(_03910_));
 sky130_fd_sc_hd__xnor2_1 _10770_ (.A(_03899_),
    .B(_03909_),
    .Y(_03911_));
 sky130_fd_sc_hd__xor2_1 _10771_ (.A(_03898_),
    .B(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__o21ba_1 _10772_ (.A1(_03764_),
    .A2(_03799_),
    .B1_N(_03801_),
    .X(_03913_));
 sky130_fd_sc_hd__a21o_1 _10773_ (.A1(_03745_),
    .A2(_03758_),
    .B1(_03756_),
    .X(_03914_));
 sky130_fd_sc_hd__a21o_1 _10774_ (.A1(_03760_),
    .A2(_03763_),
    .B1(_03762_),
    .X(_03915_));
 sky130_fd_sc_hd__o21ai_1 _10775_ (.A1(_03795_),
    .A2(_03797_),
    .B1(_03915_),
    .Y(_03916_));
 sky130_fd_sc_hd__or3_1 _10776_ (.A(_03795_),
    .B(_03797_),
    .C(_03915_),
    .X(_03917_));
 sky130_fd_sc_hd__and2_1 _10777_ (.A(_03916_),
    .B(_03917_),
    .X(_03918_));
 sky130_fd_sc_hd__xnor2_1 _10778_ (.A(_03914_),
    .B(_03918_),
    .Y(_03919_));
 sky130_fd_sc_hd__a21bo_1 _10779_ (.A1(_03804_),
    .A2(_03808_),
    .B1_N(_03807_),
    .X(_03920_));
 sky130_fd_sc_hd__and2b_1 _10780_ (.A_N(_03919_),
    .B(_03920_),
    .X(_03921_));
 sky130_fd_sc_hd__xnor2_1 _10781_ (.A(_03919_),
    .B(_03920_),
    .Y(_03922_));
 sky130_fd_sc_hd__and2b_1 _10782_ (.A_N(_03913_),
    .B(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__xnor2_1 _10783_ (.A(_03913_),
    .B(_03922_),
    .Y(_03924_));
 sky130_fd_sc_hd__and2_1 _10784_ (.A(_03912_),
    .B(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__xnor2_1 _10785_ (.A(_03912_),
    .B(_03924_),
    .Y(_03926_));
 sky130_fd_sc_hd__and2b_1 _10786_ (.A_N(_03926_),
    .B(_03862_),
    .X(_03927_));
 sky130_fd_sc_hd__xor2_1 _10787_ (.A(_03862_),
    .B(_03926_),
    .X(_03928_));
 sky130_fd_sc_hd__a21oi_2 _10788_ (.A1(_03744_),
    .A2(_03815_),
    .B1(_03814_),
    .Y(_03929_));
 sky130_fd_sc_hd__nor2_1 _10789_ (.A(_03928_),
    .B(_03929_),
    .Y(_03930_));
 sky130_fd_sc_hd__and2_1 _10790_ (.A(_03928_),
    .B(_03929_),
    .X(_03931_));
 sky130_fd_sc_hd__nor2_1 _10791_ (.A(_03930_),
    .B(_03931_),
    .Y(_03932_));
 sky130_fd_sc_hd__and3_1 _10792_ (.A(_03701_),
    .B(_03702_),
    .C(_03820_),
    .X(_03933_));
 sky130_fd_sc_hd__and2b_1 _10793_ (.A_N(_03817_),
    .B(_03699_),
    .X(_03934_));
 sky130_fd_sc_hd__and3_1 _10794_ (.A(_03701_),
    .B(_03703_),
    .C(_03820_),
    .X(_03935_));
 sky130_fd_sc_hd__a2111o_4 _10795_ (.A1(_03462_),
    .A2(_03935_),
    .B1(_03934_),
    .C1(_03933_),
    .D1(_03818_),
    .X(_03936_));
 sky130_fd_sc_hd__xnor2_2 _10796_ (.A(_03932_),
    .B(_03936_),
    .Y(_03937_));
 sky130_fd_sc_hd__a21o_1 _10797_ (.A1(_03822_),
    .A2(_03824_),
    .B1(net84),
    .X(_03938_));
 sky130_fd_sc_hd__o21ai_1 _10798_ (.A1(_03937_),
    .A2(_03938_),
    .B1(net206),
    .Y(_03939_));
 sky130_fd_sc_hd__a21o_1 _10799_ (.A1(_03937_),
    .A2(_03938_),
    .B1(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__nor3_1 _10800_ (.A(net84),
    .B(_02156_),
    .C(_02179_),
    .Y(_03941_));
 sky130_fd_sc_hd__o21a_1 _10801_ (.A1(net84),
    .A2(_02179_),
    .B1(_02156_),
    .X(_03942_));
 sky130_fd_sc_hd__o21a_1 _10802_ (.A1(_06216_),
    .A2(_03832_),
    .B1(_06198_),
    .X(_03943_));
 sky130_fd_sc_hd__and2_1 _10803_ (.A(_04504_),
    .B(_03943_),
    .X(_03944_));
 sky130_fd_sc_hd__a21oi_1 _10804_ (.A1(_06189_),
    .A2(_06323_),
    .B1(_04504_),
    .Y(_03945_));
 sky130_fd_sc_hd__o21ai_1 _10805_ (.A1(_03944_),
    .A2(_03945_),
    .B1(_06163_),
    .Y(_03946_));
 sky130_fd_sc_hd__o31a_1 _10806_ (.A1(_06163_),
    .A2(_03944_),
    .A3(_03945_),
    .B1(net251),
    .X(_03947_));
 sky130_fd_sc_hd__nand2_1 _10807_ (.A(_03946_),
    .B(_03947_),
    .Y(_03948_));
 sky130_fd_sc_hd__mux2_1 _10808_ (.A0(_02939_),
    .A1(_02941_),
    .S(net234),
    .X(_03949_));
 sky130_fd_sc_hd__or2_1 _10809_ (.A(net238),
    .B(_03949_),
    .X(_03950_));
 sky130_fd_sc_hd__o21ai_4 _10810_ (.A1(net237),
    .A2(_02806_),
    .B1(_03950_),
    .Y(_03951_));
 sky130_fd_sc_hd__or2_1 _10811_ (.A(reg1_val[12]),
    .B(curr_PC[12]),
    .X(_03952_));
 sky130_fd_sc_hd__nand2_1 _10812_ (.A(reg1_val[12]),
    .B(curr_PC[12]),
    .Y(_03953_));
 sky130_fd_sc_hd__o211a_1 _10813_ (.A1(_03837_),
    .A2(_03839_),
    .B1(_03952_),
    .C1(_03953_),
    .X(_03954_));
 sky130_fd_sc_hd__a211o_1 _10814_ (.A1(_03952_),
    .A2(_03953_),
    .B1(_03837_),
    .C1(_03839_),
    .X(_03955_));
 sky130_fd_sc_hd__nand2_1 _10815_ (.A(net263),
    .B(_03955_),
    .Y(_03956_));
 sky130_fd_sc_hd__o22a_1 _10816_ (.A1(net263),
    .A2(_03951_),
    .B1(_03954_),
    .B2(_03956_),
    .X(_03957_));
 sky130_fd_sc_hd__or2_1 _10817_ (.A(\div_res[11] ),
    .B(_03845_),
    .X(_03958_));
 sky130_fd_sc_hd__a21oi_1 _10818_ (.A1(net23),
    .A2(_03958_),
    .B1(\div_res[12] ),
    .Y(_03959_));
 sky130_fd_sc_hd__a311o_1 _10819_ (.A1(\div_res[12] ),
    .A2(net23),
    .A3(_03958_),
    .B1(_03959_),
    .C1(net202),
    .X(_03960_));
 sky130_fd_sc_hd__or2_1 _10820_ (.A(\div_shifter[43] ),
    .B(_03850_),
    .X(_03961_));
 sky130_fd_sc_hd__a21oi_1 _10821_ (.A1(net247),
    .A2(_03961_),
    .B1(\div_shifter[44] ),
    .Y(_03962_));
 sky130_fd_sc_hd__a311o_1 _10822_ (.A1(\div_shifter[44] ),
    .A2(net246),
    .A3(_03961_),
    .B1(_03962_),
    .C1(net249),
    .X(_03963_));
 sky130_fd_sc_hd__nor2_1 _10823_ (.A(_06145_),
    .B(net204),
    .Y(_03964_));
 sky130_fd_sc_hd__a211o_1 _10824_ (.A1(_06145_),
    .A2(_02294_),
    .B1(_03964_),
    .C1(net205),
    .X(_03965_));
 sky130_fd_sc_hd__a22oi_2 _10825_ (.A1(_06127_),
    .A2(net212),
    .B1(_03965_),
    .B2(_06154_),
    .Y(_03966_));
 sky130_fd_sc_hd__and3_1 _10826_ (.A(_03960_),
    .B(_03963_),
    .C(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__o21a_1 _10827_ (.A1(net238),
    .A2(_02786_),
    .B1(_02312_),
    .X(_03968_));
 sky130_fd_sc_hd__inv_2 _10828_ (.A(_03968_),
    .Y(_03969_));
 sky130_fd_sc_hd__o221a_1 _10829_ (.A1(net182),
    .A2(_03951_),
    .B1(_03969_),
    .B2(net186),
    .C1(_03967_),
    .X(_03970_));
 sky130_fd_sc_hd__o211a_1 _10830_ (.A1(net214),
    .A2(_03957_),
    .B1(_03970_),
    .C1(_03948_),
    .X(_03971_));
 sky130_fd_sc_hd__o311a_1 _10831_ (.A1(net250),
    .A2(_03941_),
    .A3(_03942_),
    .B1(_03971_),
    .C1(_03940_),
    .X(_03972_));
 sky130_fd_sc_hd__and3_2 _10832_ (.A(curr_PC[11]),
    .B(curr_PC[12]),
    .C(_03740_),
    .X(_03973_));
 sky130_fd_sc_hd__o21ai_1 _10833_ (.A1(curr_PC[12]),
    .A2(_03860_),
    .B1(net262),
    .Y(_03974_));
 sky130_fd_sc_hd__o22ai_4 _10834_ (.A1(net262),
    .A2(_03972_),
    .B1(_03973_),
    .B2(_03974_),
    .Y(dest_val[12]));
 sky130_fd_sc_hd__o22a_1 _10835_ (.A1(net129),
    .A2(net11),
    .B1(net44),
    .B2(net99),
    .X(_03975_));
 sky130_fd_sc_hd__xnor2_1 _10836_ (.A(net96),
    .B(_03975_),
    .Y(_03976_));
 sky130_fd_sc_hd__o22a_1 _10837_ (.A1(net76),
    .A2(net13),
    .B1(net47),
    .B2(net73),
    .X(_03977_));
 sky130_fd_sc_hd__xnor2_1 _10838_ (.A(net108),
    .B(_03977_),
    .Y(_03978_));
 sky130_fd_sc_hd__nand2b_1 _10839_ (.A_N(_03976_),
    .B(_03978_),
    .Y(_03979_));
 sky130_fd_sc_hd__xor2_1 _10840_ (.A(_03976_),
    .B(_03978_),
    .X(_03980_));
 sky130_fd_sc_hd__o22a_1 _10841_ (.A1(net118),
    .A2(net14),
    .B1(net52),
    .B2(net70),
    .X(_03981_));
 sky130_fd_sc_hd__xnor2_1 _10842_ (.A(net111),
    .B(_03981_),
    .Y(_03982_));
 sky130_fd_sc_hd__nand2b_1 _10843_ (.A_N(_03980_),
    .B(_03982_),
    .Y(_03983_));
 sky130_fd_sc_hd__xnor2_1 _10844_ (.A(_03980_),
    .B(_03982_),
    .Y(_03984_));
 sky130_fd_sc_hd__and3_1 _10845_ (.A(_00219_),
    .B(_00221_),
    .C(_00390_),
    .X(_03985_));
 sky130_fd_sc_hd__a21oi_1 _10846_ (.A1(_00225_),
    .A2(_00226_),
    .B1(net94),
    .Y(_03986_));
 sky130_fd_sc_hd__or3b_1 _10847_ (.A(_03985_),
    .B(_03986_),
    .C_N(net137),
    .X(_03987_));
 sky130_fd_sc_hd__o21bai_1 _10848_ (.A1(_03985_),
    .A2(_03986_),
    .B1_N(net137),
    .Y(_03988_));
 sky130_fd_sc_hd__a21o_1 _10849_ (.A1(_03987_),
    .A2(_03988_),
    .B1(_06435_),
    .X(_03989_));
 sky130_fd_sc_hd__nand3_1 _10850_ (.A(_06435_),
    .B(_03987_),
    .C(_03988_),
    .Y(_03990_));
 sky130_fd_sc_hd__and2_1 _10851_ (.A(_03989_),
    .B(_03990_),
    .X(_03991_));
 sky130_fd_sc_hd__o22a_1 _10852_ (.A1(net78),
    .A2(net9),
    .B1(net3),
    .B2(net123),
    .X(_03992_));
 sky130_fd_sc_hd__xnor2_1 _10853_ (.A(net156),
    .B(_03992_),
    .Y(_03993_));
 sky130_fd_sc_hd__nand2_1 _10854_ (.A(_03991_),
    .B(_03993_),
    .Y(_03994_));
 sky130_fd_sc_hd__or2_1 _10855_ (.A(_03991_),
    .B(_03993_),
    .X(_03995_));
 sky130_fd_sc_hd__and3_1 _10856_ (.A(_03984_),
    .B(_03994_),
    .C(_03995_),
    .X(_03996_));
 sky130_fd_sc_hd__a21oi_1 _10857_ (.A1(_03994_),
    .A2(_03995_),
    .B1(_03984_),
    .Y(_03997_));
 sky130_fd_sc_hd__o22a_1 _10858_ (.A1(net67),
    .A2(net50),
    .B1(net48),
    .B2(net64),
    .X(_03998_));
 sky130_fd_sc_hd__xnor2_1 _10859_ (.A(net105),
    .B(_03998_),
    .Y(_03999_));
 sky130_fd_sc_hd__o22a_1 _10860_ (.A1(net62),
    .A2(net37),
    .B1(net35),
    .B2(net60),
    .X(_04000_));
 sky130_fd_sc_hd__xnor2_1 _10861_ (.A(net136),
    .B(_04000_),
    .Y(_04001_));
 sky130_fd_sc_hd__and2_1 _10862_ (.A(_03999_),
    .B(_04001_),
    .X(_04002_));
 sky130_fd_sc_hd__nor2_1 _10863_ (.A(_03999_),
    .B(_04001_),
    .Y(_04003_));
 sky130_fd_sc_hd__nor2_1 _10864_ (.A(_04002_),
    .B(_04003_),
    .Y(_04004_));
 sky130_fd_sc_hd__o22a_1 _10865_ (.A1(net57),
    .A2(net41),
    .B1(net39),
    .B2(net54),
    .X(_04005_));
 sky130_fd_sc_hd__xnor2_1 _10866_ (.A(net104),
    .B(_04005_),
    .Y(_04006_));
 sky130_fd_sc_hd__xnor2_1 _10867_ (.A(_04004_),
    .B(_04006_),
    .Y(_04007_));
 sky130_fd_sc_hd__or3_1 _10868_ (.A(_03996_),
    .B(_03997_),
    .C(_04007_),
    .X(_04008_));
 sky130_fd_sc_hd__o21ai_1 _10869_ (.A1(_03996_),
    .A2(_03997_),
    .B1(_04007_),
    .Y(_04009_));
 sky130_fd_sc_hd__o22a_1 _10870_ (.A1(net81),
    .A2(net7),
    .B1(net5),
    .B2(net122),
    .X(_04010_));
 sky130_fd_sc_hd__xnor2_1 _10871_ (.A(net28),
    .B(_04010_),
    .Y(_04011_));
 sky130_fd_sc_hd__nor2_1 _10872_ (.A(_03904_),
    .B(_04011_),
    .Y(_04012_));
 sky130_fd_sc_hd__and2_1 _10873_ (.A(_03904_),
    .B(_04011_),
    .X(_04013_));
 sky130_fd_sc_hd__nor2_1 _10874_ (.A(_04012_),
    .B(_04013_),
    .Y(_04014_));
 sky130_fd_sc_hd__and3b_1 _10875_ (.A_N(net125),
    .B(net33),
    .C(_04014_),
    .X(_04015_));
 sky130_fd_sc_hd__o21ba_1 _10876_ (.A1(net125),
    .A2(net28),
    .B1_N(_04014_),
    .X(_04016_));
 sky130_fd_sc_hd__nor2_1 _10877_ (.A(_04015_),
    .B(_04016_),
    .Y(_04017_));
 sky130_fd_sc_hd__and3_1 _10878_ (.A(_04008_),
    .B(_04009_),
    .C(_04017_),
    .X(_04018_));
 sky130_fd_sc_hd__a21oi_1 _10879_ (.A1(_04008_),
    .A2(_04009_),
    .B1(_04017_),
    .Y(_04019_));
 sky130_fd_sc_hd__nor2_1 _10880_ (.A(_04018_),
    .B(_04019_),
    .Y(_04020_));
 sky130_fd_sc_hd__a21oi_2 _10881_ (.A1(_03885_),
    .A2(_03887_),
    .B1(_03884_),
    .Y(_04021_));
 sky130_fd_sc_hd__a21oi_1 _10882_ (.A1(_03873_),
    .A2(_03877_),
    .B1(_03867_),
    .Y(_04022_));
 sky130_fd_sc_hd__and3_1 _10883_ (.A(_03867_),
    .B(_03873_),
    .C(_03877_),
    .X(_04023_));
 sky130_fd_sc_hd__or2_1 _10884_ (.A(_04022_),
    .B(_04023_),
    .X(_04024_));
 sky130_fd_sc_hd__xnor2_1 _10885_ (.A(_04021_),
    .B(_04024_),
    .Y(_04025_));
 sky130_fd_sc_hd__xnor2_1 _10886_ (.A(_04020_),
    .B(_04025_),
    .Y(_04026_));
 sky130_fd_sc_hd__o21ai_1 _10887_ (.A1(_03898_),
    .A2(_03911_),
    .B1(_03896_),
    .Y(_04027_));
 sky130_fd_sc_hd__a21bo_1 _10888_ (.A1(_03914_),
    .A2(_03918_),
    .B1_N(_03916_),
    .X(_04028_));
 sky130_fd_sc_hd__a21o_1 _10889_ (.A1(_03868_),
    .A2(_03878_),
    .B1(_03889_),
    .X(_04029_));
 sky130_fd_sc_hd__nor2_1 _10890_ (.A(_03891_),
    .B(_03893_),
    .Y(_04030_));
 sky130_fd_sc_hd__o21ai_1 _10891_ (.A1(_03891_),
    .A2(_03893_),
    .B1(_04029_),
    .Y(_04031_));
 sky130_fd_sc_hd__xnor2_1 _10892_ (.A(_04029_),
    .B(_04030_),
    .Y(_04032_));
 sky130_fd_sc_hd__o21ai_1 _10893_ (.A1(_03907_),
    .A2(_03910_),
    .B1(_04032_),
    .Y(_04033_));
 sky130_fd_sc_hd__or3_1 _10894_ (.A(_03907_),
    .B(_03910_),
    .C(_04032_),
    .X(_04034_));
 sky130_fd_sc_hd__and2_1 _10895_ (.A(_04033_),
    .B(_04034_),
    .X(_04035_));
 sky130_fd_sc_hd__xnor2_1 _10896_ (.A(_04028_),
    .B(_04035_),
    .Y(_04036_));
 sky130_fd_sc_hd__nand2b_1 _10897_ (.A_N(_04036_),
    .B(_04027_),
    .Y(_04037_));
 sky130_fd_sc_hd__xnor2_1 _10898_ (.A(_04027_),
    .B(_04036_),
    .Y(_04038_));
 sky130_fd_sc_hd__xor2_1 _10899_ (.A(_04026_),
    .B(_04038_),
    .X(_04039_));
 sky130_fd_sc_hd__nor2_1 _10900_ (.A(_03921_),
    .B(_03923_),
    .Y(_04040_));
 sky130_fd_sc_hd__nand2b_1 _10901_ (.A_N(_04040_),
    .B(_04039_),
    .Y(_04041_));
 sky130_fd_sc_hd__xnor2_1 _10902_ (.A(_04039_),
    .B(_04040_),
    .Y(_04042_));
 sky130_fd_sc_hd__o21a_1 _10903_ (.A1(_03925_),
    .A2(_03927_),
    .B1(_04042_),
    .X(_04043_));
 sky130_fd_sc_hd__nor3_1 _10904_ (.A(_03925_),
    .B(_03927_),
    .C(_04042_),
    .Y(_04044_));
 sky130_fd_sc_hd__nor2_1 _10905_ (.A(_04043_),
    .B(_04044_),
    .Y(_04045_));
 sky130_fd_sc_hd__a21oi_1 _10906_ (.A1(_03932_),
    .A2(_03936_),
    .B1(_03930_),
    .Y(_04046_));
 sky130_fd_sc_hd__xor2_2 _10907_ (.A(_04045_),
    .B(_04046_),
    .X(_04047_));
 sky130_fd_sc_hd__and4b_1 _10908_ (.A_N(_03591_),
    .B(_03822_),
    .C(_03823_),
    .D(_03937_),
    .X(_04048_));
 sky130_fd_sc_hd__or2_1 _10909_ (.A(net84),
    .B(_04048_),
    .X(_04049_));
 sky130_fd_sc_hd__a21oi_1 _10910_ (.A1(_04047_),
    .A2(_04049_),
    .B1(_02214_),
    .Y(_04050_));
 sky130_fd_sc_hd__o21ai_1 _10911_ (.A1(_04047_),
    .A2(_04049_),
    .B1(_04050_),
    .Y(_04051_));
 sky130_fd_sc_hd__o21a_1 _10912_ (.A1(net84),
    .A2(_02180_),
    .B1(_02155_),
    .X(_04052_));
 sky130_fd_sc_hd__nor3_1 _10913_ (.A(net84),
    .B(_02155_),
    .C(_02180_),
    .Y(_04053_));
 sky130_fd_sc_hd__and3_1 _10914_ (.A(net305),
    .B(_06136_),
    .C(_06324_),
    .X(_04054_));
 sky130_fd_sc_hd__o21a_1 _10915_ (.A1(_06163_),
    .A2(_03943_),
    .B1(_06145_),
    .X(_04055_));
 sky130_fd_sc_hd__o21ba_1 _10916_ (.A1(net305),
    .A2(_04055_),
    .B1_N(_04054_),
    .X(_04056_));
 sky130_fd_sc_hd__nor2_1 _10917_ (.A(_06109_),
    .B(_04056_),
    .Y(_04057_));
 sky130_fd_sc_hd__a211o_1 _10918_ (.A1(_06109_),
    .A2(_04056_),
    .B1(_04057_),
    .C1(_02293_),
    .X(_04058_));
 sky130_fd_sc_hd__or2_1 _10919_ (.A(net303),
    .B(curr_PC[13]),
    .X(_04059_));
 sky130_fd_sc_hd__nand2_1 _10920_ (.A(net303),
    .B(curr_PC[13]),
    .Y(_04060_));
 sky130_fd_sc_hd__nand2_1 _10921_ (.A(_04059_),
    .B(_04060_),
    .Y(_04061_));
 sky130_fd_sc_hd__a21oi_1 _10922_ (.A1(reg1_val[12]),
    .A2(curr_PC[12]),
    .B1(_03954_),
    .Y(_04062_));
 sky130_fd_sc_hd__xnor2_1 _10923_ (.A(_04061_),
    .B(_04062_),
    .Y(_04063_));
 sky130_fd_sc_hd__mux2_1 _10924_ (.A0(_03082_),
    .A1(_03086_),
    .S(net236),
    .X(_04064_));
 sky130_fd_sc_hd__mux2_1 _10925_ (.A0(_02624_),
    .A1(_04064_),
    .S(net237),
    .X(_04065_));
 sky130_fd_sc_hd__mux2_1 _10926_ (.A0(_04063_),
    .A1(_04065_),
    .S(net241),
    .X(_04066_));
 sky130_fd_sc_hd__or2_1 _10927_ (.A(\div_res[12] ),
    .B(_03958_),
    .X(_04067_));
 sky130_fd_sc_hd__a21oi_1 _10928_ (.A1(net24),
    .A2(_04067_),
    .B1(\div_res[13] ),
    .Y(_04068_));
 sky130_fd_sc_hd__a311o_1 _10929_ (.A1(\div_res[13] ),
    .A2(net24),
    .A3(_04067_),
    .B1(_04068_),
    .C1(net203),
    .X(_04069_));
 sky130_fd_sc_hd__or2_1 _10930_ (.A(\div_shifter[44] ),
    .B(_03961_),
    .X(_04070_));
 sky130_fd_sc_hd__a21oi_1 _10931_ (.A1(net245),
    .A2(_04070_),
    .B1(\div_shifter[45] ),
    .Y(_04071_));
 sky130_fd_sc_hd__a31o_1 _10932_ (.A1(\div_shifter[45] ),
    .A2(net245),
    .A3(_04070_),
    .B1(net248),
    .X(_04072_));
 sky130_fd_sc_hd__nor2_1 _10933_ (.A(_06094_),
    .B(net204),
    .Y(_04073_));
 sky130_fd_sc_hd__a211o_1 _10934_ (.A1(_06094_),
    .A2(_02294_),
    .B1(_04073_),
    .C1(net205),
    .X(_04074_));
 sky130_fd_sc_hd__a22oi_2 _10935_ (.A1(_06082_),
    .A2(net212),
    .B1(_04074_),
    .B2(_06100_),
    .Y(_04075_));
 sky130_fd_sc_hd__o211a_1 _10936_ (.A1(_04071_),
    .A2(_04072_),
    .B1(_04075_),
    .C1(_04069_),
    .X(_04076_));
 sky130_fd_sc_hd__o21a_1 _10937_ (.A1(net238),
    .A2(_02638_),
    .B1(_02312_),
    .X(_04077_));
 sky130_fd_sc_hd__inv_2 _10938_ (.A(_04077_),
    .Y(_04078_));
 sky130_fd_sc_hd__o221a_1 _10939_ (.A1(net182),
    .A2(_04065_),
    .B1(_04078_),
    .B2(net184),
    .C1(_04076_),
    .X(_04079_));
 sky130_fd_sc_hd__o211a_1 _10940_ (.A1(net214),
    .A2(_04066_),
    .B1(_04079_),
    .C1(_04058_),
    .X(_04080_));
 sky130_fd_sc_hd__o311a_1 _10941_ (.A1(net250),
    .A2(_04052_),
    .A3(_04053_),
    .B1(_04080_),
    .C1(_04051_),
    .X(_04081_));
 sky130_fd_sc_hd__a21oi_1 _10942_ (.A1(curr_PC[13]),
    .A2(_03973_),
    .B1(net257),
    .Y(_04082_));
 sky130_fd_sc_hd__o21ai_2 _10943_ (.A1(curr_PC[13]),
    .A2(_03973_),
    .B1(_04082_),
    .Y(_04083_));
 sky130_fd_sc_hd__o21ai_4 _10944_ (.A1(net262),
    .A2(_04081_),
    .B1(_04083_),
    .Y(dest_val[13]));
 sky130_fd_sc_hd__a21bo_1 _10945_ (.A1(_04026_),
    .A2(_04038_),
    .B1_N(_04041_),
    .X(_04084_));
 sky130_fd_sc_hd__a21bo_1 _10946_ (.A1(_04028_),
    .A2(_04035_),
    .B1_N(_04037_),
    .X(_04085_));
 sky130_fd_sc_hd__a21o_1 _10947_ (.A1(_04004_),
    .A2(_04006_),
    .B1(_04002_),
    .X(_04086_));
 sky130_fd_sc_hd__and2_1 _10948_ (.A(_03989_),
    .B(_03994_),
    .X(_04087_));
 sky130_fd_sc_hd__a21oi_1 _10949_ (.A1(_03979_),
    .A2(_03983_),
    .B1(_04087_),
    .Y(_04088_));
 sky130_fd_sc_hd__and3_1 _10950_ (.A(_03979_),
    .B(_03983_),
    .C(_04087_),
    .X(_04089_));
 sky130_fd_sc_hd__nor2_1 _10951_ (.A(_04088_),
    .B(_04089_),
    .Y(_04090_));
 sky130_fd_sc_hd__xnor2_1 _10952_ (.A(_04086_),
    .B(_04090_),
    .Y(_04091_));
 sky130_fd_sc_hd__o22a_1 _10953_ (.A1(net129),
    .A2(net7),
    .B1(net5),
    .B2(net81),
    .X(_04092_));
 sky130_fd_sc_hd__xnor2_1 _10954_ (.A(net28),
    .B(_04092_),
    .Y(_04093_));
 sky130_fd_sc_hd__o22a_1 _10955_ (.A1(net99),
    .A2(net11),
    .B1(net44),
    .B2(net118),
    .X(_04094_));
 sky130_fd_sc_hd__xnor2_1 _10956_ (.A(net96),
    .B(_04094_),
    .Y(_04095_));
 sky130_fd_sc_hd__or3_1 _10957_ (.A(net122),
    .B(net28),
    .C(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__o21ai_1 _10958_ (.A1(net122),
    .A2(net28),
    .B1(_04095_),
    .Y(_04097_));
 sky130_fd_sc_hd__and2_1 _10959_ (.A(_04096_),
    .B(_04097_),
    .X(_04098_));
 sky130_fd_sc_hd__nand2b_1 _10960_ (.A_N(_04093_),
    .B(_04098_),
    .Y(_04099_));
 sky130_fd_sc_hd__xor2_1 _10961_ (.A(_04093_),
    .B(_04098_),
    .X(_04100_));
 sky130_fd_sc_hd__o22a_1 _10962_ (.A1(net60),
    .A2(net37),
    .B1(net35),
    .B2(net18),
    .X(_04101_));
 sky130_fd_sc_hd__xnor2_1 _10963_ (.A(net136),
    .B(_04101_),
    .Y(_04102_));
 sky130_fd_sc_hd__o22a_1 _10964_ (.A1(net64),
    .A2(net50),
    .B1(net48),
    .B2(net57),
    .X(_04103_));
 sky130_fd_sc_hd__xnor2_1 _10965_ (.A(net105),
    .B(_04103_),
    .Y(_04104_));
 sky130_fd_sc_hd__and2_1 _10966_ (.A(_04102_),
    .B(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__nor2_1 _10967_ (.A(_04102_),
    .B(_04104_),
    .Y(_04106_));
 sky130_fd_sc_hd__nor2_1 _10968_ (.A(_04105_),
    .B(_04106_),
    .Y(_04107_));
 sky130_fd_sc_hd__o22a_1 _10969_ (.A1(net54),
    .A2(net41),
    .B1(net39),
    .B2(net62),
    .X(_04108_));
 sky130_fd_sc_hd__xnor2_1 _10970_ (.A(net104),
    .B(_04108_),
    .Y(_04109_));
 sky130_fd_sc_hd__xor2_1 _10971_ (.A(_04107_),
    .B(_04109_),
    .X(_04110_));
 sky130_fd_sc_hd__o22a_1 _10972_ (.A1(net73),
    .A2(net13),
    .B1(net47),
    .B2(net67),
    .X(_04111_));
 sky130_fd_sc_hd__xnor2_1 _10973_ (.A(net108),
    .B(_04111_),
    .Y(_04112_));
 sky130_fd_sc_hd__o22a_1 _10974_ (.A1(net71),
    .A2(net14),
    .B1(net52),
    .B2(net76),
    .X(_04113_));
 sky130_fd_sc_hd__xnor2_1 _10975_ (.A(net111),
    .B(_04113_),
    .Y(_04114_));
 sky130_fd_sc_hd__and2_1 _10976_ (.A(_04112_),
    .B(_04114_),
    .X(_04115_));
 sky130_fd_sc_hd__nor2_1 _10977_ (.A(_04112_),
    .B(_04114_),
    .Y(_04116_));
 sky130_fd_sc_hd__nor2_1 _10978_ (.A(_04115_),
    .B(_04116_),
    .Y(_04117_));
 sky130_fd_sc_hd__o22a_1 _10979_ (.A1(net17),
    .A2(net42),
    .B1(net94),
    .B2(net10),
    .X(_04118_));
 sky130_fd_sc_hd__xnor2_1 _10980_ (.A(net137),
    .B(_04118_),
    .Y(_04119_));
 sky130_fd_sc_hd__o21a_1 _10981_ (.A1(_06476_),
    .A2(net4),
    .B1(net155),
    .X(_04120_));
 sky130_fd_sc_hd__nor2_1 _10982_ (.A(_06475_),
    .B(net4),
    .Y(_04121_));
 sky130_fd_sc_hd__nor3_2 _10983_ (.A(_04119_),
    .B(_04120_),
    .C(_04121_),
    .Y(_04122_));
 sky130_fd_sc_hd__o21a_1 _10984_ (.A1(_04120_),
    .A2(_04121_),
    .B1(_04119_),
    .X(_04123_));
 sky130_fd_sc_hd__nor2_1 _10985_ (.A(_04122_),
    .B(_04123_),
    .Y(_04124_));
 sky130_fd_sc_hd__xnor2_1 _10986_ (.A(_04117_),
    .B(_04124_),
    .Y(_04125_));
 sky130_fd_sc_hd__nand2_1 _10987_ (.A(_04110_),
    .B(_04125_),
    .Y(_04126_));
 sky130_fd_sc_hd__or2_1 _10988_ (.A(_04110_),
    .B(_04125_),
    .X(_04127_));
 sky130_fd_sc_hd__nand2_1 _10989_ (.A(_04126_),
    .B(_04127_),
    .Y(_04128_));
 sky130_fd_sc_hd__or2_1 _10990_ (.A(_04100_),
    .B(_04128_),
    .X(_04129_));
 sky130_fd_sc_hd__nand2_1 _10991_ (.A(_04100_),
    .B(_04128_),
    .Y(_04130_));
 sky130_fd_sc_hd__nand2_1 _10992_ (.A(_04129_),
    .B(_04130_),
    .Y(_04131_));
 sky130_fd_sc_hd__xor2_1 _10993_ (.A(_04091_),
    .B(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__o21ba_1 _10994_ (.A1(_04019_),
    .A2(_04025_),
    .B1_N(_04018_),
    .X(_04133_));
 sky130_fd_sc_hd__o21bai_2 _10995_ (.A1(_04021_),
    .A2(_04024_),
    .B1_N(_04022_),
    .Y(_04134_));
 sky130_fd_sc_hd__nand2b_1 _10996_ (.A_N(_03996_),
    .B(_04008_),
    .Y(_04135_));
 sky130_fd_sc_hd__nor2_1 _10997_ (.A(_04012_),
    .B(_04015_),
    .Y(_04136_));
 sky130_fd_sc_hd__o21ai_1 _10998_ (.A1(_04012_),
    .A2(_04015_),
    .B1(_04135_),
    .Y(_04137_));
 sky130_fd_sc_hd__xnor2_1 _10999_ (.A(_04135_),
    .B(_04136_),
    .Y(_04138_));
 sky130_fd_sc_hd__xnor2_1 _11000_ (.A(_04134_),
    .B(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__nand2_1 _11001_ (.A(_04031_),
    .B(_04033_),
    .Y(_04140_));
 sky130_fd_sc_hd__nand2b_1 _11002_ (.A_N(_04139_),
    .B(_04140_),
    .Y(_04141_));
 sky130_fd_sc_hd__and3_1 _11003_ (.A(_04031_),
    .B(_04033_),
    .C(_04139_),
    .X(_04142_));
 sky130_fd_sc_hd__xnor2_1 _11004_ (.A(_04139_),
    .B(_04140_),
    .Y(_04143_));
 sky130_fd_sc_hd__xnor2_1 _11005_ (.A(_04133_),
    .B(_04143_),
    .Y(_04144_));
 sky130_fd_sc_hd__nand2_1 _11006_ (.A(_04132_),
    .B(_04144_),
    .Y(_04145_));
 sky130_fd_sc_hd__or2_1 _11007_ (.A(_04132_),
    .B(_04144_),
    .X(_04146_));
 sky130_fd_sc_hd__nand2_1 _11008_ (.A(_04145_),
    .B(_04146_),
    .Y(_04147_));
 sky130_fd_sc_hd__nand2b_1 _11009_ (.A_N(_04147_),
    .B(_04085_),
    .Y(_04148_));
 sky130_fd_sc_hd__xnor2_2 _11010_ (.A(_04085_),
    .B(_04147_),
    .Y(_04149_));
 sky130_fd_sc_hd__and2_1 _11011_ (.A(_04084_),
    .B(_04149_),
    .X(_04150_));
 sky130_fd_sc_hd__xor2_2 _11012_ (.A(_04084_),
    .B(_04149_),
    .X(_04151_));
 sky130_fd_sc_hd__o21ba_1 _11013_ (.A1(_03930_),
    .A2(_04043_),
    .B1_N(_04044_),
    .X(_04152_));
 sky130_fd_sc_hd__and2_1 _11014_ (.A(_03932_),
    .B(_04045_),
    .X(_04153_));
 sky130_fd_sc_hd__a21o_1 _11015_ (.A1(_03936_),
    .A2(_04153_),
    .B1(_04152_),
    .X(_04154_));
 sky130_fd_sc_hd__xnor2_2 _11016_ (.A(_04151_),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__a21o_1 _11017_ (.A1(_04047_),
    .A2(_04048_),
    .B1(net84),
    .X(_04156_));
 sky130_fd_sc_hd__o21ai_1 _11018_ (.A1(_04155_),
    .A2(_04156_),
    .B1(net206),
    .Y(_04157_));
 sky130_fd_sc_hd__a21o_1 _11019_ (.A1(_04155_),
    .A2(_04156_),
    .B1(_04157_),
    .X(_04158_));
 sky130_fd_sc_hd__a21oi_1 _11020_ (.A1(net19),
    .A2(_02181_),
    .B1(_02183_),
    .Y(_04159_));
 sky130_fd_sc_hd__a31o_1 _11021_ (.A1(net19),
    .A2(_02181_),
    .A3(_02183_),
    .B1(net250),
    .X(_04160_));
 sky130_fd_sc_hd__or2_1 _11022_ (.A(_04159_),
    .B(_04160_),
    .X(_04161_));
 sky130_fd_sc_hd__and3_1 _11023_ (.A(net305),
    .B(_06088_),
    .C(_06325_),
    .X(_04162_));
 sky130_fd_sc_hd__o21a_1 _11024_ (.A1(_06109_),
    .A2(_04055_),
    .B1(_06094_),
    .X(_04163_));
 sky130_fd_sc_hd__o21ba_1 _11025_ (.A1(net305),
    .A2(_04163_),
    .B1_N(_04162_),
    .X(_04164_));
 sky130_fd_sc_hd__nor2_1 _11026_ (.A(_06070_),
    .B(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__a211o_1 _11027_ (.A1(_06070_),
    .A2(_04164_),
    .B1(_04165_),
    .C1(_02293_),
    .X(_04166_));
 sky130_fd_sc_hd__or2_1 _11028_ (.A(reg1_val[14]),
    .B(curr_PC[14]),
    .X(_04167_));
 sky130_fd_sc_hd__nand2_1 _11029_ (.A(reg1_val[14]),
    .B(curr_PC[14]),
    .Y(_04168_));
 sky130_fd_sc_hd__nand2_1 _11030_ (.A(_04167_),
    .B(_04168_),
    .Y(_04169_));
 sky130_fd_sc_hd__o21a_1 _11031_ (.A1(_04061_),
    .A2(_04062_),
    .B1(_04060_),
    .X(_04170_));
 sky130_fd_sc_hd__xnor2_1 _11032_ (.A(_04169_),
    .B(_04170_),
    .Y(_04171_));
 sky130_fd_sc_hd__nor2_1 _11033_ (.A(net234),
    .B(_03217_),
    .Y(_04172_));
 sky130_fd_sc_hd__a211o_1 _11034_ (.A1(net235),
    .A2(_03220_),
    .B1(_04172_),
    .C1(net238),
    .X(_04173_));
 sky130_fd_sc_hd__o21ai_2 _11035_ (.A1(net237),
    .A2(_02443_),
    .B1(_04173_),
    .Y(_04174_));
 sky130_fd_sc_hd__mux2_1 _11036_ (.A0(_04171_),
    .A1(_04174_),
    .S(net241),
    .X(_04175_));
 sky130_fd_sc_hd__or2_1 _11037_ (.A(\div_shifter[45] ),
    .B(_04070_),
    .X(_04176_));
 sky130_fd_sc_hd__a21oi_1 _11038_ (.A1(net245),
    .A2(_04176_),
    .B1(\div_shifter[46] ),
    .Y(_04177_));
 sky130_fd_sc_hd__a311o_1 _11039_ (.A1(\div_shifter[46] ),
    .A2(net245),
    .A3(_04176_),
    .B1(_04177_),
    .C1(net248),
    .X(_04178_));
 sky130_fd_sc_hd__or2_1 _11040_ (.A(\div_res[13] ),
    .B(_04067_),
    .X(_04179_));
 sky130_fd_sc_hd__a21oi_1 _11041_ (.A1(net24),
    .A2(_04179_),
    .B1(\div_res[14] ),
    .Y(_04180_));
 sky130_fd_sc_hd__a311o_1 _11042_ (.A1(\div_res[14] ),
    .A2(net23),
    .A3(_04179_),
    .B1(_04180_),
    .C1(net203),
    .X(_04181_));
 sky130_fd_sc_hd__nor2_1 _11043_ (.A(_06058_),
    .B(net204),
    .Y(_04182_));
 sky130_fd_sc_hd__a211o_1 _11044_ (.A1(_06058_),
    .A2(_02294_),
    .B1(_04182_),
    .C1(net205),
    .X(_04183_));
 sky130_fd_sc_hd__a22oi_2 _11045_ (.A1(_06046_),
    .A2(net212),
    .B1(_04183_),
    .B2(_06064_),
    .Y(_04184_));
 sky130_fd_sc_hd__o21a_1 _11046_ (.A1(net238),
    .A2(_02474_),
    .B1(_02312_),
    .X(_04185_));
 sky130_fd_sc_hd__inv_2 _11047_ (.A(_04185_),
    .Y(_04186_));
 sky130_fd_sc_hd__o2111a_1 _11048_ (.A1(net185),
    .A2(_04186_),
    .B1(_04184_),
    .C1(_04181_),
    .D1(_04178_),
    .X(_04187_));
 sky130_fd_sc_hd__o221a_1 _11049_ (.A1(net182),
    .A2(_04174_),
    .B1(_04175_),
    .B2(net214),
    .C1(_04187_),
    .X(_04188_));
 sky130_fd_sc_hd__a41o_1 _11050_ (.A1(_04158_),
    .A2(_04161_),
    .A3(_04166_),
    .A4(_04188_),
    .B1(net262),
    .X(_04189_));
 sky130_fd_sc_hd__and3_1 _11051_ (.A(curr_PC[13]),
    .B(curr_PC[14]),
    .C(_03973_),
    .X(_04190_));
 sky130_fd_sc_hd__a21oi_1 _11052_ (.A1(curr_PC[13]),
    .A2(_03973_),
    .B1(curr_PC[14]),
    .Y(_04191_));
 sky130_fd_sc_hd__o31ai_4 _11053_ (.A1(net257),
    .A2(_04190_),
    .A3(_04191_),
    .B1(_04189_),
    .Y(dest_val[14]));
 sky130_fd_sc_hd__o22a_1 _11054_ (.A1(net67),
    .A2(net13),
    .B1(net47),
    .B2(net64),
    .X(_04192_));
 sky130_fd_sc_hd__xnor2_1 _11055_ (.A(net108),
    .B(_04192_),
    .Y(_04193_));
 sky130_fd_sc_hd__o22a_1 _11056_ (.A1(net62),
    .A2(net41),
    .B1(net39),
    .B2(net60),
    .X(_04194_));
 sky130_fd_sc_hd__xnor2_1 _11057_ (.A(net102),
    .B(_04194_),
    .Y(_04195_));
 sky130_fd_sc_hd__nand2_1 _11058_ (.A(_04193_),
    .B(_04195_),
    .Y(_04196_));
 sky130_fd_sc_hd__xor2_1 _11059_ (.A(_04193_),
    .B(_04195_),
    .X(_04197_));
 sky130_fd_sc_hd__o22a_1 _11060_ (.A1(net57),
    .A2(net50),
    .B1(net48),
    .B2(net54),
    .X(_04198_));
 sky130_fd_sc_hd__xnor2_1 _11061_ (.A(net105),
    .B(_04198_),
    .Y(_04199_));
 sky130_fd_sc_hd__nand2_1 _11062_ (.A(_04197_),
    .B(_04199_),
    .Y(_04200_));
 sky130_fd_sc_hd__xor2_1 _11063_ (.A(_04197_),
    .B(_04199_),
    .X(_04201_));
 sky130_fd_sc_hd__nand2_1 _11064_ (.A(_04115_),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__or2_1 _11065_ (.A(_04115_),
    .B(_04201_),
    .X(_04203_));
 sky130_fd_sc_hd__nand2_1 _11066_ (.A(_04202_),
    .B(_04203_),
    .Y(_04204_));
 sky130_fd_sc_hd__o22a_1 _11067_ (.A1(net18),
    .A2(net37),
    .B1(net35),
    .B2(net16),
    .X(_04205_));
 sky130_fd_sc_hd__xnor2_1 _11068_ (.A(net136),
    .B(_04205_),
    .Y(_04206_));
 sky130_fd_sc_hd__and2b_1 _11069_ (.A_N(net154),
    .B(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__xnor2_1 _11070_ (.A(net154),
    .B(_04206_),
    .Y(_04208_));
 sky130_fd_sc_hd__o22a_1 _11071_ (.A1(net43),
    .A2(net9),
    .B1(net3),
    .B2(net95),
    .X(_04209_));
 sky130_fd_sc_hd__xnor2_1 _11072_ (.A(net139),
    .B(_04209_),
    .Y(_04210_));
 sky130_fd_sc_hd__xnor2_1 _11073_ (.A(_04208_),
    .B(_04210_),
    .Y(_04211_));
 sky130_fd_sc_hd__or2_1 _11074_ (.A(_04204_),
    .B(_04211_),
    .X(_04212_));
 sky130_fd_sc_hd__nand2_1 _11075_ (.A(_04204_),
    .B(_04211_),
    .Y(_04213_));
 sky130_fd_sc_hd__and2_1 _11076_ (.A(_04212_),
    .B(_04213_),
    .X(_04214_));
 sky130_fd_sc_hd__o22a_1 _11077_ (.A1(net118),
    .A2(net11),
    .B1(net44),
    .B2(net70),
    .X(_04215_));
 sky130_fd_sc_hd__xnor2_1 _11078_ (.A(net96),
    .B(_04215_),
    .Y(_04216_));
 sky130_fd_sc_hd__o22a_1 _11079_ (.A1(net99),
    .A2(net7),
    .B1(net5),
    .B2(net129),
    .X(_04217_));
 sky130_fd_sc_hd__xnor2_1 _11080_ (.A(net28),
    .B(_04217_),
    .Y(_04218_));
 sky130_fd_sc_hd__o22a_1 _11081_ (.A1(net76),
    .A2(net14),
    .B1(net52),
    .B2(net73),
    .X(_04219_));
 sky130_fd_sc_hd__xnor2_1 _11082_ (.A(net111),
    .B(_04219_),
    .Y(_04220_));
 sky130_fd_sc_hd__nand2b_1 _11083_ (.A_N(_04218_),
    .B(_04220_),
    .Y(_04221_));
 sky130_fd_sc_hd__nand2b_1 _11084_ (.A_N(_04220_),
    .B(_04218_),
    .Y(_04222_));
 sky130_fd_sc_hd__nand2_1 _11085_ (.A(_04221_),
    .B(_04222_),
    .Y(_04223_));
 sky130_fd_sc_hd__xor2_1 _11086_ (.A(_04216_),
    .B(_04223_),
    .X(_04224_));
 sky130_fd_sc_hd__and3_1 _11087_ (.A(_04212_),
    .B(_04213_),
    .C(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__or2_1 _11088_ (.A(_04214_),
    .B(_04224_),
    .X(_04226_));
 sky130_fd_sc_hd__nand2b_1 _11089_ (.A_N(_04225_),
    .B(_04226_),
    .Y(_04227_));
 sky130_fd_sc_hd__a21oi_1 _11090_ (.A1(_04107_),
    .A2(_04109_),
    .B1(_04105_),
    .Y(_04228_));
 sky130_fd_sc_hd__nand2_1 _11091_ (.A(_06459_),
    .B(net33),
    .Y(_04229_));
 sky130_fd_sc_hd__xnor2_1 _11092_ (.A(_04228_),
    .B(_04229_),
    .Y(_04230_));
 sky130_fd_sc_hd__nor2_1 _11093_ (.A(_04122_),
    .B(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__and2_1 _11094_ (.A(_04122_),
    .B(_04230_),
    .X(_04232_));
 sky130_fd_sc_hd__nor2_1 _11095_ (.A(_04231_),
    .B(_04232_),
    .Y(_04233_));
 sky130_fd_sc_hd__xnor2_2 _11096_ (.A(_04227_),
    .B(_04233_),
    .Y(_04234_));
 sky130_fd_sc_hd__o21a_1 _11097_ (.A1(_04091_),
    .A2(_04131_),
    .B1(_04129_),
    .X(_04235_));
 sky130_fd_sc_hd__a21bo_1 _11098_ (.A1(_04134_),
    .A2(_04138_),
    .B1_N(_04137_),
    .X(_04236_));
 sky130_fd_sc_hd__a21o_1 _11099_ (.A1(_04086_),
    .A2(_04090_),
    .B1(_04088_),
    .X(_04237_));
 sky130_fd_sc_hd__o31a_1 _11100_ (.A1(_04115_),
    .A2(_04116_),
    .A3(_04124_),
    .B1(_04126_),
    .X(_04238_));
 sky130_fd_sc_hd__a21oi_1 _11101_ (.A1(_04096_),
    .A2(_04099_),
    .B1(_04238_),
    .Y(_04239_));
 sky130_fd_sc_hd__and3_1 _11102_ (.A(_04096_),
    .B(_04099_),
    .C(_04238_),
    .X(_04240_));
 sky130_fd_sc_hd__nor2_1 _11103_ (.A(_04239_),
    .B(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__xnor2_1 _11104_ (.A(_04237_),
    .B(_04241_),
    .Y(_04242_));
 sky130_fd_sc_hd__nand2b_1 _11105_ (.A_N(_04242_),
    .B(_04236_),
    .Y(_04243_));
 sky130_fd_sc_hd__xnor2_1 _11106_ (.A(_04236_),
    .B(_04242_),
    .Y(_04244_));
 sky130_fd_sc_hd__nand2b_1 _11107_ (.A_N(_04235_),
    .B(_04244_),
    .Y(_04245_));
 sky130_fd_sc_hd__xnor2_1 _11108_ (.A(_04235_),
    .B(_04244_),
    .Y(_04246_));
 sky130_fd_sc_hd__nand2_1 _11109_ (.A(_04234_),
    .B(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__xnor2_1 _11110_ (.A(_04234_),
    .B(_04246_),
    .Y(_04248_));
 sky130_fd_sc_hd__o21a_1 _11111_ (.A1(_04133_),
    .A2(_04142_),
    .B1(_04141_),
    .X(_04249_));
 sky130_fd_sc_hd__or2_1 _11112_ (.A(_04248_),
    .B(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__xnor2_1 _11113_ (.A(_04248_),
    .B(_04249_),
    .Y(_04251_));
 sky130_fd_sc_hd__nand3_1 _11114_ (.A(_04145_),
    .B(_04148_),
    .C(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__a21o_1 _11115_ (.A1(_04145_),
    .A2(_04148_),
    .B1(_04251_),
    .X(_04253_));
 sky130_fd_sc_hd__nand2_1 _11116_ (.A(_04252_),
    .B(_04253_),
    .Y(_04254_));
 sky130_fd_sc_hd__a21oi_1 _11117_ (.A1(_04151_),
    .A2(_04154_),
    .B1(_04150_),
    .Y(_04255_));
 sky130_fd_sc_hd__xnor2_2 _11118_ (.A(_04254_),
    .B(_04255_),
    .Y(_04256_));
 sky130_fd_sc_hd__a31o_1 _11119_ (.A1(_04047_),
    .A2(_04048_),
    .A3(_04155_),
    .B1(net84),
    .X(_04257_));
 sky130_fd_sc_hd__o21ai_1 _11120_ (.A1(_04256_),
    .A2(_04257_),
    .B1(net206),
    .Y(_04258_));
 sky130_fd_sc_hd__a21oi_1 _11121_ (.A1(_04256_),
    .A2(_04257_),
    .B1(_04258_),
    .Y(_04259_));
 sky130_fd_sc_hd__or3_1 _11122_ (.A(net84),
    .B(_02184_),
    .C(_02186_),
    .X(_04260_));
 sky130_fd_sc_hd__o21ai_1 _11123_ (.A1(net84),
    .A2(_02184_),
    .B1(_02186_),
    .Y(_04261_));
 sky130_fd_sc_hd__or3_1 _11124_ (.A(_04504_),
    .B(_06052_),
    .C(_06326_),
    .X(_04262_));
 sky130_fd_sc_hd__o21a_1 _11125_ (.A1(_06070_),
    .A2(_04163_),
    .B1(_06058_),
    .X(_04263_));
 sky130_fd_sc_hd__o21a_1 _11126_ (.A1(net305),
    .A2(_04263_),
    .B1(_04262_),
    .X(_04264_));
 sky130_fd_sc_hd__a21oi_1 _11127_ (.A1(_06034_),
    .A2(_04264_),
    .B1(_02293_),
    .Y(_04265_));
 sky130_fd_sc_hd__o21a_1 _11128_ (.A1(_06034_),
    .A2(_04264_),
    .B1(_04265_),
    .X(_04266_));
 sky130_fd_sc_hd__nor2_1 _11129_ (.A(reg1_val[15]),
    .B(curr_PC[15]),
    .Y(_04267_));
 sky130_fd_sc_hd__nand2_1 _11130_ (.A(reg1_val[15]),
    .B(curr_PC[15]),
    .Y(_04268_));
 sky130_fd_sc_hd__and2b_1 _11131_ (.A_N(_04267_),
    .B(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__o21a_1 _11132_ (.A1(_04169_),
    .A2(_04170_),
    .B1(_04168_),
    .X(_04270_));
 sky130_fd_sc_hd__xnor2_1 _11133_ (.A(_04269_),
    .B(_04270_),
    .Y(_04271_));
 sky130_fd_sc_hd__mux2_1 _11134_ (.A0(_03345_),
    .A1(_03347_),
    .S(net235),
    .X(_04272_));
 sky130_fd_sc_hd__mux2_1 _11135_ (.A0(_02320_),
    .A1(_04272_),
    .S(net237),
    .X(_04273_));
 sky130_fd_sc_hd__mux2_1 _11136_ (.A0(_04271_),
    .A1(_04273_),
    .S(net241),
    .X(_04274_));
 sky130_fd_sc_hd__or2_1 _11137_ (.A(\div_shifter[46] ),
    .B(_04176_),
    .X(_04275_));
 sky130_fd_sc_hd__a21oi_1 _11138_ (.A1(net245),
    .A2(_04275_),
    .B1(\div_shifter[47] ),
    .Y(_04276_));
 sky130_fd_sc_hd__a31o_1 _11139_ (.A1(\div_shifter[47] ),
    .A2(net245),
    .A3(_04275_),
    .B1(net248),
    .X(_04277_));
 sky130_fd_sc_hd__or2_1 _11140_ (.A(\div_res[14] ),
    .B(_04179_),
    .X(_04278_));
 sky130_fd_sc_hd__a21oi_1 _11141_ (.A1(net24),
    .A2(_04278_),
    .B1(\div_res[15] ),
    .Y(_04279_));
 sky130_fd_sc_hd__a311o_1 _11142_ (.A1(\div_res[15] ),
    .A2(net24),
    .A3(_04278_),
    .B1(_04279_),
    .C1(net203),
    .X(_04280_));
 sky130_fd_sc_hd__mux2_1 _11143_ (.A0(_02300_),
    .A1(_02294_),
    .S(_06021_),
    .X(_04281_));
 sky130_fd_sc_hd__o21ai_1 _11144_ (.A1(net205),
    .A2(_04281_),
    .B1(_06028_),
    .Y(_04282_));
 sky130_fd_sc_hd__o211a_1 _11145_ (.A1(_05999_),
    .A2(_06426_),
    .B1(_04280_),
    .C1(_04282_),
    .X(_04283_));
 sky130_fd_sc_hd__o21ai_2 _11146_ (.A1(_04276_),
    .A2(_04277_),
    .B1(_04283_),
    .Y(_04284_));
 sky130_fd_sc_hd__o21a_1 _11147_ (.A1(net238),
    .A2(_02281_),
    .B1(_02312_),
    .X(_04285_));
 sky130_fd_sc_hd__a221o_1 _11148_ (.A1(_02288_),
    .A2(_04273_),
    .B1(_04285_),
    .B2(_02217_),
    .C1(_04284_),
    .X(_04286_));
 sky130_fd_sc_hd__a211o_1 _11149_ (.A1(_06412_),
    .A2(_04274_),
    .B1(_04286_),
    .C1(_04266_),
    .X(_04287_));
 sky130_fd_sc_hd__a311o_1 _11150_ (.A1(_02298_),
    .A2(_04260_),
    .A3(_04261_),
    .B1(_04287_),
    .C1(_04259_),
    .X(_04288_));
 sky130_fd_sc_hd__or2_1 _11151_ (.A(curr_PC[15]),
    .B(_04190_),
    .X(_04289_));
 sky130_fd_sc_hd__and2_1 _11152_ (.A(curr_PC[15]),
    .B(_04190_),
    .X(_04290_));
 sky130_fd_sc_hd__nor2_1 _11153_ (.A(net257),
    .B(_04290_),
    .Y(_04291_));
 sky130_fd_sc_hd__a22o_4 _11154_ (.A1(net257),
    .A2(_04288_),
    .B1(_04289_),
    .B2(_04291_),
    .X(dest_val[15]));
 sky130_fd_sc_hd__and3_1 _11155_ (.A(_04151_),
    .B(_04252_),
    .C(_04253_),
    .X(_04292_));
 sky130_fd_sc_hd__and2_2 _11156_ (.A(_04153_),
    .B(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__nand2_1 _11157_ (.A(_03935_),
    .B(_04293_),
    .Y(_04294_));
 sky130_fd_sc_hd__nand2_1 _11158_ (.A(_04152_),
    .B(_04292_),
    .Y(_04295_));
 sky130_fd_sc_hd__nand2_1 _11159_ (.A(_04150_),
    .B(_04252_),
    .Y(_04296_));
 sky130_fd_sc_hd__and3_1 _11160_ (.A(_04253_),
    .B(_04295_),
    .C(_04296_),
    .X(_04297_));
 sky130_fd_sc_hd__o31ai_2 _11161_ (.A1(_03818_),
    .A2(_03933_),
    .A3(_03934_),
    .B1(_04293_),
    .Y(_04298_));
 sky130_fd_sc_hd__o211a_2 _11162_ (.A1(_03460_),
    .A2(_04294_),
    .B1(_04297_),
    .C1(_04298_),
    .X(_04299_));
 sky130_fd_sc_hd__or4b_4 _11163_ (.A(_02923_),
    .B(_03455_),
    .C(_04294_),
    .D_N(_02035_),
    .X(_04300_));
 sky130_fd_sc_hd__nand2_1 _11164_ (.A(_04299_),
    .B(_04300_),
    .Y(_04301_));
 sky130_fd_sc_hd__a21oi_2 _11165_ (.A1(_04208_),
    .A2(_04210_),
    .B1(_04207_),
    .Y(_04302_));
 sky130_fd_sc_hd__o22a_1 _11166_ (.A1(net118),
    .A2(net7),
    .B1(net5),
    .B2(net99),
    .X(_04303_));
 sky130_fd_sc_hd__xnor2_1 _11167_ (.A(net28),
    .B(_04303_),
    .Y(_04304_));
 sky130_fd_sc_hd__xnor2_1 _11168_ (.A(_04302_),
    .B(_04304_),
    .Y(_04305_));
 sky130_fd_sc_hd__or3_1 _11169_ (.A(net129),
    .B(net28),
    .C(_04305_),
    .X(_04306_));
 sky130_fd_sc_hd__o21ai_1 _11170_ (.A1(net129),
    .A2(net28),
    .B1(_04305_),
    .Y(_04307_));
 sky130_fd_sc_hd__nand2_1 _11171_ (.A(_04306_),
    .B(_04307_),
    .Y(_04308_));
 sky130_fd_sc_hd__o22a_1 _11172_ (.A1(net54),
    .A2(net50),
    .B1(net48),
    .B2(net62),
    .X(_04309_));
 sky130_fd_sc_hd__xnor2_1 _11173_ (.A(net105),
    .B(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__o22a_1 _11174_ (.A1(net60),
    .A2(net41),
    .B1(net39),
    .B2(net18),
    .X(_04311_));
 sky130_fd_sc_hd__xnor2_1 _11175_ (.A(net102),
    .B(_04311_),
    .Y(_04312_));
 sky130_fd_sc_hd__nand2_1 _11176_ (.A(_04310_),
    .B(_04312_),
    .Y(_04313_));
 sky130_fd_sc_hd__or2_1 _11177_ (.A(_04310_),
    .B(_04312_),
    .X(_04314_));
 sky130_fd_sc_hd__nand2_1 _11178_ (.A(_04313_),
    .B(_04314_),
    .Y(_04315_));
 sky130_fd_sc_hd__a21o_1 _11179_ (.A1(_04196_),
    .A2(_04200_),
    .B1(_04315_),
    .X(_04316_));
 sky130_fd_sc_hd__nand3_1 _11180_ (.A(_04196_),
    .B(_04200_),
    .C(_04315_),
    .Y(_04317_));
 sky130_fd_sc_hd__and2_1 _11181_ (.A(_04316_),
    .B(_04317_),
    .X(_04318_));
 sky130_fd_sc_hd__o22a_1 _11182_ (.A1(net16),
    .A2(net36),
    .B1(net34),
    .B2(net9),
    .X(_04319_));
 sky130_fd_sc_hd__xnor2_1 _11183_ (.A(net135),
    .B(_04319_),
    .Y(_04320_));
 sky130_fd_sc_hd__or3_1 _11184_ (.A(net154),
    .B(_00386_),
    .C(net3),
    .X(_04321_));
 sky130_fd_sc_hd__a2bb2o_1 _11185_ (.A1_N(_00387_),
    .A2_N(net3),
    .B1(_04321_),
    .B2(net137),
    .X(_04322_));
 sky130_fd_sc_hd__nor2_1 _11186_ (.A(_04320_),
    .B(_04322_),
    .Y(_04323_));
 sky130_fd_sc_hd__and2_1 _11187_ (.A(_04320_),
    .B(_04322_),
    .X(_04324_));
 sky130_fd_sc_hd__o21ai_1 _11188_ (.A1(_04323_),
    .A2(_04324_),
    .B1(_04318_),
    .Y(_04325_));
 sky130_fd_sc_hd__or3_1 _11189_ (.A(_04318_),
    .B(_04323_),
    .C(_04324_),
    .X(_04326_));
 sky130_fd_sc_hd__nand2_1 _11190_ (.A(_04325_),
    .B(_04326_),
    .Y(_04327_));
 sky130_fd_sc_hd__o22a_1 _11191_ (.A1(net70),
    .A2(net11),
    .B1(net44),
    .B2(net76),
    .X(_04328_));
 sky130_fd_sc_hd__xnor2_1 _11192_ (.A(net96),
    .B(_04328_),
    .Y(_04329_));
 sky130_fd_sc_hd__inv_2 _11193_ (.A(_04329_),
    .Y(_04330_));
 sky130_fd_sc_hd__o22a_1 _11194_ (.A1(net64),
    .A2(net13),
    .B1(net47),
    .B2(net57),
    .X(_04331_));
 sky130_fd_sc_hd__xnor2_1 _11195_ (.A(net108),
    .B(_04331_),
    .Y(_04332_));
 sky130_fd_sc_hd__xor2_1 _11196_ (.A(_04329_),
    .B(_04332_),
    .X(_04333_));
 sky130_fd_sc_hd__o22a_1 _11197_ (.A1(net73),
    .A2(net14),
    .B1(net52),
    .B2(net67),
    .X(_04334_));
 sky130_fd_sc_hd__xnor2_1 _11198_ (.A(net111),
    .B(_04334_),
    .Y(_04335_));
 sky130_fd_sc_hd__and2b_1 _11199_ (.A_N(_04333_),
    .B(_04335_),
    .X(_04336_));
 sky130_fd_sc_hd__and2b_1 _11200_ (.A_N(_04335_),
    .B(_04333_),
    .X(_04337_));
 sky130_fd_sc_hd__or2_1 _11201_ (.A(_04336_),
    .B(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__nor2_1 _11202_ (.A(_04327_),
    .B(_04338_),
    .Y(_04339_));
 sky130_fd_sc_hd__and2_1 _11203_ (.A(_04327_),
    .B(_04338_),
    .X(_04341_));
 sky130_fd_sc_hd__or2_1 _11204_ (.A(_04339_),
    .B(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__nor2_1 _11205_ (.A(_04308_),
    .B(_04342_),
    .Y(_04343_));
 sky130_fd_sc_hd__and2_1 _11206_ (.A(_04308_),
    .B(_04342_),
    .X(_04344_));
 sky130_fd_sc_hd__nor2_1 _11207_ (.A(_04343_),
    .B(_04344_),
    .Y(_04345_));
 sky130_fd_sc_hd__a21o_1 _11208_ (.A1(_04226_),
    .A2(_04233_),
    .B1(_04225_),
    .X(_04346_));
 sky130_fd_sc_hd__o21bai_1 _11209_ (.A1(_04228_),
    .A2(_04229_),
    .B1_N(_04231_),
    .Y(_04347_));
 sky130_fd_sc_hd__o21a_1 _11210_ (.A1(_04216_),
    .A2(_04223_),
    .B1(_04221_),
    .X(_04348_));
 sky130_fd_sc_hd__a21oi_1 _11211_ (.A1(_04202_),
    .A2(_04212_),
    .B1(_04348_),
    .Y(_04349_));
 sky130_fd_sc_hd__and3_1 _11212_ (.A(_04202_),
    .B(_04212_),
    .C(_04348_),
    .X(_04350_));
 sky130_fd_sc_hd__nor2_1 _11213_ (.A(_04349_),
    .B(_04350_),
    .Y(_04352_));
 sky130_fd_sc_hd__xnor2_1 _11214_ (.A(_04347_),
    .B(_04352_),
    .Y(_04353_));
 sky130_fd_sc_hd__a21oi_1 _11215_ (.A1(_04237_),
    .A2(_04241_),
    .B1(_04239_),
    .Y(_04354_));
 sky130_fd_sc_hd__xnor2_1 _11216_ (.A(_04353_),
    .B(_04354_),
    .Y(_04355_));
 sky130_fd_sc_hd__and2b_1 _11217_ (.A_N(_04355_),
    .B(_04346_),
    .X(_04356_));
 sky130_fd_sc_hd__xnor2_1 _11218_ (.A(_04346_),
    .B(_04355_),
    .Y(_04357_));
 sky130_fd_sc_hd__and2_1 _11219_ (.A(_04345_),
    .B(_04357_),
    .X(_04358_));
 sky130_fd_sc_hd__nor2_1 _11220_ (.A(_04345_),
    .B(_04357_),
    .Y(_04359_));
 sky130_fd_sc_hd__or2_1 _11221_ (.A(_04358_),
    .B(_04359_),
    .X(_04360_));
 sky130_fd_sc_hd__a21oi_1 _11222_ (.A1(_04243_),
    .A2(_04245_),
    .B1(_04360_),
    .Y(_04361_));
 sky130_fd_sc_hd__and3_1 _11223_ (.A(_04243_),
    .B(_04245_),
    .C(_04360_),
    .X(_04363_));
 sky130_fd_sc_hd__or2_1 _11224_ (.A(_04361_),
    .B(_04363_),
    .X(_04364_));
 sky130_fd_sc_hd__a21o_1 _11225_ (.A1(_04247_),
    .A2(_04250_),
    .B1(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__nand3_1 _11226_ (.A(_04247_),
    .B(_04250_),
    .C(_04364_),
    .Y(_04366_));
 sky130_fd_sc_hd__and2_1 _11227_ (.A(_04365_),
    .B(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__a21bo_1 _11228_ (.A1(_04299_),
    .A2(_04300_),
    .B1_N(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__xnor2_2 _11229_ (.A(_04301_),
    .B(_04367_),
    .Y(_04369_));
 sky130_fd_sc_hd__and4_1 _11230_ (.A(_03822_),
    .B(_03937_),
    .C(_04047_),
    .D(_04155_),
    .X(_04370_));
 sky130_fd_sc_hd__and4b_4 _11231_ (.A_N(_03591_),
    .B(_03823_),
    .C(_04256_),
    .D(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__or2_1 _11232_ (.A(net84),
    .B(_04371_),
    .X(_04372_));
 sky130_fd_sc_hd__nand2_1 _11233_ (.A(_04369_),
    .B(_04372_),
    .Y(_04374_));
 sky130_fd_sc_hd__o21a_1 _11234_ (.A1(_04369_),
    .A2(_04372_),
    .B1(net206),
    .X(_04375_));
 sky130_fd_sc_hd__nor2_1 _11235_ (.A(_02137_),
    .B(_02187_),
    .Y(_04376_));
 sky130_fd_sc_hd__xnor2_1 _11236_ (.A(_02154_),
    .B(_04376_),
    .Y(_04377_));
 sky130_fd_sc_hd__o21ai_1 _11237_ (.A1(_06034_),
    .A2(_04263_),
    .B1(_06021_),
    .Y(_04378_));
 sky130_fd_sc_hd__nand3_1 _11238_ (.A(net305),
    .B(_06010_),
    .C(_06327_),
    .Y(_04379_));
 sky130_fd_sc_hd__a21boi_1 _11239_ (.A1(_04504_),
    .A2(_04378_),
    .B1_N(_04379_),
    .Y(_04380_));
 sky130_fd_sc_hd__nand2_1 _11240_ (.A(_05966_),
    .B(_04380_),
    .Y(_04381_));
 sky130_fd_sc_hd__o21a_1 _11241_ (.A1(_05966_),
    .A2(_04380_),
    .B1(net251),
    .X(_04382_));
 sky130_fd_sc_hd__o21a_1 _11242_ (.A1(_04267_),
    .A2(_04270_),
    .B1(_04268_),
    .X(_04383_));
 sky130_fd_sc_hd__nor2_1 _11243_ (.A(reg1_val[16]),
    .B(curr_PC[16]),
    .Y(_04385_));
 sky130_fd_sc_hd__nand2_1 _11244_ (.A(reg1_val[16]),
    .B(curr_PC[16]),
    .Y(_04386_));
 sky130_fd_sc_hd__and2b_1 _11245_ (.A_N(_04385_),
    .B(_04386_),
    .X(_04387_));
 sky130_fd_sc_hd__xnor2_1 _11246_ (.A(_04383_),
    .B(_04387_),
    .Y(_04388_));
 sky130_fd_sc_hd__or2_1 _11247_ (.A(net263),
    .B(_04285_),
    .X(_04389_));
 sky130_fd_sc_hd__o211a_1 _11248_ (.A1(net241),
    .A2(_04388_),
    .B1(_04389_),
    .C1(_06412_),
    .X(_04390_));
 sky130_fd_sc_hd__or2_1 _11249_ (.A(\div_res[15] ),
    .B(_04278_),
    .X(_04391_));
 sky130_fd_sc_hd__a21oi_1 _11250_ (.A1(net23),
    .A2(_04391_),
    .B1(\div_res[16] ),
    .Y(_04392_));
 sky130_fd_sc_hd__a31o_1 _11251_ (.A1(\div_res[16] ),
    .A2(net23),
    .A3(_04391_),
    .B1(net202),
    .X(_04393_));
 sky130_fd_sc_hd__or2_1 _11252_ (.A(\div_shifter[47] ),
    .B(_04275_),
    .X(_04394_));
 sky130_fd_sc_hd__a21oi_1 _11253_ (.A1(net245),
    .A2(_04394_),
    .B1(\div_shifter[48] ),
    .Y(_04396_));
 sky130_fd_sc_hd__a311o_1 _11254_ (.A1(\div_shifter[48] ),
    .A2(net245),
    .A3(_04394_),
    .B1(_04396_),
    .C1(net248),
    .X(_04397_));
 sky130_fd_sc_hd__o21ai_1 _11255_ (.A1(_05944_),
    .A2(_02295_),
    .B1(_02291_),
    .Y(_04398_));
 sky130_fd_sc_hd__a22o_1 _11256_ (.A1(_05911_),
    .A2(net212),
    .B1(_02300_),
    .B2(_05944_),
    .X(_04399_));
 sky130_fd_sc_hd__a21oi_2 _11257_ (.A1(_05955_),
    .A2(_04398_),
    .B1(_04399_),
    .Y(_04400_));
 sky130_fd_sc_hd__o211ai_2 _11258_ (.A1(_04392_),
    .A2(_04393_),
    .B1(_04397_),
    .C1(_04400_),
    .Y(_04401_));
 sky130_fd_sc_hd__a221o_1 _11259_ (.A1(_02217_),
    .A2(_04273_),
    .B1(_04285_),
    .B2(_02288_),
    .C1(_04401_),
    .X(_04402_));
 sky130_fd_sc_hd__a211o_1 _11260_ (.A1(_04381_),
    .A2(_04382_),
    .B1(_04390_),
    .C1(_04402_),
    .X(_04403_));
 sky130_fd_sc_hd__a221o_1 _11261_ (.A1(_04374_),
    .A2(_04375_),
    .B1(_04377_),
    .B2(_02298_),
    .C1(_04403_),
    .X(_04404_));
 sky130_fd_sc_hd__nand2_1 _11262_ (.A(curr_PC[16]),
    .B(_04290_),
    .Y(_04405_));
 sky130_fd_sc_hd__o21a_1 _11263_ (.A1(curr_PC[16]),
    .A2(_04290_),
    .B1(net262),
    .X(_04407_));
 sky130_fd_sc_hd__a22o_4 _11264_ (.A1(net258),
    .A2(_04404_),
    .B1(_04405_),
    .B2(_04407_),
    .X(dest_val[16]));
 sky130_fd_sc_hd__and3_1 _11265_ (.A(curr_PC[16]),
    .B(curr_PC[17]),
    .C(_04290_),
    .X(_04408_));
 sky130_fd_sc_hd__a21oi_1 _11266_ (.A1(curr_PC[16]),
    .A2(_04290_),
    .B1(curr_PC[17]),
    .Y(_04409_));
 sky130_fd_sc_hd__o21a_1 _11267_ (.A1(_04408_),
    .A2(_04409_),
    .B1(net262),
    .X(_04410_));
 sky130_fd_sc_hd__o22a_1 _11268_ (.A1(net18),
    .A2(net40),
    .B1(net38),
    .B2(net16),
    .X(_04411_));
 sky130_fd_sc_hd__xor2_1 _11269_ (.A(net102),
    .B(_04411_),
    .X(_04412_));
 sky130_fd_sc_hd__or2_1 _11270_ (.A(net137),
    .B(_04412_),
    .X(_04413_));
 sky130_fd_sc_hd__xnor2_1 _11271_ (.A(net137),
    .B(_04412_),
    .Y(_04414_));
 sky130_fd_sc_hd__o22a_1 _11272_ (.A1(net9),
    .A2(net36),
    .B1(net34),
    .B2(net3),
    .X(_04415_));
 sky130_fd_sc_hd__xnor2_1 _11273_ (.A(_00436_),
    .B(_04415_),
    .Y(_04417_));
 sky130_fd_sc_hd__or2_1 _11274_ (.A(_04414_),
    .B(_04417_),
    .X(_04418_));
 sky130_fd_sc_hd__nand2_1 _11275_ (.A(_04414_),
    .B(_04417_),
    .Y(_04419_));
 sky130_fd_sc_hd__nand2_1 _11276_ (.A(_04418_),
    .B(_04419_),
    .Y(_04420_));
 sky130_fd_sc_hd__nor2_1 _11277_ (.A(_04323_),
    .B(_04420_),
    .Y(_04421_));
 sky130_fd_sc_hd__and2_1 _11278_ (.A(_04323_),
    .B(_04420_),
    .X(_04422_));
 sky130_fd_sc_hd__nor2_1 _11279_ (.A(_04421_),
    .B(_04422_),
    .Y(_04423_));
 sky130_fd_sc_hd__xnor2_1 _11280_ (.A(_04313_),
    .B(_04423_),
    .Y(_04424_));
 sky130_fd_sc_hd__o22a_1 _11281_ (.A1(net67),
    .A2(net14),
    .B1(net52),
    .B2(net64),
    .X(_04425_));
 sky130_fd_sc_hd__xnor2_1 _11282_ (.A(net111),
    .B(_04425_),
    .Y(_04426_));
 sky130_fd_sc_hd__o22a_1 _11283_ (.A1(net62),
    .A2(net50),
    .B1(net48),
    .B2(net60),
    .X(_04428_));
 sky130_fd_sc_hd__xnor2_1 _11284_ (.A(net105),
    .B(_04428_),
    .Y(_04429_));
 sky130_fd_sc_hd__and2_1 _11285_ (.A(_04426_),
    .B(_04429_),
    .X(_04430_));
 sky130_fd_sc_hd__nor2_1 _11286_ (.A(_04426_),
    .B(_04429_),
    .Y(_04431_));
 sky130_fd_sc_hd__nor2_1 _11287_ (.A(_04430_),
    .B(_04431_),
    .Y(_04432_));
 sky130_fd_sc_hd__o22a_1 _11288_ (.A1(net57),
    .A2(net13),
    .B1(net47),
    .B2(net54),
    .X(_04433_));
 sky130_fd_sc_hd__xnor2_1 _11289_ (.A(net108),
    .B(_04433_),
    .Y(_04434_));
 sky130_fd_sc_hd__and2_1 _11290_ (.A(_04432_),
    .B(_04434_),
    .X(_04435_));
 sky130_fd_sc_hd__nor2_1 _11291_ (.A(_04432_),
    .B(_04434_),
    .Y(_04436_));
 sky130_fd_sc_hd__nor2_1 _11292_ (.A(_04435_),
    .B(_04436_),
    .Y(_04437_));
 sky130_fd_sc_hd__and2_1 _11293_ (.A(_04424_),
    .B(_04437_),
    .X(_04439_));
 sky130_fd_sc_hd__nor2_1 _11294_ (.A(_04424_),
    .B(_04437_),
    .Y(_04440_));
 sky130_fd_sc_hd__o22a_1 _11295_ (.A1(net70),
    .A2(net7),
    .B1(net5),
    .B2(net118),
    .X(_04441_));
 sky130_fd_sc_hd__xnor2_1 _11296_ (.A(net28),
    .B(_04441_),
    .Y(_04442_));
 sky130_fd_sc_hd__nor2_1 _11297_ (.A(net99),
    .B(net29),
    .Y(_04443_));
 sky130_fd_sc_hd__o22a_1 _11298_ (.A1(net76),
    .A2(net11),
    .B1(net44),
    .B2(net73),
    .X(_04444_));
 sky130_fd_sc_hd__xor2_1 _11299_ (.A(net96),
    .B(_04444_),
    .X(_04445_));
 sky130_fd_sc_hd__nand2_1 _11300_ (.A(_04443_),
    .B(_04445_),
    .Y(_04446_));
 sky130_fd_sc_hd__or2_1 _11301_ (.A(_04443_),
    .B(_04445_),
    .X(_04447_));
 sky130_fd_sc_hd__nand2_1 _11302_ (.A(_04446_),
    .B(_04447_),
    .Y(_04448_));
 sky130_fd_sc_hd__xnor2_1 _11303_ (.A(_04442_),
    .B(_04448_),
    .Y(_04450_));
 sky130_fd_sc_hd__or3_1 _11304_ (.A(_04439_),
    .B(_04440_),
    .C(_04450_),
    .X(_04451_));
 sky130_fd_sc_hd__o21ai_1 _11305_ (.A1(_04439_),
    .A2(_04440_),
    .B1(_04450_),
    .Y(_04452_));
 sky130_fd_sc_hd__nand2_1 _11306_ (.A(_04451_),
    .B(_04452_),
    .Y(_04453_));
 sky130_fd_sc_hd__o21ai_1 _11307_ (.A1(_04302_),
    .A2(_04304_),
    .B1(_04306_),
    .Y(_04454_));
 sky130_fd_sc_hd__nand2_1 _11308_ (.A(_04316_),
    .B(_04325_),
    .Y(_04455_));
 sky130_fd_sc_hd__a21oi_1 _11309_ (.A1(_04330_),
    .A2(_04332_),
    .B1(_04336_),
    .Y(_04456_));
 sky130_fd_sc_hd__inv_2 _11310_ (.A(_04456_),
    .Y(_04457_));
 sky130_fd_sc_hd__nand2_1 _11311_ (.A(_04455_),
    .B(_04457_),
    .Y(_04458_));
 sky130_fd_sc_hd__xnor2_1 _11312_ (.A(_04455_),
    .B(_04457_),
    .Y(_04459_));
 sky130_fd_sc_hd__nand2b_1 _11313_ (.A_N(_04459_),
    .B(_04454_),
    .Y(_04461_));
 sky130_fd_sc_hd__xor2_1 _11314_ (.A(_04454_),
    .B(_04459_),
    .X(_04462_));
 sky130_fd_sc_hd__a21o_1 _11315_ (.A1(_04347_),
    .A2(_04352_),
    .B1(_04349_),
    .X(_04463_));
 sky130_fd_sc_hd__and2b_1 _11316_ (.A_N(_04462_),
    .B(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__xnor2_1 _11317_ (.A(_04462_),
    .B(_04463_),
    .Y(_04465_));
 sky130_fd_sc_hd__o21a_1 _11318_ (.A1(_04339_),
    .A2(_04343_),
    .B1(_04465_),
    .X(_04466_));
 sky130_fd_sc_hd__nor3_1 _11319_ (.A(_04339_),
    .B(_04343_),
    .C(_04465_),
    .Y(_04467_));
 sky130_fd_sc_hd__or2_1 _11320_ (.A(_04466_),
    .B(_04467_),
    .X(_04468_));
 sky130_fd_sc_hd__xor2_1 _11321_ (.A(_04453_),
    .B(_04468_),
    .X(_04469_));
 sky130_fd_sc_hd__o21ba_1 _11322_ (.A1(_04353_),
    .A2(_04354_),
    .B1_N(_04356_),
    .X(_04470_));
 sky130_fd_sc_hd__nand2b_1 _11323_ (.A_N(_04470_),
    .B(_04469_),
    .Y(_04472_));
 sky130_fd_sc_hd__xnor2_1 _11324_ (.A(_04469_),
    .B(_04470_),
    .Y(_04473_));
 sky130_fd_sc_hd__o21ai_1 _11325_ (.A1(_04358_),
    .A2(_04361_),
    .B1(_04473_),
    .Y(_04474_));
 sky130_fd_sc_hd__inv_2 _11326_ (.A(_04474_),
    .Y(_04475_));
 sky130_fd_sc_hd__nor3_1 _11327_ (.A(_04358_),
    .B(_04361_),
    .C(_04473_),
    .Y(_04476_));
 sky130_fd_sc_hd__nor2_1 _11328_ (.A(_04475_),
    .B(_04476_),
    .Y(_04477_));
 sky130_fd_sc_hd__nand3_1 _11329_ (.A(_04365_),
    .B(_04368_),
    .C(_04477_),
    .Y(_04478_));
 sky130_fd_sc_hd__a21o_1 _11330_ (.A1(_04365_),
    .A2(_04368_),
    .B1(_04477_),
    .X(_04479_));
 sky130_fd_sc_hd__and2_1 _11331_ (.A(_04478_),
    .B(_04479_),
    .X(_04480_));
 sky130_fd_sc_hd__a21o_1 _11332_ (.A1(_04369_),
    .A2(_04371_),
    .B1(net84),
    .X(_04481_));
 sky130_fd_sc_hd__o21ai_1 _11333_ (.A1(_04480_),
    .A2(_04481_),
    .B1(net206),
    .Y(_04483_));
 sky130_fd_sc_hd__a21o_1 _11334_ (.A1(_04480_),
    .A2(_04481_),
    .B1(_04483_),
    .X(_04484_));
 sky130_fd_sc_hd__a21oi_1 _11335_ (.A1(net20),
    .A2(_02188_),
    .B1(_02190_),
    .Y(_04485_));
 sky130_fd_sc_hd__a31o_1 _11336_ (.A1(net20),
    .A2(_02188_),
    .A3(_02190_),
    .B1(net250),
    .X(_04486_));
 sky130_fd_sc_hd__a21o_1 _11337_ (.A1(_05955_),
    .A2(_04378_),
    .B1(_05944_),
    .X(_04487_));
 sky130_fd_sc_hd__mux2_1 _11338_ (.A0(_06329_),
    .A1(_04487_),
    .S(net299),
    .X(_04488_));
 sky130_fd_sc_hd__nor2_1 _11339_ (.A(_05887_),
    .B(_04488_),
    .Y(_04489_));
 sky130_fd_sc_hd__a21o_1 _11340_ (.A1(_05887_),
    .A2(_04488_),
    .B1(_02293_),
    .X(_04490_));
 sky130_fd_sc_hd__o21a_1 _11341_ (.A1(_04383_),
    .A2(_04385_),
    .B1(_04386_),
    .X(_04491_));
 sky130_fd_sc_hd__nor2_1 _11342_ (.A(reg1_val[17]),
    .B(curr_PC[17]),
    .Y(_04492_));
 sky130_fd_sc_hd__nand2_1 _11343_ (.A(reg1_val[17]),
    .B(curr_PC[17]),
    .Y(_04494_));
 sky130_fd_sc_hd__nand2b_1 _11344_ (.A_N(_04492_),
    .B(_04494_),
    .Y(_04495_));
 sky130_fd_sc_hd__xnor2_1 _11345_ (.A(_04491_),
    .B(_04495_),
    .Y(_04496_));
 sky130_fd_sc_hd__nor2_1 _11346_ (.A(net263),
    .B(_04185_),
    .Y(_04497_));
 sky130_fd_sc_hd__a211o_1 _11347_ (.A1(net263),
    .A2(_04496_),
    .B1(_04497_),
    .C1(net214),
    .X(_04498_));
 sky130_fd_sc_hd__or2_1 _11348_ (.A(\div_res[16] ),
    .B(_04391_),
    .X(_04499_));
 sky130_fd_sc_hd__a21oi_1 _11349_ (.A1(net23),
    .A2(_04499_),
    .B1(\div_res[17] ),
    .Y(_04500_));
 sky130_fd_sc_hd__a311o_1 _11350_ (.A1(\div_res[17] ),
    .A2(net23),
    .A3(_04499_),
    .B1(_04500_),
    .C1(net202),
    .X(_04501_));
 sky130_fd_sc_hd__o21a_1 _11351_ (.A1(_05868_),
    .A2(_02295_),
    .B1(_02291_),
    .X(_04502_));
 sky130_fd_sc_hd__a221oi_1 _11352_ (.A1(_05840_),
    .A2(net212),
    .B1(_02300_),
    .B2(_05868_),
    .C1(_06390_),
    .Y(_04503_));
 sky130_fd_sc_hd__o211a_1 _11353_ (.A1(_05875_),
    .A2(_04502_),
    .B1(_04503_),
    .C1(_04501_),
    .X(_04505_));
 sky130_fd_sc_hd__or2_1 _11354_ (.A(\div_shifter[48] ),
    .B(_04394_),
    .X(_04506_));
 sky130_fd_sc_hd__a21oi_1 _11355_ (.A1(net244),
    .A2(_04506_),
    .B1(\div_shifter[49] ),
    .Y(_04507_));
 sky130_fd_sc_hd__a31o_1 _11356_ (.A1(\div_shifter[49] ),
    .A2(net244),
    .A3(_04506_),
    .B1(net248),
    .X(_04508_));
 sky130_fd_sc_hd__o22a_1 _11357_ (.A1(net183),
    .A2(_04186_),
    .B1(_04507_),
    .B2(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__o211a_1 _11358_ (.A1(net186),
    .A2(_04174_),
    .B1(_04505_),
    .C1(_04509_),
    .X(_04510_));
 sky130_fd_sc_hd__o211a_1 _11359_ (.A1(_04489_),
    .A2(_04490_),
    .B1(_04498_),
    .C1(_04510_),
    .X(_04511_));
 sky130_fd_sc_hd__o21a_1 _11360_ (.A1(_04485_),
    .A2(_04486_),
    .B1(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__a21oi_4 _11361_ (.A1(_04484_),
    .A2(_04512_),
    .B1(_04410_),
    .Y(dest_val[17]));
 sky130_fd_sc_hd__o21ai_1 _11362_ (.A1(_04453_),
    .A2(_04468_),
    .B1(_04472_),
    .Y(_04513_));
 sky130_fd_sc_hd__o22a_1 _11363_ (.A1(net73),
    .A2(net11),
    .B1(net44),
    .B2(net67),
    .X(_04515_));
 sky130_fd_sc_hd__xnor2_1 _11364_ (.A(net96),
    .B(_04515_),
    .Y(_04516_));
 sky130_fd_sc_hd__o22a_1 _11365_ (.A1(net77),
    .A2(net7),
    .B1(net5),
    .B2(net71),
    .X(_04517_));
 sky130_fd_sc_hd__xnor2_1 _11366_ (.A(net33),
    .B(_04517_),
    .Y(_04518_));
 sky130_fd_sc_hd__o22a_1 _11367_ (.A1(net64),
    .A2(net14),
    .B1(net52),
    .B2(net57),
    .X(_04519_));
 sky130_fd_sc_hd__xnor2_1 _11368_ (.A(net111),
    .B(_04519_),
    .Y(_04520_));
 sky130_fd_sc_hd__nand2_1 _11369_ (.A(_04518_),
    .B(_04520_),
    .Y(_04521_));
 sky130_fd_sc_hd__or2_1 _11370_ (.A(_04518_),
    .B(_04520_),
    .X(_04522_));
 sky130_fd_sc_hd__nand2_1 _11371_ (.A(_04521_),
    .B(_04522_),
    .Y(_04523_));
 sky130_fd_sc_hd__xnor2_1 _11372_ (.A(_04516_),
    .B(_04523_),
    .Y(_04524_));
 sky130_fd_sc_hd__o22a_1 _11373_ (.A1(net55),
    .A2(net13),
    .B1(net47),
    .B2(net63),
    .X(_04526_));
 sky130_fd_sc_hd__xnor2_1 _11374_ (.A(net108),
    .B(_04526_),
    .Y(_04527_));
 sky130_fd_sc_hd__o22a_1 _11375_ (.A1(net17),
    .A2(net40),
    .B1(net38),
    .B2(net10),
    .X(_04528_));
 sky130_fd_sc_hd__xnor2_1 _11376_ (.A(net102),
    .B(_04528_),
    .Y(_04529_));
 sky130_fd_sc_hd__nand2_1 _11377_ (.A(_04527_),
    .B(_04529_),
    .Y(_04530_));
 sky130_fd_sc_hd__or2_1 _11378_ (.A(_04527_),
    .B(_04529_),
    .X(_04531_));
 sky130_fd_sc_hd__and2_1 _11379_ (.A(_04530_),
    .B(_04531_),
    .X(_04532_));
 sky130_fd_sc_hd__o22a_1 _11380_ (.A1(net61),
    .A2(net50),
    .B1(net48),
    .B2(net18),
    .X(_04533_));
 sky130_fd_sc_hd__xnor2_1 _11381_ (.A(net105),
    .B(_04533_),
    .Y(_04534_));
 sky130_fd_sc_hd__nand2_1 _11382_ (.A(_04532_),
    .B(_04534_),
    .Y(_04535_));
 sky130_fd_sc_hd__or2_1 _11383_ (.A(_04532_),
    .B(_04534_),
    .X(_04537_));
 sky130_fd_sc_hd__and2_1 _11384_ (.A(_04535_),
    .B(_04537_),
    .X(_04538_));
 sky130_fd_sc_hd__nand2_1 _11385_ (.A(_00454_),
    .B(_00756_),
    .Y(_04539_));
 sky130_fd_sc_hd__a22o_1 _11386_ (.A1(_00453_),
    .A2(_00756_),
    .B1(_04539_),
    .B2(net135),
    .X(_04540_));
 sky130_fd_sc_hd__or2_1 _11387_ (.A(net119),
    .B(net29),
    .X(_04541_));
 sky130_fd_sc_hd__xnor2_1 _11388_ (.A(_04540_),
    .B(_04541_),
    .Y(_04542_));
 sky130_fd_sc_hd__a21o_1 _11389_ (.A1(_04413_),
    .A2(_04418_),
    .B1(_04542_),
    .X(_04543_));
 sky130_fd_sc_hd__nand3_1 _11390_ (.A(_04413_),
    .B(_04418_),
    .C(_04542_),
    .Y(_04544_));
 sky130_fd_sc_hd__and2_1 _11391_ (.A(_04543_),
    .B(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__nand2_1 _11392_ (.A(_04538_),
    .B(_04545_),
    .Y(_04546_));
 sky130_fd_sc_hd__or2_1 _11393_ (.A(_04538_),
    .B(_04545_),
    .X(_04547_));
 sky130_fd_sc_hd__nand2_1 _11394_ (.A(_04546_),
    .B(_04547_),
    .Y(_04548_));
 sky130_fd_sc_hd__xnor2_1 _11395_ (.A(_04524_),
    .B(_04548_),
    .Y(_04549_));
 sky130_fd_sc_hd__nand2b_1 _11396_ (.A_N(_04439_),
    .B(_04451_),
    .Y(_04550_));
 sky130_fd_sc_hd__o21ai_1 _11397_ (.A1(_04442_),
    .A2(_04448_),
    .B1(_04446_),
    .Y(_04551_));
 sky130_fd_sc_hd__a31o_1 _11398_ (.A1(_04310_),
    .A2(_04312_),
    .A3(_04423_),
    .B1(_04421_),
    .X(_04552_));
 sky130_fd_sc_hd__nor2_1 _11399_ (.A(_04430_),
    .B(_04435_),
    .Y(_04553_));
 sky130_fd_sc_hd__o21ai_1 _11400_ (.A1(_04430_),
    .A2(_04435_),
    .B1(_04552_),
    .Y(_04554_));
 sky130_fd_sc_hd__xnor2_1 _11401_ (.A(_04552_),
    .B(_04553_),
    .Y(_04555_));
 sky130_fd_sc_hd__xnor2_1 _11402_ (.A(_04551_),
    .B(_04555_),
    .Y(_04556_));
 sky130_fd_sc_hd__a21o_1 _11403_ (.A1(_04458_),
    .A2(_04461_),
    .B1(_04556_),
    .X(_04557_));
 sky130_fd_sc_hd__nand3_1 _11404_ (.A(_04458_),
    .B(_04461_),
    .C(_04556_),
    .Y(_04558_));
 sky130_fd_sc_hd__and2_1 _11405_ (.A(_04557_),
    .B(_04558_),
    .X(_04559_));
 sky130_fd_sc_hd__nand2_1 _11406_ (.A(_04550_),
    .B(_04559_),
    .Y(_04560_));
 sky130_fd_sc_hd__xnor2_1 _11407_ (.A(_04550_),
    .B(_04559_),
    .Y(_04561_));
 sky130_fd_sc_hd__or2_1 _11408_ (.A(_04549_),
    .B(_04561_),
    .X(_04562_));
 sky130_fd_sc_hd__nand2_1 _11409_ (.A(_04549_),
    .B(_04561_),
    .Y(_04563_));
 sky130_fd_sc_hd__and2_1 _11410_ (.A(_04562_),
    .B(_04563_),
    .X(_04564_));
 sky130_fd_sc_hd__o21ai_1 _11411_ (.A1(_04464_),
    .A2(_04466_),
    .B1(_04564_),
    .Y(_04565_));
 sky130_fd_sc_hd__or3_1 _11412_ (.A(_04464_),
    .B(_04466_),
    .C(_04564_),
    .X(_04566_));
 sky130_fd_sc_hd__nand2_1 _11413_ (.A(_04565_),
    .B(_04566_),
    .Y(_04568_));
 sky130_fd_sc_hd__and3_1 _11414_ (.A(_04513_),
    .B(_04565_),
    .C(_04566_),
    .X(_04569_));
 sky130_fd_sc_hd__inv_2 _11415_ (.A(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__xor2_1 _11416_ (.A(_04513_),
    .B(_04568_),
    .X(_04571_));
 sky130_fd_sc_hd__a21o_1 _11417_ (.A1(_04365_),
    .A2(_04474_),
    .B1(_04476_),
    .X(_04572_));
 sky130_fd_sc_hd__nand2_1 _11418_ (.A(_04367_),
    .B(_04477_),
    .Y(_04573_));
 sky130_fd_sc_hd__a21o_1 _11419_ (.A1(_04299_),
    .A2(_04300_),
    .B1(_04573_),
    .X(_04574_));
 sky130_fd_sc_hd__a21oi_1 _11420_ (.A1(_04572_),
    .A2(_04574_),
    .B1(_04571_),
    .Y(_04575_));
 sky130_fd_sc_hd__and3_1 _11421_ (.A(_04571_),
    .B(_04572_),
    .C(_04574_),
    .X(_04576_));
 sky130_fd_sc_hd__or2_1 _11422_ (.A(_04575_),
    .B(_04576_),
    .X(_04577_));
 sky130_fd_sc_hd__a31o_1 _11423_ (.A1(_04369_),
    .A2(_04371_),
    .A3(_04480_),
    .B1(_02137_),
    .X(_04579_));
 sky130_fd_sc_hd__or2_1 _11424_ (.A(_04577_),
    .B(_04579_),
    .X(_04580_));
 sky130_fd_sc_hd__a21oi_1 _11425_ (.A1(_04577_),
    .A2(_04579_),
    .B1(_02214_),
    .Y(_04581_));
 sky130_fd_sc_hd__and3_1 _11426_ (.A(net20),
    .B(_02153_),
    .C(_02191_),
    .X(_04582_));
 sky130_fd_sc_hd__a21oi_1 _11427_ (.A1(net20),
    .A2(_02191_),
    .B1(_02153_),
    .Y(_04583_));
 sky130_fd_sc_hd__nor2_1 _11428_ (.A(_04582_),
    .B(_04583_),
    .Y(_04584_));
 sky130_fd_sc_hd__a21o_1 _11429_ (.A1(_05881_),
    .A2(_04487_),
    .B1(_05868_),
    .X(_04585_));
 sky130_fd_sc_hd__mux2_1 _11430_ (.A0(_06331_),
    .A1(_04585_),
    .S(net299),
    .X(_04586_));
 sky130_fd_sc_hd__nand2_1 _11431_ (.A(_05814_),
    .B(_04586_),
    .Y(_04587_));
 sky130_fd_sc_hd__o211a_1 _11432_ (.A1(_05814_),
    .A2(_04586_),
    .B1(_04587_),
    .C1(net251),
    .X(_04588_));
 sky130_fd_sc_hd__nor2_1 _11433_ (.A(reg1_val[18]),
    .B(curr_PC[18]),
    .Y(_04590_));
 sky130_fd_sc_hd__nand2_1 _11434_ (.A(reg1_val[18]),
    .B(curr_PC[18]),
    .Y(_04591_));
 sky130_fd_sc_hd__and2b_1 _11435_ (.A_N(_04590_),
    .B(_04591_),
    .X(_04592_));
 sky130_fd_sc_hd__o21a_1 _11436_ (.A1(_04491_),
    .A2(_04492_),
    .B1(_04494_),
    .X(_04593_));
 sky130_fd_sc_hd__xnor2_1 _11437_ (.A(_04592_),
    .B(_04593_),
    .Y(_04594_));
 sky130_fd_sc_hd__mux2_1 _11438_ (.A0(_04077_),
    .A1(_04594_),
    .S(net263),
    .X(_04595_));
 sky130_fd_sc_hd__mux2_1 _11439_ (.A0(net204),
    .A1(_02295_),
    .S(_05796_),
    .X(_04596_));
 sky130_fd_sc_hd__a2bb2o_1 _11440_ (.A1_N(reg1_val[18]),
    .A2_N(_05778_),
    .B1(_02291_),
    .B2(_04596_),
    .X(_04597_));
 sky130_fd_sc_hd__o221a_1 _11441_ (.A1(net184),
    .A2(_04065_),
    .B1(_04078_),
    .B2(net182),
    .C1(_04597_),
    .X(_04598_));
 sky130_fd_sc_hd__or2_1 _11442_ (.A(\div_shifter[49] ),
    .B(_04506_),
    .X(_04599_));
 sky130_fd_sc_hd__a21oi_1 _11443_ (.A1(net244),
    .A2(_04599_),
    .B1(\div_shifter[50] ),
    .Y(_04601_));
 sky130_fd_sc_hd__a31o_1 _11444_ (.A1(\div_shifter[50] ),
    .A2(net244),
    .A3(_04599_),
    .B1(net248),
    .X(_04602_));
 sky130_fd_sc_hd__or2_1 _11445_ (.A(\div_res[17] ),
    .B(_04499_),
    .X(_04603_));
 sky130_fd_sc_hd__and3_1 _11446_ (.A(\div_res[18] ),
    .B(net24),
    .C(_04603_),
    .X(_04604_));
 sky130_fd_sc_hd__a21oi_1 _11447_ (.A1(net25),
    .A2(_04603_),
    .B1(\div_res[18] ),
    .Y(_04605_));
 sky130_fd_sc_hd__or3_1 _11448_ (.A(net202),
    .B(_04604_),
    .C(_04605_),
    .X(_04606_));
 sky130_fd_sc_hd__o21a_1 _11449_ (.A1(_04601_),
    .A2(_04602_),
    .B1(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__nand2_1 _11450_ (.A(_04598_),
    .B(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__a211o_1 _11451_ (.A1(_06412_),
    .A2(_04595_),
    .B1(_04608_),
    .C1(_04588_),
    .X(_04609_));
 sky130_fd_sc_hd__a221o_1 _11452_ (.A1(_04580_),
    .A2(_04581_),
    .B1(_04584_),
    .B2(_02298_),
    .C1(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__a22o_1 _11453_ (.A1(_05778_),
    .A2(net212),
    .B1(_06427_),
    .B2(_04610_),
    .X(_04612_));
 sky130_fd_sc_hd__and2_1 _11454_ (.A(curr_PC[18]),
    .B(_04408_),
    .X(_04613_));
 sky130_fd_sc_hd__o21ai_1 _11455_ (.A1(curr_PC[18]),
    .A2(_04408_),
    .B1(net262),
    .Y(_04614_));
 sky130_fd_sc_hd__a2bb2o_4 _11456_ (.A1_N(_04613_),
    .A2_N(_04614_),
    .B1(net258),
    .B2(_04612_),
    .X(dest_val[18]));
 sky130_fd_sc_hd__o22a_1 _11457_ (.A1(net73),
    .A2(net7),
    .B1(net5),
    .B2(net76),
    .X(_04615_));
 sky130_fd_sc_hd__xnor2_1 _11458_ (.A(net29),
    .B(_04615_),
    .Y(_04616_));
 sky130_fd_sc_hd__and2b_1 _11459_ (.A_N(_04616_),
    .B(_04540_),
    .X(_04617_));
 sky130_fd_sc_hd__and2b_1 _11460_ (.A_N(_04540_),
    .B(_04616_),
    .X(_04618_));
 sky130_fd_sc_hd__or2_1 _11461_ (.A(_04617_),
    .B(_04618_),
    .X(_04619_));
 sky130_fd_sc_hd__nor3_1 _11462_ (.A(net70),
    .B(net30),
    .C(_04619_),
    .Y(_04620_));
 sky130_fd_sc_hd__o21a_1 _11463_ (.A1(net70),
    .A2(net30),
    .B1(_04619_),
    .X(_04622_));
 sky130_fd_sc_hd__nor2_1 _11464_ (.A(_04620_),
    .B(_04622_),
    .Y(_04623_));
 sky130_fd_sc_hd__inv_2 _11465_ (.A(_04623_),
    .Y(_04624_));
 sky130_fd_sc_hd__o22a_1 _11466_ (.A1(net18),
    .A2(net50),
    .B1(net48),
    .B2(net16),
    .X(_04625_));
 sky130_fd_sc_hd__xnor2_1 _11467_ (.A(net105),
    .B(_04625_),
    .Y(_04626_));
 sky130_fd_sc_hd__xnor2_1 _11468_ (.A(_00436_),
    .B(_04626_),
    .Y(_04627_));
 sky130_fd_sc_hd__o22a_1 _11469_ (.A1(net10),
    .A2(net41),
    .B1(net39),
    .B2(net3),
    .X(_04628_));
 sky130_fd_sc_hd__xor2_1 _11470_ (.A(net104),
    .B(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__nor2_1 _11471_ (.A(_04627_),
    .B(_04629_),
    .Y(_04630_));
 sky130_fd_sc_hd__and2_1 _11472_ (.A(_04627_),
    .B(_04629_),
    .X(_04631_));
 sky130_fd_sc_hd__or2_1 _11473_ (.A(_04630_),
    .B(_04631_),
    .X(_04633_));
 sky130_fd_sc_hd__xor2_1 _11474_ (.A(_04623_),
    .B(_04633_),
    .X(_04634_));
 sky130_fd_sc_hd__o22a_1 _11475_ (.A1(net67),
    .A2(net11),
    .B1(net44),
    .B2(net64),
    .X(_04635_));
 sky130_fd_sc_hd__xnor2_1 _11476_ (.A(net96),
    .B(_04635_),
    .Y(_04636_));
 sky130_fd_sc_hd__o22a_1 _11477_ (.A1(net62),
    .A2(net13),
    .B1(net47),
    .B2(net60),
    .X(_04637_));
 sky130_fd_sc_hd__xnor2_1 _11478_ (.A(net108),
    .B(_04637_),
    .Y(_04638_));
 sky130_fd_sc_hd__nand2b_1 _11479_ (.A_N(_04636_),
    .B(_04638_),
    .Y(_04639_));
 sky130_fd_sc_hd__xnor2_1 _11480_ (.A(_04636_),
    .B(_04638_),
    .Y(_04640_));
 sky130_fd_sc_hd__o22a_1 _11481_ (.A1(net57),
    .A2(net14),
    .B1(net52),
    .B2(net54),
    .X(_04641_));
 sky130_fd_sc_hd__xnor2_1 _11482_ (.A(net111),
    .B(_04641_),
    .Y(_04642_));
 sky130_fd_sc_hd__xnor2_1 _11483_ (.A(_04640_),
    .B(_04642_),
    .Y(_04644_));
 sky130_fd_sc_hd__or2_1 _11484_ (.A(_04634_),
    .B(_04644_),
    .X(_04645_));
 sky130_fd_sc_hd__nand2_1 _11485_ (.A(_04634_),
    .B(_04644_),
    .Y(_04646_));
 sky130_fd_sc_hd__and2_1 _11486_ (.A(_04645_),
    .B(_04646_),
    .X(_04647_));
 sky130_fd_sc_hd__o21ai_2 _11487_ (.A1(_04524_),
    .A2(_04548_),
    .B1(_04546_),
    .Y(_04648_));
 sky130_fd_sc_hd__o21ai_1 _11488_ (.A1(_04516_),
    .A2(_04523_),
    .B1(_04521_),
    .Y(_04649_));
 sky130_fd_sc_hd__o31a_1 _11489_ (.A1(net119),
    .A2(net29),
    .A3(_04540_),
    .B1(_04543_),
    .X(_04650_));
 sky130_fd_sc_hd__a21o_1 _11490_ (.A1(_04530_),
    .A2(_04535_),
    .B1(_04650_),
    .X(_04651_));
 sky130_fd_sc_hd__nand3_1 _11491_ (.A(_04530_),
    .B(_04535_),
    .C(_04650_),
    .Y(_04652_));
 sky130_fd_sc_hd__nand2_1 _11492_ (.A(_04651_),
    .B(_04652_),
    .Y(_04653_));
 sky130_fd_sc_hd__nand2b_1 _11493_ (.A_N(_04653_),
    .B(_04649_),
    .Y(_04655_));
 sky130_fd_sc_hd__xor2_1 _11494_ (.A(_04649_),
    .B(_04653_),
    .X(_04656_));
 sky130_fd_sc_hd__a21boi_1 _11495_ (.A1(_04551_),
    .A2(_04555_),
    .B1_N(_04554_),
    .Y(_04657_));
 sky130_fd_sc_hd__or2_1 _11496_ (.A(_04656_),
    .B(_04657_),
    .X(_04658_));
 sky130_fd_sc_hd__xnor2_1 _11497_ (.A(_04656_),
    .B(_04657_),
    .Y(_04659_));
 sky130_fd_sc_hd__nand2b_1 _11498_ (.A_N(_04659_),
    .B(_04648_),
    .Y(_04660_));
 sky130_fd_sc_hd__xnor2_1 _11499_ (.A(_04648_),
    .B(_04659_),
    .Y(_04661_));
 sky130_fd_sc_hd__nand2_1 _11500_ (.A(_04647_),
    .B(_04661_),
    .Y(_04662_));
 sky130_fd_sc_hd__or2_1 _11501_ (.A(_04647_),
    .B(_04661_),
    .X(_04663_));
 sky130_fd_sc_hd__nand2_1 _11502_ (.A(_04662_),
    .B(_04663_),
    .Y(_04664_));
 sky130_fd_sc_hd__a21o_1 _11503_ (.A1(_04557_),
    .A2(_04560_),
    .B1(_04664_),
    .X(_04666_));
 sky130_fd_sc_hd__nand3_1 _11504_ (.A(_04557_),
    .B(_04560_),
    .C(_04664_),
    .Y(_04667_));
 sky130_fd_sc_hd__nand2_1 _11505_ (.A(_04666_),
    .B(_04667_),
    .Y(_04668_));
 sky130_fd_sc_hd__and3_1 _11506_ (.A(_04562_),
    .B(_04565_),
    .C(_04668_),
    .X(_04669_));
 sky130_fd_sc_hd__a21o_1 _11507_ (.A1(_04562_),
    .A2(_04565_),
    .B1(_04668_),
    .X(_04670_));
 sky130_fd_sc_hd__nand2b_1 _11508_ (.A_N(_04669_),
    .B(_04670_),
    .Y(_04671_));
 sky130_fd_sc_hd__or3_1 _11509_ (.A(_04569_),
    .B(_04575_),
    .C(_04671_),
    .X(_04672_));
 sky130_fd_sc_hd__o21ai_1 _11510_ (.A1(_04569_),
    .A2(_04575_),
    .B1(_04671_),
    .Y(_04673_));
 sky130_fd_sc_hd__nand2_1 _11511_ (.A(_04672_),
    .B(_04673_),
    .Y(_04674_));
 sky130_fd_sc_hd__o2111a_1 _11512_ (.A1(_04575_),
    .A2(_04576_),
    .B1(_04369_),
    .C1(_04478_),
    .D1(_04479_),
    .X(_04675_));
 sky130_fd_sc_hd__nand2_1 _11513_ (.A(_04371_),
    .B(_04675_),
    .Y(_04677_));
 sky130_fd_sc_hd__nand3_1 _11514_ (.A(net27),
    .B(_04674_),
    .C(_04677_),
    .Y(_04678_));
 sky130_fd_sc_hd__a21o_1 _11515_ (.A1(net27),
    .A2(_04677_),
    .B1(_04674_),
    .X(_04679_));
 sky130_fd_sc_hd__a21oi_1 _11516_ (.A1(net20),
    .A2(_02192_),
    .B1(_02194_),
    .Y(_04680_));
 sky130_fd_sc_hd__a31o_1 _11517_ (.A1(net20),
    .A2(_02192_),
    .A3(_02194_),
    .B1(_02299_),
    .X(_04681_));
 sky130_fd_sc_hd__a21bo_1 _11518_ (.A1(_05814_),
    .A2(_04585_),
    .B1_N(_05796_),
    .X(_04682_));
 sky130_fd_sc_hd__and2_1 _11519_ (.A(net299),
    .B(_04682_),
    .X(_04683_));
 sky130_fd_sc_hd__a31o_1 _11520_ (.A1(net305),
    .A2(_05787_),
    .A3(_06332_),
    .B1(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__nand2_1 _11521_ (.A(_05741_),
    .B(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__o211a_1 _11522_ (.A1(_05741_),
    .A2(_04684_),
    .B1(_04685_),
    .C1(net251),
    .X(_04686_));
 sky130_fd_sc_hd__nor2_1 _11523_ (.A(reg1_val[19]),
    .B(curr_PC[19]),
    .Y(_04688_));
 sky130_fd_sc_hd__nand2_1 _11524_ (.A(reg1_val[19]),
    .B(curr_PC[19]),
    .Y(_04689_));
 sky130_fd_sc_hd__and2b_1 _11525_ (.A_N(_04688_),
    .B(_04689_),
    .X(_04690_));
 sky130_fd_sc_hd__o21a_1 _11526_ (.A1(_04590_),
    .A2(_04593_),
    .B1(_04591_),
    .X(_04691_));
 sky130_fd_sc_hd__xnor2_1 _11527_ (.A(_04690_),
    .B(_04691_),
    .Y(_04692_));
 sky130_fd_sc_hd__mux2_1 _11528_ (.A0(_03968_),
    .A1(_04692_),
    .S(net263),
    .X(_04693_));
 sky130_fd_sc_hd__or2_1 _11529_ (.A(\div_res[18] ),
    .B(_04603_),
    .X(_04694_));
 sky130_fd_sc_hd__a21oi_1 _11530_ (.A1(net24),
    .A2(_04694_),
    .B1(\div_res[19] ),
    .Y(_04695_));
 sky130_fd_sc_hd__a311o_1 _11531_ (.A1(\div_res[19] ),
    .A2(net24),
    .A3(_04694_),
    .B1(_04695_),
    .C1(net202),
    .X(_04696_));
 sky130_fd_sc_hd__or2_1 _11532_ (.A(\div_shifter[50] ),
    .B(_04599_),
    .X(_04697_));
 sky130_fd_sc_hd__a21oi_1 _11533_ (.A1(net244),
    .A2(_04697_),
    .B1(\div_shifter[51] ),
    .Y(_04699_));
 sky130_fd_sc_hd__a31o_1 _11534_ (.A1(\div_shifter[51] ),
    .A2(net244),
    .A3(_04697_),
    .B1(net248),
    .X(_04700_));
 sky130_fd_sc_hd__nor2_1 _11535_ (.A(_05723_),
    .B(net204),
    .Y(_04701_));
 sky130_fd_sc_hd__a211o_1 _11536_ (.A1(_05723_),
    .A2(_02294_),
    .B1(_04701_),
    .C1(net205),
    .X(_04702_));
 sky130_fd_sc_hd__o2bb2a_1 _11537_ (.A1_N(_05732_),
    .A2_N(_04702_),
    .B1(_03969_),
    .B2(net182),
    .X(_04703_));
 sky130_fd_sc_hd__o211a_1 _11538_ (.A1(net186),
    .A2(_03951_),
    .B1(_04696_),
    .C1(_04703_),
    .X(_04704_));
 sky130_fd_sc_hd__o21ai_2 _11539_ (.A1(_04699_),
    .A2(_04700_),
    .B1(_04704_),
    .Y(_04705_));
 sky130_fd_sc_hd__a211oi_2 _11540_ (.A1(_06412_),
    .A2(_04693_),
    .B1(_04705_),
    .C1(_04686_),
    .Y(_04706_));
 sky130_fd_sc_hd__o21ai_1 _11541_ (.A1(_04680_),
    .A2(_04681_),
    .B1(_04706_),
    .Y(_04707_));
 sky130_fd_sc_hd__a31o_1 _11542_ (.A1(net206),
    .A2(_04678_),
    .A3(_04679_),
    .B1(_04707_),
    .X(_04708_));
 sky130_fd_sc_hd__a22o_1 _11543_ (.A1(_05696_),
    .A2(net212),
    .B1(_06427_),
    .B2(_04708_),
    .X(_04710_));
 sky130_fd_sc_hd__or2_1 _11544_ (.A(curr_PC[19]),
    .B(_04613_),
    .X(_04711_));
 sky130_fd_sc_hd__a21oi_1 _11545_ (.A1(curr_PC[19]),
    .A2(_04613_),
    .B1(net258),
    .Y(_04712_));
 sky130_fd_sc_hd__a22o_4 _11546_ (.A1(net258),
    .A2(_04710_),
    .B1(_04711_),
    .B2(_04712_),
    .X(dest_val[19]));
 sky130_fd_sc_hd__or2_1 _11547_ (.A(_04571_),
    .B(_04671_),
    .X(_04713_));
 sky130_fd_sc_hd__a211o_1 _11548_ (.A1(_04299_),
    .A2(_04300_),
    .B1(_04573_),
    .C1(_04713_),
    .X(_04714_));
 sky130_fd_sc_hd__o221a_1 _11549_ (.A1(_04570_),
    .A2(_04669_),
    .B1(_04713_),
    .B2(_04572_),
    .C1(_04670_),
    .X(_04715_));
 sky130_fd_sc_hd__o22a_1 _11550_ (.A1(net64),
    .A2(net11),
    .B1(net44),
    .B2(net57),
    .X(_04716_));
 sky130_fd_sc_hd__xnor2_1 _11551_ (.A(net96),
    .B(_04716_),
    .Y(_04717_));
 sky130_fd_sc_hd__a22o_1 _11552_ (.A1(_00197_),
    .A2(_00307_),
    .B1(_00308_),
    .B2(_00222_),
    .X(_04718_));
 sky130_fd_sc_hd__xor2_1 _11553_ (.A(net108),
    .B(_04718_),
    .X(_04720_));
 sky130_fd_sc_hd__nand2b_1 _11554_ (.A_N(_04717_),
    .B(_04720_),
    .Y(_04721_));
 sky130_fd_sc_hd__nand2b_1 _11555_ (.A_N(_04720_),
    .B(_04717_),
    .Y(_04722_));
 sky130_fd_sc_hd__nand2_1 _11556_ (.A(_04721_),
    .B(_04722_),
    .Y(_04723_));
 sky130_fd_sc_hd__o22a_1 _11557_ (.A1(net54),
    .A2(net14),
    .B1(net52),
    .B2(net62),
    .X(_04724_));
 sky130_fd_sc_hd__xnor2_1 _11558_ (.A(net111),
    .B(_04724_),
    .Y(_04725_));
 sky130_fd_sc_hd__nand2b_1 _11559_ (.A_N(_04723_),
    .B(_04725_),
    .Y(_04726_));
 sky130_fd_sc_hd__nand2b_1 _11560_ (.A_N(_04725_),
    .B(_04723_),
    .Y(_04727_));
 sky130_fd_sc_hd__nand2_1 _11561_ (.A(_04726_),
    .B(_04727_),
    .Y(_04728_));
 sky130_fd_sc_hd__o22a_1 _11562_ (.A1(net17),
    .A2(net50),
    .B1(net48),
    .B2(_00408_),
    .X(_04729_));
 sky130_fd_sc_hd__xnor2_1 _11563_ (.A(net105),
    .B(_04729_),
    .Y(_04731_));
 sky130_fd_sc_hd__nor2_1 _11564_ (.A(net40),
    .B(net3),
    .Y(_04732_));
 sky130_fd_sc_hd__xnor2_1 _11565_ (.A(net102),
    .B(_04732_),
    .Y(_04733_));
 sky130_fd_sc_hd__and2b_1 _11566_ (.A_N(_04731_),
    .B(_04733_),
    .X(_04734_));
 sky130_fd_sc_hd__and2b_1 _11567_ (.A_N(_04733_),
    .B(_04731_),
    .X(_04735_));
 sky130_fd_sc_hd__or2_1 _11568_ (.A(_04734_),
    .B(_04735_),
    .X(_04736_));
 sky130_fd_sc_hd__o22a_1 _11569_ (.A1(net67),
    .A2(net7),
    .B1(net5),
    .B2(net73),
    .X(_04737_));
 sky130_fd_sc_hd__nor2_1 _11570_ (.A(_06503_),
    .B(net30),
    .Y(_04738_));
 sky130_fd_sc_hd__xnor2_1 _11571_ (.A(_04737_),
    .B(_04738_),
    .Y(_04739_));
 sky130_fd_sc_hd__nand2_1 _11572_ (.A(_04736_),
    .B(_04739_),
    .Y(_04740_));
 sky130_fd_sc_hd__xnor2_1 _11573_ (.A(_04736_),
    .B(_04739_),
    .Y(_04742_));
 sky130_fd_sc_hd__xor2_1 _11574_ (.A(_04728_),
    .B(_04742_),
    .X(_04743_));
 sky130_fd_sc_hd__o21a_1 _11575_ (.A1(_04624_),
    .A2(_04633_),
    .B1(_04645_),
    .X(_04744_));
 sky130_fd_sc_hd__a21bo_1 _11576_ (.A1(_04640_),
    .A2(_04642_),
    .B1_N(_04639_),
    .X(_04745_));
 sky130_fd_sc_hd__a21oi_1 _11577_ (.A1(_00436_),
    .A2(_04626_),
    .B1(_04630_),
    .Y(_04746_));
 sky130_fd_sc_hd__o21ba_1 _11578_ (.A1(_04617_),
    .A2(_04620_),
    .B1_N(_04746_),
    .X(_04747_));
 sky130_fd_sc_hd__or3b_1 _11579_ (.A(_04617_),
    .B(_04620_),
    .C_N(_04746_),
    .X(_04748_));
 sky130_fd_sc_hd__and2b_1 _11580_ (.A_N(_04747_),
    .B(_04748_),
    .X(_04749_));
 sky130_fd_sc_hd__and2_1 _11581_ (.A(_04745_),
    .B(_04749_),
    .X(_04750_));
 sky130_fd_sc_hd__or2_1 _11582_ (.A(_04745_),
    .B(_04749_),
    .X(_04751_));
 sky130_fd_sc_hd__nand2b_1 _11583_ (.A_N(_04750_),
    .B(_04751_),
    .Y(_04753_));
 sky130_fd_sc_hd__a21oi_1 _11584_ (.A1(_04651_),
    .A2(_04655_),
    .B1(_04753_),
    .Y(_04754_));
 sky130_fd_sc_hd__and3_1 _11585_ (.A(_04651_),
    .B(_04655_),
    .C(_04753_),
    .X(_04755_));
 sky130_fd_sc_hd__nor2_1 _11586_ (.A(_04754_),
    .B(_04755_),
    .Y(_04756_));
 sky130_fd_sc_hd__and2b_1 _11587_ (.A_N(_04744_),
    .B(_04756_),
    .X(_04757_));
 sky130_fd_sc_hd__xnor2_1 _11588_ (.A(_04744_),
    .B(_04756_),
    .Y(_04758_));
 sky130_fd_sc_hd__and2_1 _11589_ (.A(_04743_),
    .B(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__nor2_1 _11590_ (.A(_04743_),
    .B(_04758_),
    .Y(_04760_));
 sky130_fd_sc_hd__or2_1 _11591_ (.A(_04759_),
    .B(_04760_),
    .X(_04761_));
 sky130_fd_sc_hd__a21oi_1 _11592_ (.A1(_04658_),
    .A2(_04660_),
    .B1(_04761_),
    .Y(_04762_));
 sky130_fd_sc_hd__and3_1 _11593_ (.A(_04658_),
    .B(_04660_),
    .C(_04761_),
    .X(_04764_));
 sky130_fd_sc_hd__or2_1 _11594_ (.A(_04762_),
    .B(_04764_),
    .X(_04765_));
 sky130_fd_sc_hd__a21oi_1 _11595_ (.A1(_04662_),
    .A2(_04666_),
    .B1(_04765_),
    .Y(_04766_));
 sky130_fd_sc_hd__and3_1 _11596_ (.A(_04662_),
    .B(_04666_),
    .C(_04765_),
    .X(_04767_));
 sky130_fd_sc_hd__or2_1 _11597_ (.A(_04766_),
    .B(_04767_),
    .X(_04768_));
 sky130_fd_sc_hd__a21oi_1 _11598_ (.A1(_04714_),
    .A2(_04715_),
    .B1(_04768_),
    .Y(_04769_));
 sky130_fd_sc_hd__a21o_1 _11599_ (.A1(_04714_),
    .A2(_04715_),
    .B1(_04768_),
    .X(_04770_));
 sky130_fd_sc_hd__and3_1 _11600_ (.A(_04714_),
    .B(_04715_),
    .C(_04768_),
    .X(_04771_));
 sky130_fd_sc_hd__nor2_1 _11601_ (.A(_04769_),
    .B(_04771_),
    .Y(_04772_));
 sky130_fd_sc_hd__inv_2 _11602_ (.A(_04772_),
    .Y(_04773_));
 sky130_fd_sc_hd__and3_1 _11603_ (.A(_04672_),
    .B(_04673_),
    .C(_04675_),
    .X(_04775_));
 sky130_fd_sc_hd__a21o_1 _11604_ (.A1(_04371_),
    .A2(_04775_),
    .B1(net84),
    .X(_04776_));
 sky130_fd_sc_hd__o21ai_1 _11605_ (.A1(_04773_),
    .A2(_04776_),
    .B1(net206),
    .Y(_04777_));
 sky130_fd_sc_hd__a21oi_1 _11606_ (.A1(_04773_),
    .A2(_04776_),
    .B1(_04777_),
    .Y(_04778_));
 sky130_fd_sc_hd__a21o_1 _11607_ (.A1(net20),
    .A2(_02195_),
    .B1(_02196_),
    .X(_04779_));
 sky130_fd_sc_hd__nand3_1 _11608_ (.A(net20),
    .B(_02195_),
    .C(_02196_),
    .Y(_04780_));
 sky130_fd_sc_hd__a21bo_1 _11609_ (.A1(_05741_),
    .A2(_04682_),
    .B1_N(_05723_),
    .X(_04781_));
 sky130_fd_sc_hd__mux2_1 _11610_ (.A0(_06334_),
    .A1(_04781_),
    .S(net299),
    .X(_04782_));
 sky130_fd_sc_hd__o21ai_1 _11611_ (.A1(_05668_),
    .A2(_04782_),
    .B1(net251),
    .Y(_04783_));
 sky130_fd_sc_hd__a21o_1 _11612_ (.A1(_05668_),
    .A2(_04782_),
    .B1(_04783_),
    .X(_04784_));
 sky130_fd_sc_hd__or2_1 _11613_ (.A(reg1_val[20]),
    .B(curr_PC[20]),
    .X(_04786_));
 sky130_fd_sc_hd__nand2_1 _11614_ (.A(reg1_val[20]),
    .B(curr_PC[20]),
    .Y(_04787_));
 sky130_fd_sc_hd__nand2_1 _11615_ (.A(_04786_),
    .B(_04787_),
    .Y(_04788_));
 sky130_fd_sc_hd__o21a_1 _11616_ (.A1(_04688_),
    .A2(_04691_),
    .B1(_04689_),
    .X(_04789_));
 sky130_fd_sc_hd__xnor2_1 _11617_ (.A(_04788_),
    .B(_04789_),
    .Y(_04790_));
 sky130_fd_sc_hd__mux2_1 _11618_ (.A0(_03855_),
    .A1(_04790_),
    .S(net263),
    .X(_04791_));
 sky130_fd_sc_hd__or2_1 _11619_ (.A(\div_res[19] ),
    .B(_04694_),
    .X(_04792_));
 sky130_fd_sc_hd__and3_1 _11620_ (.A(\div_res[20] ),
    .B(net24),
    .C(_04792_),
    .X(_04793_));
 sky130_fd_sc_hd__a21oi_1 _11621_ (.A1(net23),
    .A2(_04792_),
    .B1(\div_res[20] ),
    .Y(_04794_));
 sky130_fd_sc_hd__or2_1 _11622_ (.A(\div_shifter[51] ),
    .B(_04697_),
    .X(_04795_));
 sky130_fd_sc_hd__and3_1 _11623_ (.A(\div_shifter[52] ),
    .B(net244),
    .C(_04795_),
    .X(_04797_));
 sky130_fd_sc_hd__a21oi_1 _11624_ (.A1(net244),
    .A2(_04795_),
    .B1(\div_shifter[52] ),
    .Y(_04798_));
 sky130_fd_sc_hd__or2_1 _11625_ (.A(_05639_),
    .B(net204),
    .X(_04799_));
 sky130_fd_sc_hd__o211a_1 _11626_ (.A1(_05649_),
    .A2(_02295_),
    .B1(_04799_),
    .C1(_02291_),
    .X(_04800_));
 sky130_fd_sc_hd__o22a_1 _11627_ (.A1(_05611_),
    .A2(_06426_),
    .B1(_04800_),
    .B2(_05658_),
    .X(_04801_));
 sky130_fd_sc_hd__o221a_1 _11628_ (.A1(net186),
    .A2(_03842_),
    .B1(_03855_),
    .B2(net182),
    .C1(_04801_),
    .X(_04802_));
 sky130_fd_sc_hd__o31a_1 _11629_ (.A1(net248),
    .A2(_04797_),
    .A3(_04798_),
    .B1(_04802_),
    .X(_04803_));
 sky130_fd_sc_hd__o31a_1 _11630_ (.A1(net202),
    .A2(_04793_),
    .A3(_04794_),
    .B1(_04803_),
    .X(_04804_));
 sky130_fd_sc_hd__o211ai_2 _11631_ (.A1(net214),
    .A2(_04791_),
    .B1(_04804_),
    .C1(_04784_),
    .Y(_04805_));
 sky130_fd_sc_hd__a311o_1 _11632_ (.A1(_02298_),
    .A2(_04779_),
    .A3(_04780_),
    .B1(_04805_),
    .C1(_04778_),
    .X(_04806_));
 sky130_fd_sc_hd__and3_1 _11633_ (.A(curr_PC[19]),
    .B(curr_PC[20]),
    .C(_04613_),
    .X(_04808_));
 sky130_fd_sc_hd__a21oi_1 _11634_ (.A1(curr_PC[19]),
    .A2(_04613_),
    .B1(curr_PC[20]),
    .Y(_04809_));
 sky130_fd_sc_hd__nor2_1 _11635_ (.A(_04808_),
    .B(_04809_),
    .Y(_04810_));
 sky130_fd_sc_hd__mux2_8 _11636_ (.A0(_04806_),
    .A1(_04810_),
    .S(net262),
    .X(dest_val[20]));
 sky130_fd_sc_hd__o22a_1 _11637_ (.A1(net57),
    .A2(net12),
    .B1(net44),
    .B2(net55),
    .X(_04811_));
 sky130_fd_sc_hd__xnor2_1 _11638_ (.A(net96),
    .B(_04811_),
    .Y(_04812_));
 sky130_fd_sc_hd__o22a_1 _11639_ (.A1(net65),
    .A2(net8),
    .B1(net6),
    .B2(net68),
    .X(_04813_));
 sky130_fd_sc_hd__xnor2_1 _11640_ (.A(net31),
    .B(_04813_),
    .Y(_04814_));
 sky130_fd_sc_hd__o22a_1 _11641_ (.A1(net63),
    .A2(net15),
    .B1(net53),
    .B2(net60),
    .X(_04815_));
 sky130_fd_sc_hd__xnor2_1 _11642_ (.A(net111),
    .B(_04815_),
    .Y(_04816_));
 sky130_fd_sc_hd__nand2b_1 _11643_ (.A_N(_04814_),
    .B(_04816_),
    .Y(_04818_));
 sky130_fd_sc_hd__nand2b_1 _11644_ (.A_N(_04816_),
    .B(_04814_),
    .Y(_04819_));
 sky130_fd_sc_hd__nand2_1 _11645_ (.A(_04818_),
    .B(_04819_),
    .Y(_04820_));
 sky130_fd_sc_hd__or2_1 _11646_ (.A(_04812_),
    .B(_04820_),
    .X(_04821_));
 sky130_fd_sc_hd__nand2_1 _11647_ (.A(_04812_),
    .B(_04820_),
    .Y(_04822_));
 sky130_fd_sc_hd__and2_1 _11648_ (.A(_04821_),
    .B(_04822_),
    .X(_04823_));
 sky130_fd_sc_hd__and3_1 _11649_ (.A(_06503_),
    .B(net33),
    .C(_04737_),
    .X(_04824_));
 sky130_fd_sc_hd__xnor2_1 _11650_ (.A(_04823_),
    .B(_04824_),
    .Y(_04825_));
 sky130_fd_sc_hd__a22o_1 _11651_ (.A1(_00222_),
    .A2(_00307_),
    .B1(_00308_),
    .B2(_00228_),
    .X(_04826_));
 sky130_fd_sc_hd__xor2_1 _11652_ (.A(_00255_),
    .B(_04826_),
    .X(_04827_));
 sky130_fd_sc_hd__and2b_1 _11653_ (.A_N(net102),
    .B(_04827_),
    .X(_04829_));
 sky130_fd_sc_hd__xnor2_1 _11654_ (.A(net102),
    .B(_04827_),
    .Y(_04830_));
 sky130_fd_sc_hd__o22a_1 _11655_ (.A1(net51),
    .A2(net10),
    .B1(net3),
    .B2(_00291_),
    .X(_04831_));
 sky130_fd_sc_hd__xnor2_1 _11656_ (.A(net105),
    .B(_04831_),
    .Y(_04832_));
 sky130_fd_sc_hd__xnor2_1 _11657_ (.A(_04830_),
    .B(_04832_),
    .Y(_04833_));
 sky130_fd_sc_hd__or2_1 _11658_ (.A(_04825_),
    .B(_04833_),
    .X(_04834_));
 sky130_fd_sc_hd__nand2_1 _11659_ (.A(_04825_),
    .B(_04833_),
    .Y(_04835_));
 sky130_fd_sc_hd__nand2_1 _11660_ (.A(_04834_),
    .B(_04835_),
    .Y(_04836_));
 sky130_fd_sc_hd__o21a_1 _11661_ (.A1(_04728_),
    .A2(_04742_),
    .B1(_04740_),
    .X(_04837_));
 sky130_fd_sc_hd__nand2_1 _11662_ (.A(_04721_),
    .B(_04726_),
    .Y(_04838_));
 sky130_fd_sc_hd__nor2_1 _11663_ (.A(net73),
    .B(net30),
    .Y(_04840_));
 sky130_fd_sc_hd__nand2_1 _11664_ (.A(_04838_),
    .B(_04840_),
    .Y(_04841_));
 sky130_fd_sc_hd__xnor2_1 _11665_ (.A(_04838_),
    .B(_04840_),
    .Y(_04842_));
 sky130_fd_sc_hd__xor2_1 _11666_ (.A(_04734_),
    .B(_04842_),
    .X(_04843_));
 sky130_fd_sc_hd__o21ai_1 _11667_ (.A1(_04747_),
    .A2(_04750_),
    .B1(_04843_),
    .Y(_04844_));
 sky130_fd_sc_hd__or3_1 _11668_ (.A(_04747_),
    .B(_04750_),
    .C(_04843_),
    .X(_04845_));
 sky130_fd_sc_hd__and2_1 _11669_ (.A(_04844_),
    .B(_04845_),
    .X(_04846_));
 sky130_fd_sc_hd__nand2b_1 _11670_ (.A_N(_04837_),
    .B(_04846_),
    .Y(_04847_));
 sky130_fd_sc_hd__xnor2_1 _11671_ (.A(_04837_),
    .B(_04846_),
    .Y(_04848_));
 sky130_fd_sc_hd__xnor2_1 _11672_ (.A(_04836_),
    .B(_04848_),
    .Y(_04849_));
 sky130_fd_sc_hd__o21a_1 _11673_ (.A1(_04754_),
    .A2(_04757_),
    .B1(_04849_),
    .X(_04851_));
 sky130_fd_sc_hd__nor3_1 _11674_ (.A(_04754_),
    .B(_04757_),
    .C(_04849_),
    .Y(_04852_));
 sky130_fd_sc_hd__nor2_1 _11675_ (.A(_04851_),
    .B(_04852_),
    .Y(_04853_));
 sky130_fd_sc_hd__o21a_1 _11676_ (.A1(_04759_),
    .A2(_04762_),
    .B1(_04853_),
    .X(_04854_));
 sky130_fd_sc_hd__nor3_1 _11677_ (.A(_04759_),
    .B(_04762_),
    .C(_04853_),
    .Y(_04855_));
 sky130_fd_sc_hd__or2_2 _11678_ (.A(_04854_),
    .B(_04855_),
    .X(_04856_));
 sky130_fd_sc_hd__nor2_1 _11679_ (.A(_04766_),
    .B(_04769_),
    .Y(_04857_));
 sky130_fd_sc_hd__xnor2_1 _11680_ (.A(_04856_),
    .B(_04857_),
    .Y(_04858_));
 sky130_fd_sc_hd__xor2_1 _11681_ (.A(_04856_),
    .B(_04857_),
    .X(_04859_));
 sky130_fd_sc_hd__a31oi_1 _11682_ (.A1(_04371_),
    .A2(_04773_),
    .A3(_04775_),
    .B1(net86),
    .Y(_04860_));
 sky130_fd_sc_hd__nand2_1 _11683_ (.A(_04859_),
    .B(_04860_),
    .Y(_04862_));
 sky130_fd_sc_hd__o21a_1 _11684_ (.A1(_04859_),
    .A2(_04860_),
    .B1(_02213_),
    .X(_04863_));
 sky130_fd_sc_hd__a21o_1 _11685_ (.A1(net20),
    .A2(_02197_),
    .B1(_02151_),
    .X(_04864_));
 sky130_fd_sc_hd__a31oi_1 _11686_ (.A1(net20),
    .A2(_02151_),
    .A3(_02197_),
    .B1(net250),
    .Y(_04865_));
 sky130_fd_sc_hd__a21o_1 _11687_ (.A1(_05668_),
    .A2(_04781_),
    .B1(_05649_),
    .X(_04866_));
 sky130_fd_sc_hd__mux2_1 _11688_ (.A0(_06336_),
    .A1(_04866_),
    .S(net299),
    .X(_04867_));
 sky130_fd_sc_hd__nand2_1 _11689_ (.A(_05582_),
    .B(_04867_),
    .Y(_04868_));
 sky130_fd_sc_hd__o211a_1 _11690_ (.A1(_05582_),
    .A2(_04867_),
    .B1(_04868_),
    .C1(net251),
    .X(_04869_));
 sky130_fd_sc_hd__nor2_1 _11691_ (.A(reg1_val[21]),
    .B(curr_PC[21]),
    .Y(_04870_));
 sky130_fd_sc_hd__nand2_1 _11692_ (.A(reg1_val[21]),
    .B(curr_PC[21]),
    .Y(_04871_));
 sky130_fd_sc_hd__and2b_1 _11693_ (.A_N(_04870_),
    .B(_04871_),
    .X(_04873_));
 sky130_fd_sc_hd__o21a_1 _11694_ (.A1(_04788_),
    .A2(_04789_),
    .B1(_04787_),
    .X(_04874_));
 sky130_fd_sc_hd__xnor2_1 _11695_ (.A(_04873_),
    .B(_04874_),
    .Y(_04875_));
 sky130_fd_sc_hd__nand2_1 _11696_ (.A(net241),
    .B(_03736_),
    .Y(_04876_));
 sky130_fd_sc_hd__o211a_1 _11697_ (.A1(net241),
    .A2(_04875_),
    .B1(_04876_),
    .C1(net215),
    .X(_04877_));
 sky130_fd_sc_hd__or2_1 _11698_ (.A(\div_shifter[52] ),
    .B(_04795_),
    .X(_04878_));
 sky130_fd_sc_hd__a21oi_1 _11699_ (.A1(net244),
    .A2(_04878_),
    .B1(\div_shifter[53] ),
    .Y(_04879_));
 sky130_fd_sc_hd__a311o_1 _11700_ (.A1(\div_shifter[53] ),
    .A2(net244),
    .A3(_04878_),
    .B1(_04879_),
    .C1(net248),
    .X(_04880_));
 sky130_fd_sc_hd__or2_1 _11701_ (.A(\div_res[20] ),
    .B(_04792_),
    .X(_04881_));
 sky130_fd_sc_hd__a21oi_1 _11702_ (.A1(net23),
    .A2(_04881_),
    .B1(\div_res[21] ),
    .Y(_04882_));
 sky130_fd_sc_hd__a31o_1 _11703_ (.A1(\div_res[21] ),
    .A2(net23),
    .A3(_04881_),
    .B1(net202),
    .X(_04884_));
 sky130_fd_sc_hd__mux2_1 _11704_ (.A0(_02295_),
    .A1(net204),
    .S(_05563_),
    .X(_04885_));
 sky130_fd_sc_hd__a21o_1 _11705_ (.A1(_02291_),
    .A2(_04885_),
    .B1(_05572_),
    .X(_04886_));
 sky130_fd_sc_hd__o221a_1 _11706_ (.A1(net185),
    .A2(_03724_),
    .B1(_03736_),
    .B2(net182),
    .C1(_04886_),
    .X(_04887_));
 sky130_fd_sc_hd__o21ai_1 _11707_ (.A1(_04882_),
    .A2(_04884_),
    .B1(_04887_),
    .Y(_04888_));
 sky130_fd_sc_hd__or4b_2 _11708_ (.A(_04869_),
    .B(_04877_),
    .C(_04888_),
    .D_N(_04880_),
    .X(_04889_));
 sky130_fd_sc_hd__a221o_1 _11709_ (.A1(_04862_),
    .A2(_04863_),
    .B1(_04864_),
    .B2(_04865_),
    .C1(_04889_),
    .X(_04890_));
 sky130_fd_sc_hd__a22o_1 _11710_ (.A1(_05544_),
    .A2(net212),
    .B1(_06427_),
    .B2(_04890_),
    .X(_04891_));
 sky130_fd_sc_hd__or2_1 _11711_ (.A(curr_PC[21]),
    .B(_04808_),
    .X(_04892_));
 sky130_fd_sc_hd__and2_1 _11712_ (.A(curr_PC[21]),
    .B(_04808_),
    .X(_04893_));
 sky130_fd_sc_hd__nor2_1 _11713_ (.A(net258),
    .B(_04893_),
    .Y(_04895_));
 sky130_fd_sc_hd__a22o_4 _11714_ (.A1(net257),
    .A2(_04891_),
    .B1(_04892_),
    .B2(_04895_),
    .X(dest_val[21]));
 sky130_fd_sc_hd__o22a_1 _11715_ (.A1(net55),
    .A2(net12),
    .B1(net45),
    .B2(net63),
    .X(_04896_));
 sky130_fd_sc_hd__xnor2_1 _11716_ (.A(net97),
    .B(_04896_),
    .Y(_04897_));
 sky130_fd_sc_hd__o22a_1 _11717_ (.A1(net61),
    .A2(net15),
    .B1(net53),
    .B2(_00223_),
    .X(_04898_));
 sky130_fd_sc_hd__xnor2_1 _11718_ (.A(net111),
    .B(_04898_),
    .Y(_04899_));
 sky130_fd_sc_hd__nand2b_1 _11719_ (.A_N(_04897_),
    .B(_04899_),
    .Y(_04900_));
 sky130_fd_sc_hd__nand2b_1 _11720_ (.A_N(_04899_),
    .B(_04897_),
    .Y(_04901_));
 sky130_fd_sc_hd__nand2_1 _11721_ (.A(_04900_),
    .B(_04901_),
    .Y(_04902_));
 sky130_fd_sc_hd__a21o_1 _11722_ (.A1(_04818_),
    .A2(_04821_),
    .B1(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__nand3_1 _11723_ (.A(_04818_),
    .B(_04821_),
    .C(_04902_),
    .Y(_04905_));
 sky130_fd_sc_hd__nand2_1 _11724_ (.A(_04903_),
    .B(_04905_),
    .Y(_04906_));
 sky130_fd_sc_hd__o22a_1 _11725_ (.A1(net17),
    .A2(net13),
    .B1(_00309_),
    .B2(net10),
    .X(_04907_));
 sky130_fd_sc_hd__xnor2_1 _11726_ (.A(net109),
    .B(_04907_),
    .Y(_04908_));
 sky130_fd_sc_hd__or2_1 _11727_ (.A(_00287_),
    .B(net3),
    .X(_04909_));
 sky130_fd_sc_hd__a22o_1 _11728_ (.A1(_00286_),
    .A2(_00756_),
    .B1(_04909_),
    .B2(net106),
    .X(_04910_));
 sky130_fd_sc_hd__or2_1 _11729_ (.A(_04908_),
    .B(_04910_),
    .X(_04911_));
 sky130_fd_sc_hd__nand2_1 _11730_ (.A(_04908_),
    .B(_04910_),
    .Y(_04912_));
 sky130_fd_sc_hd__and2_1 _11731_ (.A(_04911_),
    .B(_04912_),
    .X(_04913_));
 sky130_fd_sc_hd__xor2_1 _11732_ (.A(_04906_),
    .B(_04913_),
    .X(_04914_));
 sky130_fd_sc_hd__a21bo_1 _11733_ (.A1(_04823_),
    .A2(_04824_),
    .B1_N(_04834_),
    .X(_04916_));
 sky130_fd_sc_hd__a21o_1 _11734_ (.A1(_04830_),
    .A2(_04832_),
    .B1(_04829_),
    .X(_04917_));
 sky130_fd_sc_hd__o22a_1 _11735_ (.A1(net57),
    .A2(net7),
    .B1(net5),
    .B2(net64),
    .X(_04918_));
 sky130_fd_sc_hd__xnor2_1 _11736_ (.A(net30),
    .B(_04918_),
    .Y(_04919_));
 sky130_fd_sc_hd__and2b_1 _11737_ (.A_N(_04919_),
    .B(_04917_),
    .X(_04920_));
 sky130_fd_sc_hd__xnor2_1 _11738_ (.A(_04917_),
    .B(_04919_),
    .Y(_04921_));
 sky130_fd_sc_hd__nor2_1 _11739_ (.A(net67),
    .B(net30),
    .Y(_04922_));
 sky130_fd_sc_hd__and2_1 _11740_ (.A(_04921_),
    .B(_04922_),
    .X(_04923_));
 sky130_fd_sc_hd__xnor2_1 _11741_ (.A(_04921_),
    .B(_04922_),
    .Y(_04924_));
 sky130_fd_sc_hd__o21a_1 _11742_ (.A1(_04734_),
    .A2(_04842_),
    .B1(_04841_),
    .X(_04925_));
 sky130_fd_sc_hd__xnor2_1 _11743_ (.A(_04924_),
    .B(_04925_),
    .Y(_04927_));
 sky130_fd_sc_hd__nand2b_1 _11744_ (.A_N(_04927_),
    .B(_04916_),
    .Y(_04928_));
 sky130_fd_sc_hd__xnor2_1 _11745_ (.A(_04916_),
    .B(_04927_),
    .Y(_04929_));
 sky130_fd_sc_hd__nand2_1 _11746_ (.A(_04914_),
    .B(_04929_),
    .Y(_04930_));
 sky130_fd_sc_hd__or2_1 _11747_ (.A(_04914_),
    .B(_04929_),
    .X(_04931_));
 sky130_fd_sc_hd__nand2_1 _11748_ (.A(_04930_),
    .B(_04931_),
    .Y(_04932_));
 sky130_fd_sc_hd__and2_1 _11749_ (.A(_04844_),
    .B(_04847_),
    .X(_04933_));
 sky130_fd_sc_hd__or2_1 _11750_ (.A(_04932_),
    .B(_04933_),
    .X(_04934_));
 sky130_fd_sc_hd__nand2_1 _11751_ (.A(_04932_),
    .B(_04933_),
    .Y(_04935_));
 sky130_fd_sc_hd__nand2_1 _11752_ (.A(_04934_),
    .B(_04935_),
    .Y(_04936_));
 sky130_fd_sc_hd__a31oi_1 _11753_ (.A1(_04834_),
    .A2(_04835_),
    .A3(_04848_),
    .B1(_04851_),
    .Y(_04938_));
 sky130_fd_sc_hd__nor2_1 _11754_ (.A(_04936_),
    .B(_04938_),
    .Y(_04939_));
 sky130_fd_sc_hd__and2_1 _11755_ (.A(_04936_),
    .B(_04938_),
    .X(_04940_));
 sky130_fd_sc_hd__nor2_2 _11756_ (.A(_04939_),
    .B(_04940_),
    .Y(_04941_));
 sky130_fd_sc_hd__nor2_1 _11757_ (.A(_04766_),
    .B(_04854_),
    .Y(_04942_));
 sky130_fd_sc_hd__a21oi_2 _11758_ (.A1(_04770_),
    .A2(_04942_),
    .B1(_04855_),
    .Y(_04943_));
 sky130_fd_sc_hd__xnor2_2 _11759_ (.A(_04941_),
    .B(_04943_),
    .Y(_04944_));
 sky130_fd_sc_hd__a41o_1 _11760_ (.A1(_04371_),
    .A2(_04773_),
    .A3(_04775_),
    .A4(_04858_),
    .B1(net86),
    .X(_04945_));
 sky130_fd_sc_hd__nand2_1 _11761_ (.A(_04944_),
    .B(_04945_),
    .Y(_04946_));
 sky130_fd_sc_hd__o21a_1 _11762_ (.A1(_04944_),
    .A2(_04945_),
    .B1(_02213_),
    .X(_04947_));
 sky130_fd_sc_hd__a21o_1 _11763_ (.A1(net20),
    .A2(_02198_),
    .B1(_02149_),
    .X(_04949_));
 sky130_fd_sc_hd__a31oi_1 _11764_ (.A1(net20),
    .A2(_02149_),
    .A3(_02198_),
    .B1(_02299_),
    .Y(_04950_));
 sky130_fd_sc_hd__a21o_1 _11765_ (.A1(_05582_),
    .A2(_04866_),
    .B1(_05563_),
    .X(_04951_));
 sky130_fd_sc_hd__mux2_1 _11766_ (.A0(_06338_),
    .A1(_04951_),
    .S(net299),
    .X(_04952_));
 sky130_fd_sc_hd__nand2_1 _11767_ (.A(_05501_),
    .B(_04952_),
    .Y(_04953_));
 sky130_fd_sc_hd__o211a_1 _11768_ (.A1(_05501_),
    .A2(_04952_),
    .B1(_04953_),
    .C1(net251),
    .X(_04954_));
 sky130_fd_sc_hd__nor2_1 _11769_ (.A(reg1_val[22]),
    .B(curr_PC[22]),
    .Y(_04955_));
 sky130_fd_sc_hd__nand2_1 _11770_ (.A(reg1_val[22]),
    .B(curr_PC[22]),
    .Y(_04956_));
 sky130_fd_sc_hd__and2b_1 _11771_ (.A_N(_04955_),
    .B(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__o21a_1 _11772_ (.A1(_04870_),
    .A2(_04874_),
    .B1(_04871_),
    .X(_04958_));
 sky130_fd_sc_hd__xnor2_1 _11773_ (.A(_04957_),
    .B(_04958_),
    .Y(_04960_));
 sky130_fd_sc_hd__nand2_1 _11774_ (.A(net242),
    .B(_03619_),
    .Y(_04961_));
 sky130_fd_sc_hd__o211a_1 _11775_ (.A1(net241),
    .A2(_04960_),
    .B1(_04961_),
    .C1(net215),
    .X(_04962_));
 sky130_fd_sc_hd__or2_1 _11776_ (.A(\div_shifter[53] ),
    .B(_04878_),
    .X(_04963_));
 sky130_fd_sc_hd__a21oi_1 _11777_ (.A1(net244),
    .A2(_04963_),
    .B1(\div_shifter[54] ),
    .Y(_04964_));
 sky130_fd_sc_hd__a311o_1 _11778_ (.A1(\div_shifter[54] ),
    .A2(net244),
    .A3(_04963_),
    .B1(_04964_),
    .C1(net248),
    .X(_04965_));
 sky130_fd_sc_hd__or2_1 _11779_ (.A(\div_res[21] ),
    .B(_04881_),
    .X(_04966_));
 sky130_fd_sc_hd__a21o_1 _11780_ (.A1(net23),
    .A2(_04966_),
    .B1(\div_res[22] ),
    .X(_04967_));
 sky130_fd_sc_hd__nand3_1 _11781_ (.A(\div_res[22] ),
    .B(net23),
    .C(_04966_),
    .Y(_04968_));
 sky130_fd_sc_hd__mux2_1 _11782_ (.A0(_02295_),
    .A1(net204),
    .S(_05479_),
    .X(_04969_));
 sky130_fd_sc_hd__a21oi_1 _11783_ (.A1(_02291_),
    .A2(_04969_),
    .B1(_05490_),
    .Y(_04971_));
 sky130_fd_sc_hd__a221o_1 _11784_ (.A1(_02217_),
    .A2(_03607_),
    .B1(_03620_),
    .B2(_02288_),
    .C1(_04971_),
    .X(_04972_));
 sky130_fd_sc_hd__a31o_1 _11785_ (.A1(_02305_),
    .A2(_04967_),
    .A3(_04968_),
    .B1(_04972_),
    .X(_04973_));
 sky130_fd_sc_hd__or4b_2 _11786_ (.A(_04954_),
    .B(_04962_),
    .C(_04973_),
    .D_N(_04965_),
    .X(_04974_));
 sky130_fd_sc_hd__a221o_1 _11787_ (.A1(_04946_),
    .A2(_04947_),
    .B1(_04949_),
    .B2(_04950_),
    .C1(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__a22o_1 _11788_ (.A1(_05458_),
    .A2(net212),
    .B1(_06427_),
    .B2(_04975_),
    .X(_04976_));
 sky130_fd_sc_hd__nand2_1 _11789_ (.A(curr_PC[22]),
    .B(_04893_),
    .Y(_04977_));
 sky130_fd_sc_hd__o21a_1 _11790_ (.A1(curr_PC[22]),
    .A2(_04893_),
    .B1(_06390_),
    .X(_04978_));
 sky130_fd_sc_hd__a22o_4 _11791_ (.A1(net258),
    .A2(_04976_),
    .B1(_04977_),
    .B2(_04978_),
    .X(dest_val[22]));
 sky130_fd_sc_hd__o21ai_1 _11792_ (.A1(_04924_),
    .A2(_04925_),
    .B1(_04928_),
    .Y(_04979_));
 sky130_fd_sc_hd__o22a_1 _11793_ (.A1(net18),
    .A2(net15),
    .B1(_00265_),
    .B2(net17),
    .X(_04981_));
 sky130_fd_sc_hd__xor2_1 _11794_ (.A(net112),
    .B(_04981_),
    .X(_04982_));
 sky130_fd_sc_hd__or2_1 _11795_ (.A(net106),
    .B(_04982_),
    .X(_04983_));
 sky130_fd_sc_hd__nand2_1 _11796_ (.A(net106),
    .B(_04982_),
    .Y(_04984_));
 sky130_fd_sc_hd__nand2_1 _11797_ (.A(_04983_),
    .B(_04984_),
    .Y(_04985_));
 sky130_fd_sc_hd__o22a_1 _11798_ (.A1(net13),
    .A2(net10),
    .B1(net4),
    .B2(net47),
    .X(_04986_));
 sky130_fd_sc_hd__xor2_1 _11799_ (.A(net108),
    .B(_04986_),
    .X(_04987_));
 sky130_fd_sc_hd__or2_1 _11800_ (.A(_04985_),
    .B(_04987_),
    .X(_04988_));
 sky130_fd_sc_hd__nand2_1 _11801_ (.A(_04985_),
    .B(_04987_),
    .Y(_04989_));
 sky130_fd_sc_hd__nand2_1 _11802_ (.A(_04988_),
    .B(_04989_),
    .Y(_04990_));
 sky130_fd_sc_hd__xor2_1 _11803_ (.A(_04911_),
    .B(_04990_),
    .X(_04992_));
 sky130_fd_sc_hd__nor2_1 _11804_ (.A(_04900_),
    .B(_04992_),
    .Y(_04993_));
 sky130_fd_sc_hd__and2_1 _11805_ (.A(_04900_),
    .B(_04992_),
    .X(_04994_));
 sky130_fd_sc_hd__nor2_1 _11806_ (.A(_04993_),
    .B(_04994_),
    .Y(_04995_));
 sky130_fd_sc_hd__o21a_1 _11807_ (.A1(_04906_),
    .A2(_04913_),
    .B1(_04903_),
    .X(_04996_));
 sky130_fd_sc_hd__o22a_1 _11808_ (.A1(net55),
    .A2(net8),
    .B1(net6),
    .B2(net58),
    .X(_04997_));
 sky130_fd_sc_hd__xnor2_1 _11809_ (.A(net31),
    .B(_04997_),
    .Y(_04998_));
 sky130_fd_sc_hd__o22a_1 _11810_ (.A1(net63),
    .A2(net11),
    .B1(net44),
    .B2(net61),
    .X(_04999_));
 sky130_fd_sc_hd__xor2_1 _11811_ (.A(net97),
    .B(_04999_),
    .X(_05000_));
 sky130_fd_sc_hd__and3b_1 _11812_ (.A_N(net65),
    .B(net33),
    .C(_05000_),
    .X(_05001_));
 sky130_fd_sc_hd__o21ba_1 _11813_ (.A1(net65),
    .A2(net31),
    .B1_N(_05000_),
    .X(_05003_));
 sky130_fd_sc_hd__or2_1 _11814_ (.A(_05001_),
    .B(_05003_),
    .X(_05004_));
 sky130_fd_sc_hd__nor2_1 _11815_ (.A(_04998_),
    .B(_05004_),
    .Y(_05005_));
 sky130_fd_sc_hd__and2_1 _11816_ (.A(_04998_),
    .B(_05004_),
    .X(_05006_));
 sky130_fd_sc_hd__nor2_1 _11817_ (.A(_05005_),
    .B(_05006_),
    .Y(_05007_));
 sky130_fd_sc_hd__o21a_1 _11818_ (.A1(_04920_),
    .A2(_04923_),
    .B1(_05007_),
    .X(_05008_));
 sky130_fd_sc_hd__nor3_1 _11819_ (.A(_04920_),
    .B(_04923_),
    .C(_05007_),
    .Y(_05009_));
 sky130_fd_sc_hd__nor2_1 _11820_ (.A(_05008_),
    .B(_05009_),
    .Y(_05010_));
 sky130_fd_sc_hd__and2b_1 _11821_ (.A_N(_04996_),
    .B(_05010_),
    .X(_05011_));
 sky130_fd_sc_hd__xnor2_1 _11822_ (.A(_04996_),
    .B(_05010_),
    .Y(_05012_));
 sky130_fd_sc_hd__and2_1 _11823_ (.A(_04995_),
    .B(_05012_),
    .X(_05014_));
 sky130_fd_sc_hd__nor2_1 _11824_ (.A(_04995_),
    .B(_05012_),
    .Y(_05015_));
 sky130_fd_sc_hd__or2_1 _11825_ (.A(_05014_),
    .B(_05015_),
    .X(_05016_));
 sky130_fd_sc_hd__and2b_1 _11826_ (.A_N(_05016_),
    .B(_04979_),
    .X(_05017_));
 sky130_fd_sc_hd__xor2_1 _11827_ (.A(_04979_),
    .B(_05016_),
    .X(_05018_));
 sky130_fd_sc_hd__nand3_1 _11828_ (.A(_04930_),
    .B(_04934_),
    .C(_05018_),
    .Y(_05019_));
 sky130_fd_sc_hd__a21oi_1 _11829_ (.A1(_04930_),
    .A2(_04934_),
    .B1(_05018_),
    .Y(_05020_));
 sky130_fd_sc_hd__inv_2 _11830_ (.A(_05020_),
    .Y(_05021_));
 sky130_fd_sc_hd__nand2_1 _11831_ (.A(_05019_),
    .B(_05021_),
    .Y(_05022_));
 sky130_fd_sc_hd__a21oi_1 _11832_ (.A1(_04941_),
    .A2(_04943_),
    .B1(_04939_),
    .Y(_05023_));
 sky130_fd_sc_hd__xnor2_2 _11833_ (.A(_05022_),
    .B(_05023_),
    .Y(_05025_));
 sky130_fd_sc_hd__and4_1 _11834_ (.A(_04773_),
    .B(_04775_),
    .C(_04858_),
    .D(_04944_),
    .X(_05026_));
 sky130_fd_sc_hd__a21o_1 _11835_ (.A1(_04371_),
    .A2(_05026_),
    .B1(net86),
    .X(_05027_));
 sky130_fd_sc_hd__nor2_1 _11836_ (.A(_05025_),
    .B(_05027_),
    .Y(_05028_));
 sky130_fd_sc_hd__a21o_1 _11837_ (.A1(_05025_),
    .A2(_05027_),
    .B1(_02214_),
    .X(_05029_));
 sky130_fd_sc_hd__and3_1 _11838_ (.A(net20),
    .B(_02148_),
    .C(_02199_),
    .X(_05030_));
 sky130_fd_sc_hd__a21oi_1 _11839_ (.A1(net20),
    .A2(_02199_),
    .B1(_02148_),
    .Y(_05031_));
 sky130_fd_sc_hd__or2_1 _11840_ (.A(_05030_),
    .B(_05031_),
    .X(_05032_));
 sky130_fd_sc_hd__a21o_1 _11841_ (.A1(_05501_),
    .A2(_04951_),
    .B1(_05479_),
    .X(_05033_));
 sky130_fd_sc_hd__mux2_1 _11842_ (.A0(_06340_),
    .A1(_05033_),
    .S(net299),
    .X(_05034_));
 sky130_fd_sc_hd__o21ai_1 _11843_ (.A1(_05425_),
    .A2(_05034_),
    .B1(_02292_),
    .Y(_05036_));
 sky130_fd_sc_hd__a21o_1 _11844_ (.A1(_05425_),
    .A2(_05034_),
    .B1(_05036_),
    .X(_05037_));
 sky130_fd_sc_hd__or2_1 _11845_ (.A(reg1_val[23]),
    .B(curr_PC[23]),
    .X(_05038_));
 sky130_fd_sc_hd__nand2_1 _11846_ (.A(reg1_val[23]),
    .B(curr_PC[23]),
    .Y(_05039_));
 sky130_fd_sc_hd__nand2_1 _11847_ (.A(_05038_),
    .B(_05039_),
    .Y(_05040_));
 sky130_fd_sc_hd__o21a_1 _11848_ (.A1(_04955_),
    .A2(_04958_),
    .B1(_04956_),
    .X(_05041_));
 sky130_fd_sc_hd__xnor2_1 _11849_ (.A(_05040_),
    .B(_05041_),
    .Y(_05042_));
 sky130_fd_sc_hd__mux2_1 _11850_ (.A0(_03495_),
    .A1(_05042_),
    .S(net264),
    .X(_05043_));
 sky130_fd_sc_hd__or2_1 _11851_ (.A(\div_shifter[54] ),
    .B(_04963_),
    .X(_05044_));
 sky130_fd_sc_hd__a21oi_1 _11852_ (.A1(net244),
    .A2(_05044_),
    .B1(\div_shifter[55] ),
    .Y(_05045_));
 sky130_fd_sc_hd__a31o_1 _11853_ (.A1(\div_shifter[55] ),
    .A2(net244),
    .A3(_05044_),
    .B1(net248),
    .X(_05047_));
 sky130_fd_sc_hd__or2_1 _11854_ (.A(\div_res[22] ),
    .B(_04966_),
    .X(_05048_));
 sky130_fd_sc_hd__a21oi_1 _11855_ (.A1(net24),
    .A2(_05048_),
    .B1(\div_res[23] ),
    .Y(_05049_));
 sky130_fd_sc_hd__a31o_1 _11856_ (.A1(\div_res[23] ),
    .A2(net24),
    .A3(_05048_),
    .B1(net202),
    .X(_05050_));
 sky130_fd_sc_hd__or2_1 _11857_ (.A(_05049_),
    .B(_05050_),
    .X(_05051_));
 sky130_fd_sc_hd__mux2_1 _11858_ (.A0(_02295_),
    .A1(net204),
    .S(_05404_),
    .X(_05052_));
 sky130_fd_sc_hd__a2bb2o_1 _11859_ (.A1_N(reg1_val[23]),
    .A2_N(_05382_),
    .B1(_02291_),
    .B2(_05052_),
    .X(_05053_));
 sky130_fd_sc_hd__o221a_1 _11860_ (.A1(net186),
    .A2(_03485_),
    .B1(_03495_),
    .B2(net182),
    .C1(_05053_),
    .X(_05054_));
 sky130_fd_sc_hd__o211a_1 _11861_ (.A1(_05045_),
    .A2(_05047_),
    .B1(_05051_),
    .C1(_05054_),
    .X(_05055_));
 sky130_fd_sc_hd__o211a_1 _11862_ (.A1(net214),
    .A2(_05043_),
    .B1(_05055_),
    .C1(_05037_),
    .X(_05056_));
 sky130_fd_sc_hd__o221a_1 _11863_ (.A1(_05028_),
    .A2(_05029_),
    .B1(_05032_),
    .B2(net250),
    .C1(_05056_),
    .X(_05058_));
 sky130_fd_sc_hd__o22a_1 _11864_ (.A1(_05371_),
    .A2(_06426_),
    .B1(_06428_),
    .B2(_05058_),
    .X(_05059_));
 sky130_fd_sc_hd__a21oi_1 _11865_ (.A1(curr_PC[22]),
    .A2(_04893_),
    .B1(curr_PC[23]),
    .Y(_05060_));
 sky130_fd_sc_hd__and3_1 _11866_ (.A(curr_PC[22]),
    .B(curr_PC[23]),
    .C(_04893_),
    .X(_05061_));
 sky130_fd_sc_hd__or3_1 _11867_ (.A(net261),
    .B(_05060_),
    .C(_05061_),
    .X(_05062_));
 sky130_fd_sc_hd__o21ai_4 _11868_ (.A1(_06390_),
    .A2(_05059_),
    .B1(_05062_),
    .Y(dest_val[23]));
 sky130_fd_sc_hd__nand3_1 _11869_ (.A(_04941_),
    .B(_05019_),
    .C(_05021_),
    .Y(_05063_));
 sky130_fd_sc_hd__a2111o_1 _11870_ (.A1(_04714_),
    .A2(_04715_),
    .B1(_04768_),
    .C1(_04856_),
    .D1(_05063_),
    .X(_05064_));
 sky130_fd_sc_hd__nand2_1 _11871_ (.A(_04939_),
    .B(_05019_),
    .Y(_05065_));
 sky130_fd_sc_hd__o311a_1 _11872_ (.A1(_04855_),
    .A2(_04942_),
    .A3(_05063_),
    .B1(_05065_),
    .C1(_05021_),
    .X(_05066_));
 sky130_fd_sc_hd__nand2_1 _11873_ (.A(_05064_),
    .B(_05066_),
    .Y(_05068_));
 sky130_fd_sc_hd__o21ai_1 _11874_ (.A1(_00305_),
    .A2(net4),
    .B1(net109),
    .Y(_05069_));
 sky130_fd_sc_hd__o31a_1 _11875_ (.A1(net109),
    .A2(_00303_),
    .A3(net4),
    .B1(_05069_),
    .X(_05070_));
 sky130_fd_sc_hd__nor2_1 _11876_ (.A(net57),
    .B(net32),
    .Y(_05071_));
 sky130_fd_sc_hd__xnor2_1 _11877_ (.A(_05070_),
    .B(_05071_),
    .Y(_05072_));
 sky130_fd_sc_hd__a21oi_1 _11878_ (.A1(_04983_),
    .A2(_04988_),
    .B1(_05072_),
    .Y(_05073_));
 sky130_fd_sc_hd__and3_1 _11879_ (.A(_04983_),
    .B(_04988_),
    .C(_05072_),
    .X(_05074_));
 sky130_fd_sc_hd__or2_1 _11880_ (.A(_05073_),
    .B(_05074_),
    .X(_05075_));
 sky130_fd_sc_hd__a31o_1 _11881_ (.A1(_04911_),
    .A2(_04988_),
    .A3(_04989_),
    .B1(_04993_),
    .X(_05076_));
 sky130_fd_sc_hd__o22a_1 _11882_ (.A1(net61),
    .A2(net12),
    .B1(net45),
    .B2(net18),
    .X(_05077_));
 sky130_fd_sc_hd__xnor2_1 _11883_ (.A(net97),
    .B(_05077_),
    .Y(_05079_));
 sky130_fd_sc_hd__o22a_1 _11884_ (.A1(net62),
    .A2(net8),
    .B1(net6),
    .B2(net54),
    .X(_05080_));
 sky130_fd_sc_hd__xnor2_1 _11885_ (.A(net31),
    .B(_05080_),
    .Y(_05081_));
 sky130_fd_sc_hd__o22a_1 _11886_ (.A1(net16),
    .A2(net15),
    .B1(net53),
    .B2(net10),
    .X(_05082_));
 sky130_fd_sc_hd__xor2_1 _11887_ (.A(_00248_),
    .B(_05082_),
    .X(_05083_));
 sky130_fd_sc_hd__nor2_1 _11888_ (.A(_05081_),
    .B(_05083_),
    .Y(_05084_));
 sky130_fd_sc_hd__and2_1 _11889_ (.A(_05081_),
    .B(_05083_),
    .X(_05085_));
 sky130_fd_sc_hd__or2_1 _11890_ (.A(_05084_),
    .B(_05085_),
    .X(_05086_));
 sky130_fd_sc_hd__nor2_1 _11891_ (.A(_05079_),
    .B(_05086_),
    .Y(_05087_));
 sky130_fd_sc_hd__and2_1 _11892_ (.A(_05079_),
    .B(_05086_),
    .X(_05088_));
 sky130_fd_sc_hd__nor2_1 _11893_ (.A(_05087_),
    .B(_05088_),
    .Y(_05090_));
 sky130_fd_sc_hd__o21a_1 _11894_ (.A1(_05001_),
    .A2(_05005_),
    .B1(_05090_),
    .X(_05091_));
 sky130_fd_sc_hd__nor3_1 _11895_ (.A(_05001_),
    .B(_05005_),
    .C(_05090_),
    .Y(_05092_));
 sky130_fd_sc_hd__nor2_1 _11896_ (.A(_05091_),
    .B(_05092_),
    .Y(_05093_));
 sky130_fd_sc_hd__xnor2_1 _11897_ (.A(_05076_),
    .B(_05093_),
    .Y(_05094_));
 sky130_fd_sc_hd__or2_1 _11898_ (.A(_05075_),
    .B(_05094_),
    .X(_05095_));
 sky130_fd_sc_hd__nand2_1 _11899_ (.A(_05075_),
    .B(_05094_),
    .Y(_05096_));
 sky130_fd_sc_hd__and2_1 _11900_ (.A(_05095_),
    .B(_05096_),
    .X(_05097_));
 sky130_fd_sc_hd__o21ai_1 _11901_ (.A1(_05008_),
    .A2(_05011_),
    .B1(_05097_),
    .Y(_05098_));
 sky130_fd_sc_hd__or3_1 _11902_ (.A(_05008_),
    .B(_05011_),
    .C(_05097_),
    .X(_05099_));
 sky130_fd_sc_hd__and2_1 _11903_ (.A(_05098_),
    .B(_05099_),
    .X(_05101_));
 sky130_fd_sc_hd__o21ai_4 _11904_ (.A1(_05014_),
    .A2(_05017_),
    .B1(_05101_),
    .Y(_05102_));
 sky130_fd_sc_hd__or3_1 _11905_ (.A(_05014_),
    .B(_05017_),
    .C(_05101_),
    .X(_05103_));
 sky130_fd_sc_hd__and2_1 _11906_ (.A(_05102_),
    .B(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__inv_2 _11907_ (.A(_05104_),
    .Y(_05105_));
 sky130_fd_sc_hd__a21o_1 _11908_ (.A1(_05064_),
    .A2(_05066_),
    .B1(_05105_),
    .X(_05106_));
 sky130_fd_sc_hd__xnor2_2 _11909_ (.A(_05068_),
    .B(_05104_),
    .Y(_05107_));
 sky130_fd_sc_hd__and3_1 _11910_ (.A(_04371_),
    .B(_05025_),
    .C(_05026_),
    .X(_05108_));
 sky130_fd_sc_hd__o21ai_1 _11911_ (.A1(net85),
    .A2(_05108_),
    .B1(_05107_),
    .Y(_05109_));
 sky130_fd_sc_hd__o31a_1 _11912_ (.A1(net85),
    .A2(_05107_),
    .A3(_05108_),
    .B1(_02213_),
    .X(_05110_));
 sky130_fd_sc_hd__nand2_1 _11913_ (.A(_05109_),
    .B(_05110_),
    .Y(_05112_));
 sky130_fd_sc_hd__and3_1 _11914_ (.A(net21),
    .B(_02200_),
    .C(_02202_),
    .X(_05113_));
 sky130_fd_sc_hd__a21oi_1 _11915_ (.A1(net21),
    .A2(_02200_),
    .B1(_02202_),
    .Y(_05114_));
 sky130_fd_sc_hd__a21o_1 _11916_ (.A1(_05425_),
    .A2(_05033_),
    .B1(_05404_),
    .X(_05115_));
 sky130_fd_sc_hd__mux2_1 _11917_ (.A0(_06342_),
    .A1(_05115_),
    .S(net300),
    .X(_05116_));
 sky130_fd_sc_hd__nor2_1 _11918_ (.A(_05154_),
    .B(_05116_),
    .Y(_05117_));
 sky130_fd_sc_hd__a21o_1 _11919_ (.A1(_05154_),
    .A2(_05116_),
    .B1(_02293_),
    .X(_05118_));
 sky130_fd_sc_hd__o21a_1 _11920_ (.A1(_05040_),
    .A2(_05041_),
    .B1(_05039_),
    .X(_05119_));
 sky130_fd_sc_hd__nor2_1 _11921_ (.A(reg1_val[24]),
    .B(curr_PC[24]),
    .Y(_05120_));
 sky130_fd_sc_hd__nand2_1 _11922_ (.A(reg1_val[24]),
    .B(curr_PC[24]),
    .Y(_05121_));
 sky130_fd_sc_hd__and2b_1 _11923_ (.A_N(_05120_),
    .B(_05121_),
    .X(_05123_));
 sky130_fd_sc_hd__xnor2_1 _11924_ (.A(_05119_),
    .B(_05123_),
    .Y(_05124_));
 sky130_fd_sc_hd__nor2_1 _11925_ (.A(net242),
    .B(_05124_),
    .Y(_05125_));
 sky130_fd_sc_hd__a211o_1 _11926_ (.A1(net242),
    .A2(_03364_),
    .B1(_05125_),
    .C1(net214),
    .X(_05126_));
 sky130_fd_sc_hd__or2_1 _11927_ (.A(\div_res[23] ),
    .B(_05048_),
    .X(_05127_));
 sky130_fd_sc_hd__a21oi_1 _11928_ (.A1(net24),
    .A2(_05127_),
    .B1(\div_res[24] ),
    .Y(_05128_));
 sky130_fd_sc_hd__a31o_1 _11929_ (.A1(\div_res[24] ),
    .A2(net24),
    .A3(_05127_),
    .B1(net202),
    .X(_05129_));
 sky130_fd_sc_hd__or2_1 _11930_ (.A(_05128_),
    .B(_05129_),
    .X(_05130_));
 sky130_fd_sc_hd__or3_1 _11931_ (.A(\div_shifter[55] ),
    .B(\div_shifter[54] ),
    .C(_04963_),
    .X(_05131_));
 sky130_fd_sc_hd__a21oi_1 _11932_ (.A1(net244),
    .A2(_05131_),
    .B1(\div_shifter[56] ),
    .Y(_05132_));
 sky130_fd_sc_hd__a31o_1 _11933_ (.A1(\div_shifter[56] ),
    .A2(net244),
    .A3(_05131_),
    .B1(net248),
    .X(_05134_));
 sky130_fd_sc_hd__a21o_1 _11934_ (.A1(_05133_),
    .A2(_02294_),
    .B1(net205),
    .X(_05135_));
 sky130_fd_sc_hd__nand2_1 _11935_ (.A(_05144_),
    .B(_05135_),
    .Y(_05136_));
 sky130_fd_sc_hd__o221a_1 _11936_ (.A1(_05111_),
    .A2(_06426_),
    .B1(net204),
    .B2(_05133_),
    .C1(_05136_),
    .X(_05137_));
 sky130_fd_sc_hd__o221a_1 _11937_ (.A1(net186),
    .A2(_03350_),
    .B1(_03364_),
    .B2(net183),
    .C1(_05137_),
    .X(_05138_));
 sky130_fd_sc_hd__o211a_1 _11938_ (.A1(_05132_),
    .A2(_05134_),
    .B1(_05138_),
    .C1(_05130_),
    .X(_05139_));
 sky130_fd_sc_hd__o211a_1 _11939_ (.A1(_05117_),
    .A2(_05118_),
    .B1(_05126_),
    .C1(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__o311a_1 _11940_ (.A1(net250),
    .A2(_05113_),
    .A3(_05114_),
    .B1(_05140_),
    .C1(_05112_),
    .X(_05141_));
 sky130_fd_sc_hd__and2_2 _11941_ (.A(curr_PC[24]),
    .B(_05061_),
    .X(_05142_));
 sky130_fd_sc_hd__o21ai_1 _11942_ (.A1(curr_PC[24]),
    .A2(_05061_),
    .B1(net262),
    .Y(_05143_));
 sky130_fd_sc_hd__o22ai_4 _11943_ (.A1(_06390_),
    .A2(_05141_),
    .B1(_05142_),
    .B2(_05143_),
    .Y(dest_val[24]));
 sky130_fd_sc_hd__a21o_1 _11944_ (.A1(_05076_),
    .A2(_05093_),
    .B1(_05091_),
    .X(_05145_));
 sky130_fd_sc_hd__o22a_1 _11945_ (.A1(net60),
    .A2(net7),
    .B1(net5),
    .B2(net62),
    .X(_05146_));
 sky130_fd_sc_hd__xnor2_1 _11946_ (.A(net30),
    .B(_05146_),
    .Y(_05147_));
 sky130_fd_sc_hd__nor2_1 _11947_ (.A(_05070_),
    .B(_05147_),
    .Y(_05148_));
 sky130_fd_sc_hd__and2_1 _11948_ (.A(_05070_),
    .B(_05147_),
    .X(_05149_));
 sky130_fd_sc_hd__nor2_1 _11949_ (.A(_05148_),
    .B(_05149_),
    .Y(_05150_));
 sky130_fd_sc_hd__nor2_1 _11950_ (.A(net54),
    .B(net30),
    .Y(_05151_));
 sky130_fd_sc_hd__xnor2_1 _11951_ (.A(_05150_),
    .B(_05151_),
    .Y(_05152_));
 sky130_fd_sc_hd__a21o_1 _11952_ (.A1(_05070_),
    .A2(_05071_),
    .B1(_05073_),
    .X(_05153_));
 sky130_fd_sc_hd__o22a_1 _11953_ (.A1(net18),
    .A2(net11),
    .B1(net46),
    .B2(net16),
    .X(_05155_));
 sky130_fd_sc_hd__xnor2_1 _11954_ (.A(net96),
    .B(_05155_),
    .Y(_05156_));
 sky130_fd_sc_hd__nor2_1 _11955_ (.A(net110),
    .B(_05156_),
    .Y(_05157_));
 sky130_fd_sc_hd__and2_1 _11956_ (.A(_00255_),
    .B(_05156_),
    .X(_05158_));
 sky130_fd_sc_hd__nor2_1 _11957_ (.A(_05157_),
    .B(_05158_),
    .Y(_05159_));
 sky130_fd_sc_hd__o22a_1 _11958_ (.A1(net15),
    .A2(net10),
    .B1(_00757_),
    .B2(net53),
    .X(_05160_));
 sky130_fd_sc_hd__xnor2_1 _11959_ (.A(net113),
    .B(_05160_),
    .Y(_05161_));
 sky130_fd_sc_hd__and2_1 _11960_ (.A(_05159_),
    .B(_05161_),
    .X(_05162_));
 sky130_fd_sc_hd__nor2_1 _11961_ (.A(_05159_),
    .B(_05161_),
    .Y(_05163_));
 sky130_fd_sc_hd__nor2_1 _11962_ (.A(_05162_),
    .B(_05163_),
    .Y(_05164_));
 sky130_fd_sc_hd__o21a_1 _11963_ (.A1(_05084_),
    .A2(_05087_),
    .B1(_05164_),
    .X(_05166_));
 sky130_fd_sc_hd__nor3_1 _11964_ (.A(_05084_),
    .B(_05087_),
    .C(_05164_),
    .Y(_05167_));
 sky130_fd_sc_hd__nor2_1 _11965_ (.A(_05166_),
    .B(_05167_),
    .Y(_05168_));
 sky130_fd_sc_hd__xnor2_1 _11966_ (.A(_05153_),
    .B(_05168_),
    .Y(_05169_));
 sky130_fd_sc_hd__nor2_1 _11967_ (.A(_05152_),
    .B(_05169_),
    .Y(_05170_));
 sky130_fd_sc_hd__and2_1 _11968_ (.A(_05152_),
    .B(_05169_),
    .X(_05171_));
 sky130_fd_sc_hd__nor2_1 _11969_ (.A(_05170_),
    .B(_05171_),
    .Y(_05172_));
 sky130_fd_sc_hd__xnor2_1 _11970_ (.A(_05145_),
    .B(_05172_),
    .Y(_05173_));
 sky130_fd_sc_hd__a21o_1 _11971_ (.A1(_05095_),
    .A2(_05098_),
    .B1(_05173_),
    .X(_05174_));
 sky130_fd_sc_hd__inv_2 _11972_ (.A(_05174_),
    .Y(_05175_));
 sky130_fd_sc_hd__and3_1 _11973_ (.A(_05095_),
    .B(_05098_),
    .C(_05173_),
    .X(_05177_));
 sky130_fd_sc_hd__nor2_1 _11974_ (.A(_05175_),
    .B(_05177_),
    .Y(_05178_));
 sky130_fd_sc_hd__inv_2 _11975_ (.A(_05178_),
    .Y(_05179_));
 sky130_fd_sc_hd__nand3_1 _11976_ (.A(_05102_),
    .B(_05106_),
    .C(_05178_),
    .Y(_05180_));
 sky130_fd_sc_hd__a21o_1 _11977_ (.A1(_05102_),
    .A2(_05106_),
    .B1(_05178_),
    .X(_05181_));
 sky130_fd_sc_hd__and2_1 _11978_ (.A(_05180_),
    .B(_05181_),
    .X(_05182_));
 sky130_fd_sc_hd__a21o_1 _11979_ (.A1(_05107_),
    .A2(_05108_),
    .B1(net85),
    .X(_05183_));
 sky130_fd_sc_hd__or2_1 _11980_ (.A(_05182_),
    .B(_05183_),
    .X(_05184_));
 sky130_fd_sc_hd__a21oi_1 _11981_ (.A1(_05182_),
    .A2(_05183_),
    .B1(_02214_),
    .Y(_05185_));
 sky130_fd_sc_hd__a21oi_1 _11982_ (.A1(net21),
    .A2(_02203_),
    .B1(_02145_),
    .Y(_05186_));
 sky130_fd_sc_hd__and3_1 _11983_ (.A(net21),
    .B(_02145_),
    .C(_02203_),
    .X(_05188_));
 sky130_fd_sc_hd__nor2_1 _11984_ (.A(_05186_),
    .B(_05188_),
    .Y(_05189_));
 sky130_fd_sc_hd__a21bo_1 _11985_ (.A1(_05144_),
    .A2(_05115_),
    .B1_N(_05133_),
    .X(_05190_));
 sky130_fd_sc_hd__and2_1 _11986_ (.A(net299),
    .B(_05190_),
    .X(_05191_));
 sky130_fd_sc_hd__a31o_1 _11987_ (.A1(net305),
    .A2(_06350_),
    .A3(_06358_),
    .B1(_05191_),
    .X(_05192_));
 sky130_fd_sc_hd__nor2_1 _11988_ (.A(_05013_),
    .B(_05192_),
    .Y(_05193_));
 sky130_fd_sc_hd__a21o_1 _11989_ (.A1(_05013_),
    .A2(_05192_),
    .B1(_02293_),
    .X(_05194_));
 sky130_fd_sc_hd__o21a_1 _11990_ (.A1(_05119_),
    .A2(_05120_),
    .B1(_05121_),
    .X(_05195_));
 sky130_fd_sc_hd__nor2_1 _11991_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .Y(_05196_));
 sky130_fd_sc_hd__nand2_1 _11992_ (.A(reg1_val[25]),
    .B(curr_PC[25]),
    .Y(_05197_));
 sky130_fd_sc_hd__and2b_1 _11993_ (.A_N(_05196_),
    .B(_05197_),
    .X(_05199_));
 sky130_fd_sc_hd__nor2_1 _11994_ (.A(_05195_),
    .B(_05199_),
    .Y(_05200_));
 sky130_fd_sc_hd__a21o_1 _11995_ (.A1(_05195_),
    .A2(_05199_),
    .B1(net242),
    .X(_05201_));
 sky130_fd_sc_hd__a21oi_1 _11996_ (.A1(net242),
    .A2(_03235_),
    .B1(net214),
    .Y(_05202_));
 sky130_fd_sc_hd__o21ai_1 _11997_ (.A1(_05200_),
    .A2(_05201_),
    .B1(_05202_),
    .Y(_05203_));
 sky130_fd_sc_hd__or2_1 _11998_ (.A(\div_shifter[56] ),
    .B(_05131_),
    .X(_05204_));
 sky130_fd_sc_hd__a21oi_1 _11999_ (.A1(net245),
    .A2(_05204_),
    .B1(\div_shifter[57] ),
    .Y(_05205_));
 sky130_fd_sc_hd__a311o_1 _12000_ (.A1(\div_shifter[57] ),
    .A2(net245),
    .A3(_05204_),
    .B1(_05205_),
    .C1(net248),
    .X(_05206_));
 sky130_fd_sc_hd__or2_1 _12001_ (.A(\div_res[24] ),
    .B(_05127_),
    .X(_05207_));
 sky130_fd_sc_hd__a21oi_1 _12002_ (.A1(net24),
    .A2(_05207_),
    .B1(\div_res[25] ),
    .Y(_05208_));
 sky130_fd_sc_hd__a311o_1 _12003_ (.A1(\div_res[25] ),
    .A2(net24),
    .A3(_05207_),
    .B1(_05208_),
    .C1(net203),
    .X(_05210_));
 sky130_fd_sc_hd__a21o_1 _12004_ (.A1(_04991_),
    .A2(_02294_),
    .B1(net205),
    .X(_05211_));
 sky130_fd_sc_hd__nand2_1 _12005_ (.A(_05002_),
    .B(_05211_),
    .Y(_05212_));
 sky130_fd_sc_hd__o221a_1 _12006_ (.A1(_04980_),
    .A2(_06426_),
    .B1(net204),
    .B2(_04991_),
    .C1(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__o221a_1 _12007_ (.A1(net186),
    .A2(_03222_),
    .B1(_03235_),
    .B2(net183),
    .C1(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__and4_1 _12008_ (.A(_05203_),
    .B(_05206_),
    .C(_05210_),
    .D(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__o21ai_2 _12009_ (.A1(_05193_),
    .A2(_05194_),
    .B1(_05215_),
    .Y(_05216_));
 sky130_fd_sc_hd__a221o_1 _12010_ (.A1(_05184_),
    .A2(_05185_),
    .B1(_05189_),
    .B2(_02298_),
    .C1(_05216_),
    .X(_05217_));
 sky130_fd_sc_hd__or2_1 _12011_ (.A(curr_PC[25]),
    .B(_05142_),
    .X(_05218_));
 sky130_fd_sc_hd__a21oi_1 _12012_ (.A1(curr_PC[25]),
    .A2(_05142_),
    .B1(net261),
    .Y(_05219_));
 sky130_fd_sc_hd__a22o_4 _12013_ (.A1(net261),
    .A2(_05217_),
    .B1(_05218_),
    .B2(_05219_),
    .X(dest_val[25]));
 sky130_fd_sc_hd__a21o_1 _12014_ (.A1(_05150_),
    .A2(_05151_),
    .B1(_05148_),
    .X(_05221_));
 sky130_fd_sc_hd__o22a_1 _12015_ (.A1(net16),
    .A2(net11),
    .B1(net46),
    .B2(net10),
    .X(_05222_));
 sky130_fd_sc_hd__xnor2_1 _12016_ (.A(net98),
    .B(_05222_),
    .Y(_05223_));
 sky130_fd_sc_hd__o31ai_1 _12017_ (.A1(net110),
    .A2(_00256_),
    .A3(net4),
    .B1(_00248_),
    .Y(_05224_));
 sky130_fd_sc_hd__o21a_1 _12018_ (.A1(_00257_),
    .A2(net4),
    .B1(_05224_),
    .X(_05225_));
 sky130_fd_sc_hd__nand2_1 _12019_ (.A(_05223_),
    .B(_05225_),
    .Y(_05226_));
 sky130_fd_sc_hd__or2_1 _12020_ (.A(_05223_),
    .B(_05225_),
    .X(_05227_));
 sky130_fd_sc_hd__nand2_1 _12021_ (.A(_05226_),
    .B(_05227_),
    .Y(_05228_));
 sky130_fd_sc_hd__o21a_1 _12022_ (.A1(_05157_),
    .A2(_05162_),
    .B1(_05228_),
    .X(_05229_));
 sky130_fd_sc_hd__nor3_1 _12023_ (.A(_05157_),
    .B(_05162_),
    .C(_05228_),
    .Y(_05231_));
 sky130_fd_sc_hd__nor2_1 _12024_ (.A(_05229_),
    .B(_05231_),
    .Y(_05232_));
 sky130_fd_sc_hd__and2_1 _12025_ (.A(_05221_),
    .B(_05232_),
    .X(_05233_));
 sky130_fd_sc_hd__or2_1 _12026_ (.A(_05221_),
    .B(_05232_),
    .X(_05234_));
 sky130_fd_sc_hd__and2b_1 _12027_ (.A_N(_05233_),
    .B(_05234_),
    .X(_05235_));
 sky130_fd_sc_hd__o22a_1 _12028_ (.A1(net18),
    .A2(net8),
    .B1(net5),
    .B2(net61),
    .X(_05236_));
 sky130_fd_sc_hd__nand2_1 _12029_ (.A(net62),
    .B(net33),
    .Y(_05237_));
 sky130_fd_sc_hd__xor2_1 _12030_ (.A(_05236_),
    .B(_05237_),
    .X(_05238_));
 sky130_fd_sc_hd__nand2_1 _12031_ (.A(_05235_),
    .B(_05238_),
    .Y(_05239_));
 sky130_fd_sc_hd__or2_1 _12032_ (.A(_05235_),
    .B(_05238_),
    .X(_05240_));
 sky130_fd_sc_hd__nand2_1 _12033_ (.A(_05239_),
    .B(_05240_),
    .Y(_05242_));
 sky130_fd_sc_hd__a21oi_1 _12034_ (.A1(_05153_),
    .A2(_05168_),
    .B1(_05166_),
    .Y(_05243_));
 sky130_fd_sc_hd__or2_1 _12035_ (.A(_05242_),
    .B(_05243_),
    .X(_05244_));
 sky130_fd_sc_hd__nand2_1 _12036_ (.A(_05242_),
    .B(_05243_),
    .Y(_05245_));
 sky130_fd_sc_hd__nand2_1 _12037_ (.A(_05244_),
    .B(_05245_),
    .Y(_05246_));
 sky130_fd_sc_hd__a21oi_1 _12038_ (.A1(_05145_),
    .A2(_05172_),
    .B1(_05170_),
    .Y(_05247_));
 sky130_fd_sc_hd__nor2_1 _12039_ (.A(_05246_),
    .B(_05247_),
    .Y(_05248_));
 sky130_fd_sc_hd__and2_1 _12040_ (.A(_05246_),
    .B(_05247_),
    .X(_05249_));
 sky130_fd_sc_hd__or2_1 _12041_ (.A(_05248_),
    .B(_05249_),
    .X(_05250_));
 sky130_fd_sc_hd__a21o_1 _12042_ (.A1(_05102_),
    .A2(_05174_),
    .B1(_05177_),
    .X(_05251_));
 sky130_fd_sc_hd__a311oi_2 _12043_ (.A1(_05102_),
    .A2(_05106_),
    .A3(_05174_),
    .B1(_05177_),
    .C1(_05250_),
    .Y(_05253_));
 sky130_fd_sc_hd__o211a_1 _12044_ (.A1(_05106_),
    .A2(_05179_),
    .B1(_05250_),
    .C1(_05251_),
    .X(_05254_));
 sky130_fd_sc_hd__or2_1 _12045_ (.A(_05253_),
    .B(_05254_),
    .X(_05255_));
 sky130_fd_sc_hd__a31o_1 _12046_ (.A1(_05107_),
    .A2(_05108_),
    .A3(_05182_),
    .B1(net85),
    .X(_05256_));
 sky130_fd_sc_hd__nand2_1 _12047_ (.A(_05255_),
    .B(_05256_),
    .Y(_05257_));
 sky130_fd_sc_hd__o21a_1 _12048_ (.A1(_05255_),
    .A2(_05256_),
    .B1(_02213_),
    .X(_05258_));
 sky130_fd_sc_hd__a21oi_1 _12049_ (.A1(net22),
    .A2(_02205_),
    .B1(_02141_),
    .Y(_05259_));
 sky130_fd_sc_hd__a31o_1 _12050_ (.A1(net22),
    .A2(_02141_),
    .A3(_02205_),
    .B1(net250),
    .X(_05260_));
 sky130_fd_sc_hd__nor2_1 _12051_ (.A(_05259_),
    .B(_05260_),
    .Y(_05261_));
 sky130_fd_sc_hd__a21bo_1 _12052_ (.A1(_05002_),
    .A2(_05190_),
    .B1_N(_04991_),
    .X(_05262_));
 sky130_fd_sc_hd__and2_1 _12053_ (.A(net299),
    .B(_05262_),
    .X(_05264_));
 sky130_fd_sc_hd__a31o_1 _12054_ (.A1(net306),
    .A2(_06349_),
    .A3(_06359_),
    .B1(_05264_),
    .X(_05265_));
 sky130_fd_sc_hd__nand2_1 _12055_ (.A(_04861_),
    .B(_05265_),
    .Y(_05266_));
 sky130_fd_sc_hd__or2_1 _12056_ (.A(_04861_),
    .B(_05265_),
    .X(_05267_));
 sky130_fd_sc_hd__o21a_1 _12057_ (.A1(_05195_),
    .A2(_05196_),
    .B1(_05197_),
    .X(_05268_));
 sky130_fd_sc_hd__nor2_1 _12058_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .Y(_05269_));
 sky130_fd_sc_hd__nand2_1 _12059_ (.A(reg1_val[26]),
    .B(curr_PC[26]),
    .Y(_05270_));
 sky130_fd_sc_hd__nand2b_1 _12060_ (.A_N(_05269_),
    .B(_05270_),
    .Y(_05271_));
 sky130_fd_sc_hd__xnor2_1 _12061_ (.A(_05268_),
    .B(_05271_),
    .Y(_05272_));
 sky130_fd_sc_hd__mux2_1 _12062_ (.A0(_03100_),
    .A1(_05272_),
    .S(net264),
    .X(_05273_));
 sky130_fd_sc_hd__or2_1 _12063_ (.A(\div_shifter[57] ),
    .B(_05204_),
    .X(_05275_));
 sky130_fd_sc_hd__a21oi_1 _12064_ (.A1(net247),
    .A2(_05275_),
    .B1(\div_shifter[58] ),
    .Y(_05276_));
 sky130_fd_sc_hd__a31o_1 _12065_ (.A1(\div_shifter[58] ),
    .A2(net247),
    .A3(_05275_),
    .B1(net248),
    .X(_05277_));
 sky130_fd_sc_hd__or2_1 _12066_ (.A(_05276_),
    .B(_05277_),
    .X(_05278_));
 sky130_fd_sc_hd__or2_1 _12067_ (.A(\div_res[25] ),
    .B(_05207_),
    .X(_05279_));
 sky130_fd_sc_hd__a21oi_1 _12068_ (.A1(net26),
    .A2(_05279_),
    .B1(\div_res[26] ),
    .Y(_05280_));
 sky130_fd_sc_hd__a31o_1 _12069_ (.A1(\div_res[26] ),
    .A2(net26),
    .A3(_05279_),
    .B1(net203),
    .X(_05281_));
 sky130_fd_sc_hd__a21o_1 _12070_ (.A1(_04839_),
    .A2(_02294_),
    .B1(net205),
    .X(_05282_));
 sky130_fd_sc_hd__a2bb2o_1 _12071_ (.A1_N(_04839_),
    .A2_N(_02301_),
    .B1(net212),
    .B2(_04828_),
    .X(_05283_));
 sky130_fd_sc_hd__a21oi_1 _12072_ (.A1(_04850_),
    .A2(_05282_),
    .B1(_05283_),
    .Y(_05284_));
 sky130_fd_sc_hd__o221a_1 _12073_ (.A1(net186),
    .A2(_03088_),
    .B1(_03100_),
    .B2(net183),
    .C1(_05284_),
    .X(_05286_));
 sky130_fd_sc_hd__o211a_1 _12074_ (.A1(_05280_),
    .A2(_05281_),
    .B1(_05286_),
    .C1(_05278_),
    .X(_05287_));
 sky130_fd_sc_hd__o21ai_1 _12075_ (.A1(_06413_),
    .A2(_05273_),
    .B1(_05287_),
    .Y(_05288_));
 sky130_fd_sc_hd__a31o_1 _12076_ (.A1(net251),
    .A2(_05266_),
    .A3(_05267_),
    .B1(_05288_),
    .X(_05289_));
 sky130_fd_sc_hd__a211o_1 _12077_ (.A1(_05257_),
    .A2(_05258_),
    .B1(_05261_),
    .C1(_05289_),
    .X(_05290_));
 sky130_fd_sc_hd__a21oi_1 _12078_ (.A1(curr_PC[25]),
    .A2(_05142_),
    .B1(curr_PC[26]),
    .Y(_05291_));
 sky130_fd_sc_hd__and3_1 _12079_ (.A(curr_PC[25]),
    .B(curr_PC[26]),
    .C(_05142_),
    .X(_05292_));
 sky130_fd_sc_hd__or2_1 _12080_ (.A(net261),
    .B(_05292_),
    .X(_05293_));
 sky130_fd_sc_hd__a2bb2o_4 _12081_ (.A1_N(_05291_),
    .A2_N(_05293_),
    .B1(net261),
    .B2(_05290_),
    .X(dest_val[26]));
 sky130_fd_sc_hd__xor2_1 _12082_ (.A(curr_PC[27]),
    .B(_05292_),
    .X(_05294_));
 sky130_fd_sc_hd__o22a_1 _12083_ (.A1(net16),
    .A2(net8),
    .B1(net6),
    .B2(net18),
    .X(_05296_));
 sky130_fd_sc_hd__xnor2_1 _12084_ (.A(net32),
    .B(_05296_),
    .Y(_05297_));
 sky130_fd_sc_hd__or2_1 _12085_ (.A(net113),
    .B(_05297_),
    .X(_05298_));
 sky130_fd_sc_hd__nand2_1 _12086_ (.A(net111),
    .B(_05297_),
    .Y(_05299_));
 sky130_fd_sc_hd__and2_1 _12087_ (.A(_05298_),
    .B(_05299_),
    .X(_05300_));
 sky130_fd_sc_hd__o22a_1 _12088_ (.A1(net12),
    .A2(net10),
    .B1(net3),
    .B2(net44),
    .X(_05301_));
 sky130_fd_sc_hd__xnor2_1 _12089_ (.A(net96),
    .B(_05301_),
    .Y(_05302_));
 sky130_fd_sc_hd__inv_2 _12090_ (.A(_05302_),
    .Y(_05303_));
 sky130_fd_sc_hd__nand2_1 _12091_ (.A(_05300_),
    .B(_05303_),
    .Y(_05304_));
 sky130_fd_sc_hd__or2_1 _12092_ (.A(_05300_),
    .B(_05303_),
    .X(_05305_));
 sky130_fd_sc_hd__and2_1 _12093_ (.A(_05304_),
    .B(_05305_),
    .X(_05307_));
 sky130_fd_sc_hd__nor2_1 _12094_ (.A(net61),
    .B(net30),
    .Y(_05308_));
 sky130_fd_sc_hd__or3b_1 _12095_ (.A(net62),
    .B(net32),
    .C_N(_05236_),
    .X(_05309_));
 sky130_fd_sc_hd__mux2_1 _12096_ (.A0(net61),
    .A1(_05308_),
    .S(_05309_),
    .X(_05310_));
 sky130_fd_sc_hd__xor2_1 _12097_ (.A(_05226_),
    .B(_05310_),
    .X(_05311_));
 sky130_fd_sc_hd__and3_1 _12098_ (.A(_05304_),
    .B(_05305_),
    .C(_05311_),
    .X(_05312_));
 sky130_fd_sc_hd__nor2_1 _12099_ (.A(_05307_),
    .B(_05311_),
    .Y(_05313_));
 sky130_fd_sc_hd__nor2_1 _12100_ (.A(_05312_),
    .B(_05313_),
    .Y(_05314_));
 sky130_fd_sc_hd__o21a_1 _12101_ (.A1(_05229_),
    .A2(_05233_),
    .B1(_05314_),
    .X(_05315_));
 sky130_fd_sc_hd__nor3_1 _12102_ (.A(_05229_),
    .B(_05233_),
    .C(_05314_),
    .Y(_05316_));
 sky130_fd_sc_hd__or2_1 _12103_ (.A(_05315_),
    .B(_05316_),
    .X(_05318_));
 sky130_fd_sc_hd__nand3_1 _12104_ (.A(_05239_),
    .B(_05244_),
    .C(_05318_),
    .Y(_05319_));
 sky130_fd_sc_hd__a21o_1 _12105_ (.A1(_05239_),
    .A2(_05244_),
    .B1(_05318_),
    .X(_05320_));
 sky130_fd_sc_hd__nand2_1 _12106_ (.A(_05319_),
    .B(_05320_),
    .Y(_05321_));
 sky130_fd_sc_hd__nor2_1 _12107_ (.A(_05248_),
    .B(_05253_),
    .Y(_05322_));
 sky130_fd_sc_hd__xnor2_2 _12108_ (.A(_05321_),
    .B(_05322_),
    .Y(_05323_));
 sky130_fd_sc_hd__o2111a_1 _12109_ (.A1(_05253_),
    .A2(_05254_),
    .B1(_05107_),
    .C1(_05180_),
    .D1(_05181_),
    .X(_05324_));
 sky130_fd_sc_hd__and4_2 _12110_ (.A(_04371_),
    .B(_05025_),
    .C(_05026_),
    .D(_05324_),
    .X(_05325_));
 sky130_fd_sc_hd__o21ai_1 _12111_ (.A1(net85),
    .A2(_05325_),
    .B1(_05323_),
    .Y(_05326_));
 sky130_fd_sc_hd__or3_1 _12112_ (.A(net85),
    .B(_05323_),
    .C(_05325_),
    .X(_05327_));
 sky130_fd_sc_hd__and3_1 _12113_ (.A(_02213_),
    .B(_05326_),
    .C(_05327_),
    .X(_05329_));
 sky130_fd_sc_hd__a21bo_1 _12114_ (.A1(_04850_),
    .A2(_05262_),
    .B1_N(_04839_),
    .X(_05330_));
 sky130_fd_sc_hd__and3_1 _12115_ (.A(net306),
    .B(_06348_),
    .C(_06360_),
    .X(_05331_));
 sky130_fd_sc_hd__a21oi_1 _12116_ (.A1(net299),
    .A2(_05330_),
    .B1(_05331_),
    .Y(_05332_));
 sky130_fd_sc_hd__xnor2_1 _12117_ (.A(_04948_),
    .B(_05332_),
    .Y(_05333_));
 sky130_fd_sc_hd__o21ai_1 _12118_ (.A1(net85),
    .A2(_02206_),
    .B1(_02208_),
    .Y(_05334_));
 sky130_fd_sc_hd__o311a_1 _12119_ (.A1(net85),
    .A2(_02206_),
    .A3(_02208_),
    .B1(_02298_),
    .C1(_05334_),
    .X(_05335_));
 sky130_fd_sc_hd__o21a_1 _12120_ (.A1(_05268_),
    .A2(_05269_),
    .B1(_05270_),
    .X(_05336_));
 sky130_fd_sc_hd__nor2_1 _12121_ (.A(reg1_val[27]),
    .B(curr_PC[27]),
    .Y(_05337_));
 sky130_fd_sc_hd__nand2_1 _12122_ (.A(reg1_val[27]),
    .B(curr_PC[27]),
    .Y(_05338_));
 sky130_fd_sc_hd__nand2b_1 _12123_ (.A_N(_05337_),
    .B(_05338_),
    .Y(_05340_));
 sky130_fd_sc_hd__xnor2_1 _12124_ (.A(_05336_),
    .B(_05340_),
    .Y(_05341_));
 sky130_fd_sc_hd__mux2_1 _12125_ (.A0(_02964_),
    .A1(_05341_),
    .S(net263),
    .X(_05342_));
 sky130_fd_sc_hd__or2_1 _12126_ (.A(\div_shifter[58] ),
    .B(_05275_),
    .X(_05343_));
 sky130_fd_sc_hd__a21oi_1 _12127_ (.A1(net247),
    .A2(_05343_),
    .B1(\div_shifter[59] ),
    .Y(_05344_));
 sky130_fd_sc_hd__a311o_1 _12128_ (.A1(\div_shifter[59] ),
    .A2(net247),
    .A3(_05343_),
    .B1(_05344_),
    .C1(net249),
    .X(_05345_));
 sky130_fd_sc_hd__or2_1 _12129_ (.A(\div_res[26] ),
    .B(_05279_),
    .X(_05346_));
 sky130_fd_sc_hd__a21oi_1 _12130_ (.A1(net26),
    .A2(_05346_),
    .B1(\div_res[27] ),
    .Y(_05347_));
 sky130_fd_sc_hd__a31o_1 _12131_ (.A1(\div_res[27] ),
    .A2(net26),
    .A3(_05346_),
    .B1(net203),
    .X(_05348_));
 sky130_fd_sc_hd__o21ai_1 _12132_ (.A1(_04915_),
    .A2(_02295_),
    .B1(_02291_),
    .Y(_05349_));
 sky130_fd_sc_hd__a221o_1 _12133_ (.A1(_04894_),
    .A2(net213),
    .B1(_02300_),
    .B2(_04915_),
    .C1(_06390_),
    .X(_05351_));
 sky130_fd_sc_hd__a21oi_1 _12134_ (.A1(_04937_),
    .A2(_05349_),
    .B1(_05351_),
    .Y(_05352_));
 sky130_fd_sc_hd__o221a_1 _12135_ (.A1(net186),
    .A2(_02944_),
    .B1(_02964_),
    .B2(net182),
    .C1(_05352_),
    .X(_05353_));
 sky130_fd_sc_hd__o211a_1 _12136_ (.A1(_05347_),
    .A2(_05348_),
    .B1(_05353_),
    .C1(_05345_),
    .X(_05354_));
 sky130_fd_sc_hd__o21ai_1 _12137_ (.A1(_06413_),
    .A2(_05342_),
    .B1(_05354_),
    .Y(_05355_));
 sky130_fd_sc_hd__a211o_1 _12138_ (.A1(net251),
    .A2(_05333_),
    .B1(_05335_),
    .C1(_05355_),
    .X(_05356_));
 sky130_fd_sc_hd__o22a_4 _12139_ (.A1(net261),
    .A2(_05294_),
    .B1(_05329_),
    .B2(_05356_),
    .X(dest_val[27]));
 sky130_fd_sc_hd__a2bb2o_1 _12140_ (.A1_N(net61),
    .A2_N(_05309_),
    .B1(_05310_),
    .B2(_05226_),
    .X(_05357_));
 sky130_fd_sc_hd__nor2_1 _12141_ (.A(net12),
    .B(net4),
    .Y(_05358_));
 sky130_fd_sc_hd__xnor2_1 _12142_ (.A(net98),
    .B(_05358_),
    .Y(_05359_));
 sky130_fd_sc_hd__o22a_1 _12143_ (.A1(net10),
    .A2(net7),
    .B1(net6),
    .B2(net16),
    .X(_05361_));
 sky130_fd_sc_hd__xnor2_1 _12144_ (.A(net30),
    .B(_05361_),
    .Y(_05362_));
 sky130_fd_sc_hd__a21o_1 _12145_ (.A1(_05298_),
    .A2(_05304_),
    .B1(_05362_),
    .X(_05363_));
 sky130_fd_sc_hd__nand3_1 _12146_ (.A(_05298_),
    .B(_05304_),
    .C(_05362_),
    .Y(_05364_));
 sky130_fd_sc_hd__nand2_1 _12147_ (.A(_05363_),
    .B(_05364_),
    .Y(_05365_));
 sky130_fd_sc_hd__or3_1 _12148_ (.A(net18),
    .B(net30),
    .C(_05365_),
    .X(_05366_));
 sky130_fd_sc_hd__o21ai_1 _12149_ (.A1(net18),
    .A2(net30),
    .B1(_05365_),
    .Y(_05367_));
 sky130_fd_sc_hd__nand2_1 _12150_ (.A(_05366_),
    .B(_05367_),
    .Y(_05368_));
 sky130_fd_sc_hd__or2_1 _12151_ (.A(_05359_),
    .B(_05368_),
    .X(_05369_));
 sky130_fd_sc_hd__nand2_1 _12152_ (.A(_05359_),
    .B(_05368_),
    .Y(_05370_));
 sky130_fd_sc_hd__nand2_1 _12153_ (.A(_05369_),
    .B(_05370_),
    .Y(_05372_));
 sky130_fd_sc_hd__nand2b_1 _12154_ (.A_N(_05372_),
    .B(_05357_),
    .Y(_05373_));
 sky130_fd_sc_hd__xor2_1 _12155_ (.A(_05357_),
    .B(_05372_),
    .X(_05374_));
 sky130_fd_sc_hd__o21ba_1 _12156_ (.A1(_05312_),
    .A2(_05315_),
    .B1_N(_05374_),
    .X(_05375_));
 sky130_fd_sc_hd__or3b_1 _12157_ (.A(_05312_),
    .B(_05315_),
    .C_N(_05374_),
    .X(_05376_));
 sky130_fd_sc_hd__and2b_1 _12158_ (.A_N(_05375_),
    .B(_05376_),
    .X(_05377_));
 sky130_fd_sc_hd__inv_2 _12159_ (.A(_05377_),
    .Y(_05378_));
 sky130_fd_sc_hd__nor2_1 _12160_ (.A(_05250_),
    .B(_05321_),
    .Y(_05379_));
 sky130_fd_sc_hd__inv_2 _12161_ (.A(_05379_),
    .Y(_05380_));
 sky130_fd_sc_hd__a2111o_1 _12162_ (.A1(_05064_),
    .A2(_05066_),
    .B1(_05105_),
    .C1(_05179_),
    .D1(_05380_),
    .X(_05381_));
 sky130_fd_sc_hd__a21boi_1 _12163_ (.A1(_05248_),
    .A2(_05319_),
    .B1_N(_05320_),
    .Y(_05383_));
 sky130_fd_sc_hd__o21ai_1 _12164_ (.A1(_05251_),
    .A2(_05380_),
    .B1(_05383_),
    .Y(_05384_));
 sky130_fd_sc_hd__inv_2 _12165_ (.A(_05384_),
    .Y(_05385_));
 sky130_fd_sc_hd__a21oi_1 _12166_ (.A1(_05381_),
    .A2(_05385_),
    .B1(_05378_),
    .Y(_05386_));
 sky130_fd_sc_hd__and3_1 _12167_ (.A(_05378_),
    .B(_05381_),
    .C(_05385_),
    .X(_05387_));
 sky130_fd_sc_hd__or2_1 _12168_ (.A(_05386_),
    .B(_05387_),
    .X(_05388_));
 sky130_fd_sc_hd__and2_1 _12169_ (.A(_05323_),
    .B(_05325_),
    .X(_05389_));
 sky130_fd_sc_hd__o21ai_1 _12170_ (.A1(net85),
    .A2(_05389_),
    .B1(_05388_),
    .Y(_05390_));
 sky130_fd_sc_hd__o31a_1 _12171_ (.A1(net85),
    .A2(_05388_),
    .A3(_05389_),
    .B1(net206),
    .X(_05391_));
 sky130_fd_sc_hd__a21o_1 _12172_ (.A1(_04937_),
    .A2(_05330_),
    .B1(_04915_),
    .X(_05392_));
 sky130_fd_sc_hd__and2_1 _12173_ (.A(net300),
    .B(_05392_),
    .X(_05394_));
 sky130_fd_sc_hd__a31o_1 _12174_ (.A1(net306),
    .A2(_06347_),
    .A3(_06361_),
    .B1(_05394_),
    .X(_05395_));
 sky130_fd_sc_hd__nand2_1 _12175_ (.A(_05306_),
    .B(_05395_),
    .Y(_05396_));
 sky130_fd_sc_hd__o211a_1 _12176_ (.A1(_05306_),
    .A2(_05395_),
    .B1(_05396_),
    .C1(net251),
    .X(_05397_));
 sky130_fd_sc_hd__a21oi_1 _12177_ (.A1(_02206_),
    .A2(_02208_),
    .B1(net86),
    .Y(_05398_));
 sky130_fd_sc_hd__xnor2_1 _12178_ (.A(_02139_),
    .B(_05398_),
    .Y(_05399_));
 sky130_fd_sc_hd__nor2_1 _12179_ (.A(net250),
    .B(_05399_),
    .Y(_05400_));
 sky130_fd_sc_hd__o21ai_2 _12180_ (.A1(_05336_),
    .A2(_05337_),
    .B1(_05338_),
    .Y(_05401_));
 sky130_fd_sc_hd__xor2_1 _12181_ (.A(reg1_val[28]),
    .B(_05401_),
    .X(_05402_));
 sky130_fd_sc_hd__nand2_1 _12182_ (.A(net242),
    .B(_02807_),
    .Y(_05403_));
 sky130_fd_sc_hd__o211a_1 _12183_ (.A1(net242),
    .A2(_05402_),
    .B1(_05403_),
    .C1(net215),
    .X(_05405_));
 sky130_fd_sc_hd__or2_1 _12184_ (.A(\div_shifter[59] ),
    .B(_05343_),
    .X(_05406_));
 sky130_fd_sc_hd__a21oi_1 _12185_ (.A1(net247),
    .A2(_05406_),
    .B1(\div_shifter[60] ),
    .Y(_05407_));
 sky130_fd_sc_hd__a31o_1 _12186_ (.A1(\div_shifter[60] ),
    .A2(net247),
    .A3(_05406_),
    .B1(net249),
    .X(_05408_));
 sky130_fd_sc_hd__nor2_1 _12187_ (.A(_05407_),
    .B(_05408_),
    .Y(_05409_));
 sky130_fd_sc_hd__or2_1 _12188_ (.A(\div_res[27] ),
    .B(_05346_),
    .X(_05410_));
 sky130_fd_sc_hd__a21o_1 _12189_ (.A1(net26),
    .A2(_05410_),
    .B1(\div_res[28] ),
    .X(_05411_));
 sky130_fd_sc_hd__nand3_1 _12190_ (.A(\div_res[28] ),
    .B(net26),
    .C(_05410_),
    .Y(_05412_));
 sky130_fd_sc_hd__o21ai_1 _12191_ (.A1(_05285_),
    .A2(_02295_),
    .B1(_02291_),
    .Y(_05413_));
 sky130_fd_sc_hd__a221o_1 _12192_ (.A1(_05285_),
    .A2(_02300_),
    .B1(_05413_),
    .B2(_05295_),
    .C1(net212),
    .X(_05414_));
 sky130_fd_sc_hd__a221o_1 _12193_ (.A1(_02217_),
    .A2(_02787_),
    .B1(_02808_),
    .B2(_02288_),
    .C1(_05414_),
    .X(_05416_));
 sky130_fd_sc_hd__a31o_1 _12194_ (.A1(_02305_),
    .A2(_05411_),
    .A3(_05412_),
    .B1(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__or4_1 _12195_ (.A(_05397_),
    .B(_05405_),
    .C(_05409_),
    .D(_05417_),
    .X(_05418_));
 sky130_fd_sc_hd__a211o_1 _12196_ (.A1(_05390_),
    .A2(_05391_),
    .B1(_05400_),
    .C1(_05418_),
    .X(_05419_));
 sky130_fd_sc_hd__o211a_4 _12197_ (.A1(_05263_),
    .A2(_06426_),
    .B1(_05419_),
    .C1(net261),
    .X(dest_val[28]));
 sky130_fd_sc_hd__o22a_1 _12198_ (.A1(net10),
    .A2(net5),
    .B1(net4),
    .B2(net7),
    .X(_05420_));
 sky130_fd_sc_hd__xnor2_1 _12199_ (.A(net30),
    .B(_05420_),
    .Y(_05421_));
 sky130_fd_sc_hd__a21o_1 _12200_ (.A1(_00228_),
    .A2(net33),
    .B1(net98),
    .X(_05422_));
 sky130_fd_sc_hd__or3b_1 _12201_ (.A(net16),
    .B(net30),
    .C_N(net98),
    .X(_05423_));
 sky130_fd_sc_hd__nand2_1 _12202_ (.A(_05422_),
    .B(_05423_),
    .Y(_05424_));
 sky130_fd_sc_hd__xor2_1 _12203_ (.A(_05421_),
    .B(_05424_),
    .X(_05426_));
 sky130_fd_sc_hd__nand2_1 _12204_ (.A(_05359_),
    .B(_05426_),
    .Y(_05427_));
 sky130_fd_sc_hd__or2_1 _12205_ (.A(_05359_),
    .B(_05426_),
    .X(_05428_));
 sky130_fd_sc_hd__nand2_1 _12206_ (.A(_05427_),
    .B(_05428_),
    .Y(_05429_));
 sky130_fd_sc_hd__a21o_1 _12207_ (.A1(_05363_),
    .A2(_05366_),
    .B1(_05429_),
    .X(_05430_));
 sky130_fd_sc_hd__nand3_1 _12208_ (.A(_05363_),
    .B(_05366_),
    .C(_05429_),
    .Y(_05431_));
 sky130_fd_sc_hd__nand2_1 _12209_ (.A(_05430_),
    .B(_05431_),
    .Y(_05432_));
 sky130_fd_sc_hd__a21o_1 _12210_ (.A1(_05369_),
    .A2(_05373_),
    .B1(_05432_),
    .X(_05433_));
 sky130_fd_sc_hd__nand3_1 _12211_ (.A(_05369_),
    .B(_05373_),
    .C(_05432_),
    .Y(_05434_));
 sky130_fd_sc_hd__and2_1 _12212_ (.A(_05433_),
    .B(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__o21ai_2 _12213_ (.A1(_05375_),
    .A2(_05386_),
    .B1(_05435_),
    .Y(_05437_));
 sky130_fd_sc_hd__or3_1 _12214_ (.A(_05375_),
    .B(_05386_),
    .C(_05435_),
    .X(_05438_));
 sky130_fd_sc_hd__nand2_1 _12215_ (.A(_05437_),
    .B(_05438_),
    .Y(_05439_));
 sky130_fd_sc_hd__a31o_1 _12216_ (.A1(_05323_),
    .A2(_05325_),
    .A3(_05388_),
    .B1(net85),
    .X(_05440_));
 sky130_fd_sc_hd__or2_1 _12217_ (.A(_05439_),
    .B(_05440_),
    .X(_05441_));
 sky130_fd_sc_hd__nand2_1 _12218_ (.A(_05439_),
    .B(_05440_),
    .Y(_05442_));
 sky130_fd_sc_hd__a21o_1 _12219_ (.A1(_05295_),
    .A2(_05392_),
    .B1(_05285_),
    .X(_05443_));
 sky130_fd_sc_hd__mux2_1 _12220_ (.A0(_06363_),
    .A1(_05443_),
    .S(net300),
    .X(_05444_));
 sky130_fd_sc_hd__nand2_1 _12221_ (.A(_05230_),
    .B(_05444_),
    .Y(_05445_));
 sky130_fd_sc_hd__o211a_1 _12222_ (.A1(_05230_),
    .A2(_05444_),
    .B1(_05445_),
    .C1(net251),
    .X(_05446_));
 sky130_fd_sc_hd__and3_1 _12223_ (.A(net27),
    .B(_02209_),
    .C(_02210_),
    .X(_05448_));
 sky130_fd_sc_hd__a21oi_1 _12224_ (.A1(net27),
    .A2(_02209_),
    .B1(_02210_),
    .Y(_05449_));
 sky130_fd_sc_hd__nor2_1 _12225_ (.A(_05448_),
    .B(_05449_),
    .Y(_05450_));
 sky130_fd_sc_hd__and3_1 _12226_ (.A(reg1_val[28]),
    .B(reg1_val[29]),
    .C(_05401_),
    .X(_05451_));
 sky130_fd_sc_hd__a21oi_1 _12227_ (.A1(reg1_val[28]),
    .A2(_05401_),
    .B1(reg1_val[29]),
    .Y(_05452_));
 sky130_fd_sc_hd__o21ai_1 _12228_ (.A1(_05451_),
    .A2(_05452_),
    .B1(net264),
    .Y(_05453_));
 sky130_fd_sc_hd__o211a_1 _12229_ (.A1(net264),
    .A2(_02625_),
    .B1(_05453_),
    .C1(net215),
    .X(_05454_));
 sky130_fd_sc_hd__nor2_1 _12230_ (.A(\div_shifter[60] ),
    .B(_05406_),
    .Y(_05455_));
 sky130_fd_sc_hd__o21a_1 _12231_ (.A1(\div_shifter[60] ),
    .A2(_05406_),
    .B1(net247),
    .X(_05456_));
 sky130_fd_sc_hd__o21ai_1 _12232_ (.A1(\div_shifter[61] ),
    .A2(_05456_),
    .B1(_02303_),
    .Y(_05457_));
 sky130_fd_sc_hd__a21oi_1 _12233_ (.A1(\div_shifter[61] ),
    .A2(_05456_),
    .B1(_05457_),
    .Y(_05459_));
 sky130_fd_sc_hd__o21a_1 _12234_ (.A1(\div_res[28] ),
    .A2(_05410_),
    .B1(net26),
    .X(_05460_));
 sky130_fd_sc_hd__o21ai_1 _12235_ (.A1(\div_res[29] ),
    .A2(_05460_),
    .B1(_02305_),
    .Y(_05461_));
 sky130_fd_sc_hd__a21o_1 _12236_ (.A1(\div_res[29] ),
    .A2(_05460_),
    .B1(_05461_),
    .X(_05462_));
 sky130_fd_sc_hd__o21ai_1 _12237_ (.A1(_05209_),
    .A2(_02295_),
    .B1(_02291_),
    .Y(_05463_));
 sky130_fd_sc_hd__a221o_1 _12238_ (.A1(_05209_),
    .A2(_02300_),
    .B1(_05463_),
    .B2(_05220_),
    .C1(net213),
    .X(_05464_));
 sky130_fd_sc_hd__a221o_1 _12239_ (.A1(_02288_),
    .A2(_02625_),
    .B1(_02639_),
    .B2(_02217_),
    .C1(_05464_),
    .X(_05465_));
 sky130_fd_sc_hd__or4b_1 _12240_ (.A(_05454_),
    .B(_05459_),
    .C(_05465_),
    .D_N(_05462_),
    .X(_05466_));
 sky130_fd_sc_hd__a211o_1 _12241_ (.A1(_02298_),
    .A2(_05450_),
    .B1(_05466_),
    .C1(_05446_),
    .X(_05467_));
 sky130_fd_sc_hd__a31o_1 _12242_ (.A1(net206),
    .A2(_05441_),
    .A3(_05442_),
    .B1(_05467_),
    .X(_05468_));
 sky130_fd_sc_hd__o211a_4 _12243_ (.A1(_05198_),
    .A2(_06426_),
    .B1(_05468_),
    .C1(net261),
    .X(dest_val[29]));
 sky130_fd_sc_hd__o21ai_1 _12244_ (.A1(_05421_),
    .A2(_05424_),
    .B1(_05423_),
    .Y(_05470_));
 sky130_fd_sc_hd__or3_1 _12245_ (.A(_00420_),
    .B(net30),
    .C(_00757_),
    .X(_05471_));
 sky130_fd_sc_hd__o21a_1 _12246_ (.A1(_00419_),
    .A2(_00757_),
    .B1(net30),
    .X(_05472_));
 sky130_fd_sc_hd__mux2_1 _12247_ (.A0(_00408_),
    .A1(_05472_),
    .S(_05471_),
    .X(_05473_));
 sky130_fd_sc_hd__and3b_1 _12248_ (.A_N(_00408_),
    .B(_00728_),
    .C(_05471_),
    .X(_05474_));
 sky130_fd_sc_hd__o21a_1 _12249_ (.A1(_05473_),
    .A2(_05474_),
    .B1(_05470_),
    .X(_05475_));
 sky130_fd_sc_hd__nor3_1 _12250_ (.A(_05470_),
    .B(_05473_),
    .C(_05474_),
    .Y(_05476_));
 sky130_fd_sc_hd__or2_1 _12251_ (.A(_05475_),
    .B(_05476_),
    .X(_05477_));
 sky130_fd_sc_hd__a21o_1 _12252_ (.A1(_05427_),
    .A2(_05430_),
    .B1(_05477_),
    .X(_05478_));
 sky130_fd_sc_hd__nand3_1 _12253_ (.A(_05427_),
    .B(_05430_),
    .C(_05477_),
    .Y(_05480_));
 sky130_fd_sc_hd__nand2_1 _12254_ (.A(_05478_),
    .B(_05480_),
    .Y(_05481_));
 sky130_fd_sc_hd__a21o_1 _12255_ (.A1(_05433_),
    .A2(_05437_),
    .B1(_05481_),
    .X(_05482_));
 sky130_fd_sc_hd__nand3_1 _12256_ (.A(_05433_),
    .B(_05437_),
    .C(_05481_),
    .Y(_05483_));
 sky130_fd_sc_hd__nand2_1 _12257_ (.A(_05482_),
    .B(_05483_),
    .Y(_05484_));
 sky130_fd_sc_hd__and4_1 _12258_ (.A(_05323_),
    .B(_05325_),
    .C(_05388_),
    .D(_05439_),
    .X(_05485_));
 sky130_fd_sc_hd__o21ai_1 _12259_ (.A1(net85),
    .A2(_05485_),
    .B1(_05484_),
    .Y(_05486_));
 sky130_fd_sc_hd__o31a_1 _12260_ (.A1(net85),
    .A2(_05484_),
    .A3(_05485_),
    .B1(net206),
    .X(_05487_));
 sky130_fd_sc_hd__and2_1 _12261_ (.A(_05486_),
    .B(_05487_),
    .X(_05488_));
 sky130_fd_sc_hd__a21o_1 _12262_ (.A1(_05220_),
    .A2(_05443_),
    .B1(_05209_),
    .X(_05489_));
 sky130_fd_sc_hd__mux2_1 _12263_ (.A0(_06365_),
    .A1(_05489_),
    .S(net300),
    .X(_05491_));
 sky130_fd_sc_hd__nand2_1 _12264_ (.A(_05078_),
    .B(_05491_),
    .Y(_05492_));
 sky130_fd_sc_hd__o211a_1 _12265_ (.A1(_05078_),
    .A2(_05491_),
    .B1(_05492_),
    .C1(net251),
    .X(_05493_));
 sky130_fd_sc_hd__o21ai_1 _12266_ (.A1(_02209_),
    .A2(_02210_),
    .B1(net27),
    .Y(_05494_));
 sky130_fd_sc_hd__xnor2_1 _12267_ (.A(_02138_),
    .B(_05494_),
    .Y(_05495_));
 sky130_fd_sc_hd__nand2_1 _12268_ (.A(reg1_val[30]),
    .B(_05451_),
    .Y(_05496_));
 sky130_fd_sc_hd__or2_1 _12269_ (.A(reg1_val[30]),
    .B(_05451_),
    .X(_05497_));
 sky130_fd_sc_hd__nand2_1 _12270_ (.A(_05496_),
    .B(_05497_),
    .Y(_05498_));
 sky130_fd_sc_hd__mux2_1 _12271_ (.A0(_02444_),
    .A1(_05498_),
    .S(net264),
    .X(_05499_));
 sky130_fd_sc_hd__nand2_1 _12272_ (.A(_04351_),
    .B(_05455_),
    .Y(_05500_));
 sky130_fd_sc_hd__a21oi_1 _12273_ (.A1(net247),
    .A2(_05500_),
    .B1(\div_shifter[62] ),
    .Y(_05502_));
 sky130_fd_sc_hd__a311o_1 _12274_ (.A1(\div_shifter[62] ),
    .A2(net247),
    .A3(_05500_),
    .B1(_05502_),
    .C1(net249),
    .X(_05503_));
 sky130_fd_sc_hd__or3_1 _12275_ (.A(\div_res[29] ),
    .B(\div_res[28] ),
    .C(_05410_),
    .X(_05504_));
 sky130_fd_sc_hd__a21oi_1 _12276_ (.A1(net26),
    .A2(_05504_),
    .B1(\div_res[30] ),
    .Y(_05505_));
 sky130_fd_sc_hd__a31o_1 _12277_ (.A1(\div_res[30] ),
    .A2(net26),
    .A3(_05504_),
    .B1(net203),
    .X(_05506_));
 sky130_fd_sc_hd__mux2_1 _12278_ (.A0(_02295_),
    .A1(_02301_),
    .S(_05057_),
    .X(_05507_));
 sky130_fd_sc_hd__a21oi_1 _12279_ (.A1(_02291_),
    .A2(_05507_),
    .B1(_05067_),
    .Y(_05508_));
 sky130_fd_sc_hd__nor2_1 _12280_ (.A(net212),
    .B(_05508_),
    .Y(_05509_));
 sky130_fd_sc_hd__o221a_1 _12281_ (.A1(net182),
    .A2(_02444_),
    .B1(_02476_),
    .B2(net186),
    .C1(_05509_),
    .X(_05510_));
 sky130_fd_sc_hd__o211a_1 _12282_ (.A1(_05505_),
    .A2(_05506_),
    .B1(_05510_),
    .C1(_05503_),
    .X(_05511_));
 sky130_fd_sc_hd__o21ai_1 _12283_ (.A1(net214),
    .A2(_05499_),
    .B1(_05511_),
    .Y(_05513_));
 sky130_fd_sc_hd__a211o_1 _12284_ (.A1(_02298_),
    .A2(_05495_),
    .B1(_05513_),
    .C1(_05493_),
    .X(_05514_));
 sky130_fd_sc_hd__o221a_4 _12285_ (.A1(_05046_),
    .A2(_06426_),
    .B1(_05488_),
    .B2(_05514_),
    .C1(net261),
    .X(dest_val[30]));
 sky130_fd_sc_hd__a21oi_1 _12286_ (.A1(_05484_),
    .A2(_05485_),
    .B1(net85),
    .Y(_05515_));
 sky130_fd_sc_hd__a21oi_1 _12287_ (.A1(net33),
    .A2(net4),
    .B1(_05473_),
    .Y(_05516_));
 sky130_fd_sc_hd__xnor2_2 _12288_ (.A(_05475_),
    .B(_05516_),
    .Y(_05517_));
 sky130_fd_sc_hd__and3_1 _12289_ (.A(_05478_),
    .B(_05482_),
    .C(_05517_),
    .X(_05518_));
 sky130_fd_sc_hd__nand3_1 _12290_ (.A(_05478_),
    .B(_05482_),
    .C(_05517_),
    .Y(_05519_));
 sky130_fd_sc_hd__a21oi_1 _12291_ (.A1(_05478_),
    .A2(_05482_),
    .B1(_05517_),
    .Y(_05520_));
 sky130_fd_sc_hd__a21o_1 _12292_ (.A1(_05478_),
    .A2(_05482_),
    .B1(_05517_),
    .X(_05521_));
 sky130_fd_sc_hd__a221o_1 _12293_ (.A1(_05484_),
    .A2(_05485_),
    .B1(_05519_),
    .B2(_05521_),
    .C1(net85),
    .X(_05523_));
 sky130_fd_sc_hd__o311a_1 _12294_ (.A1(_05515_),
    .A2(_05518_),
    .A3(_05520_),
    .B1(_05523_),
    .C1(net206),
    .X(_05524_));
 sky130_fd_sc_hd__a211oi_1 _12295_ (.A1(_05078_),
    .A2(_05489_),
    .B1(net306),
    .C1(_05057_),
    .Y(_05525_));
 sky130_fd_sc_hd__a21oi_1 _12296_ (.A1(net306),
    .A2(_06367_),
    .B1(_05525_),
    .Y(_05526_));
 sky130_fd_sc_hd__xnor2_1 _12297_ (.A(_04785_),
    .B(_05526_),
    .Y(_05527_));
 sky130_fd_sc_hd__o31a_1 _12298_ (.A1(_02138_),
    .A2(_02209_),
    .A3(_02210_),
    .B1(net27),
    .X(_05528_));
 sky130_fd_sc_hd__and2_1 _12299_ (.A(_02211_),
    .B(_05528_),
    .X(_05529_));
 sky130_fd_sc_hd__o21ai_1 _12300_ (.A1(_02211_),
    .A2(_05528_),
    .B1(_02298_),
    .Y(_05530_));
 sky130_fd_sc_hd__o21a_1 _12301_ (.A1(net242),
    .A2(_05496_),
    .B1(_02321_),
    .X(_05531_));
 sky130_fd_sc_hd__nor3_1 _12302_ (.A(net242),
    .B(_02321_),
    .C(_05496_),
    .Y(_05532_));
 sky130_fd_sc_hd__or3_1 _12303_ (.A(net214),
    .B(_05531_),
    .C(_05532_),
    .X(_05534_));
 sky130_fd_sc_hd__o21a_1 _12304_ (.A1(\div_shifter[62] ),
    .A2(_05500_),
    .B1(net247),
    .X(_05535_));
 sky130_fd_sc_hd__xnor2_1 _12305_ (.A(\div_shifter[63] ),
    .B(_05535_),
    .Y(_05536_));
 sky130_fd_sc_hd__o21a_1 _12306_ (.A1(\div_res[30] ),
    .A2(_05504_),
    .B1(net26),
    .X(_05537_));
 sky130_fd_sc_hd__o21ai_1 _12307_ (.A1(\div_res[31] ),
    .A2(_05537_),
    .B1(_02305_),
    .Y(_05538_));
 sky130_fd_sc_hd__a21o_1 _12308_ (.A1(\div_res[31] ),
    .A2(_05537_),
    .B1(_05538_),
    .X(_05539_));
 sky130_fd_sc_hd__o21a_1 _12309_ (.A1(reg1_val[31]),
    .A2(_04752_),
    .B1(net205),
    .X(_05540_));
 sky130_fd_sc_hd__a311o_1 _12310_ (.A1(reg1_val[31]),
    .A2(_04752_),
    .A3(_02300_),
    .B1(_05540_),
    .C1(net212),
    .X(_05541_));
 sky130_fd_sc_hd__a21oi_1 _12311_ (.A1(_04785_),
    .A2(_02294_),
    .B1(_05541_),
    .Y(_05542_));
 sky130_fd_sc_hd__o221a_1 _12312_ (.A1(net186),
    .A2(_02283_),
    .B1(net182),
    .B2(_02321_),
    .C1(_05542_),
    .X(_05543_));
 sky130_fd_sc_hd__o211a_1 _12313_ (.A1(net248),
    .A2(_05536_),
    .B1(_05539_),
    .C1(_05543_),
    .X(_05545_));
 sky130_fd_sc_hd__o211a_1 _12314_ (.A1(_05529_),
    .A2(_05530_),
    .B1(_05534_),
    .C1(_05545_),
    .X(_05546_));
 sky130_fd_sc_hd__o21ai_1 _12315_ (.A1(_02293_),
    .A2(_05527_),
    .B1(_05546_),
    .Y(_05547_));
 sky130_fd_sc_hd__o221a_4 _12316_ (.A1(_04752_),
    .A2(_06426_),
    .B1(_05524_),
    .B2(_05547_),
    .C1(net261),
    .X(dest_val[31]));
 sky130_fd_sc_hd__mux2_1 _12317_ (.A0(net304),
    .A1(curr_PC[0]),
    .S(net259),
    .X(_05548_));
 sky130_fd_sc_hd__nand2_1 _12318_ (.A(_04654_),
    .B(_05548_),
    .Y(_05549_));
 sky130_fd_sc_hd__or2_1 _12319_ (.A(_04654_),
    .B(_05548_),
    .X(_05550_));
 sky130_fd_sc_hd__and2_4 _12320_ (.A(_05549_),
    .B(_05550_),
    .X(new_PC[0]));
 sky130_fd_sc_hd__mux2_1 _12321_ (.A0(reg1_val[1]),
    .A1(curr_PC[1]),
    .S(net259),
    .X(_05551_));
 sky130_fd_sc_hd__nand2_1 _12322_ (.A(_05893_),
    .B(_05551_),
    .Y(_05552_));
 sky130_fd_sc_hd__or2_1 _12323_ (.A(_05893_),
    .B(_05551_),
    .X(_05554_));
 sky130_fd_sc_hd__nand2_1 _12324_ (.A(_05552_),
    .B(_05554_),
    .Y(_05555_));
 sky130_fd_sc_hd__or2_1 _12325_ (.A(_05549_),
    .B(_05555_),
    .X(_05556_));
 sky130_fd_sc_hd__nand2_1 _12326_ (.A(_05549_),
    .B(_05555_),
    .Y(_05557_));
 sky130_fd_sc_hd__and2_4 _12327_ (.A(_05556_),
    .B(_05557_),
    .X(new_PC[1]));
 sky130_fd_sc_hd__mux2_1 _12328_ (.A0(reg1_val[2]),
    .A1(curr_PC[2]),
    .S(net259),
    .X(_05558_));
 sky130_fd_sc_hd__nand2_1 _12329_ (.A(_05823_),
    .B(_05558_),
    .Y(_05559_));
 sky130_fd_sc_hd__or2_1 _12330_ (.A(_05823_),
    .B(_05558_),
    .X(_05560_));
 sky130_fd_sc_hd__nand2_1 _12331_ (.A(_05559_),
    .B(_05560_),
    .Y(_05561_));
 sky130_fd_sc_hd__a21o_1 _12332_ (.A1(_05552_),
    .A2(_05556_),
    .B1(_05561_),
    .X(_05562_));
 sky130_fd_sc_hd__nand3_1 _12333_ (.A(_05552_),
    .B(_05556_),
    .C(_05561_),
    .Y(_05564_));
 sky130_fd_sc_hd__and2_4 _12334_ (.A(_05562_),
    .B(_05564_),
    .X(new_PC[2]));
 sky130_fd_sc_hd__mux2_1 _12335_ (.A0(reg1_val[3]),
    .A1(curr_PC[3]),
    .S(net259),
    .X(_05565_));
 sky130_fd_sc_hd__nand2_1 _12336_ (.A(_05750_),
    .B(_05565_),
    .Y(_05566_));
 sky130_fd_sc_hd__or2_1 _12337_ (.A(_05750_),
    .B(_05565_),
    .X(_05567_));
 sky130_fd_sc_hd__nand2_1 _12338_ (.A(_05566_),
    .B(_05567_),
    .Y(_05568_));
 sky130_fd_sc_hd__a21o_1 _12339_ (.A1(_05559_),
    .A2(_05562_),
    .B1(_05568_),
    .X(_05569_));
 sky130_fd_sc_hd__nand3_1 _12340_ (.A(_05559_),
    .B(_05562_),
    .C(_05568_),
    .Y(_05570_));
 sky130_fd_sc_hd__and2_4 _12341_ (.A(_05569_),
    .B(_05570_),
    .X(new_PC[3]));
 sky130_fd_sc_hd__mux2_1 _12342_ (.A0(reg1_val[4]),
    .A1(curr_PC[4]),
    .S(net259),
    .X(_05571_));
 sky130_fd_sc_hd__nand2_1 _12343_ (.A(_05677_),
    .B(_05571_),
    .Y(_05573_));
 sky130_fd_sc_hd__or2_1 _12344_ (.A(_05677_),
    .B(_05571_),
    .X(_05574_));
 sky130_fd_sc_hd__nand2_1 _12345_ (.A(_05573_),
    .B(_05574_),
    .Y(_05575_));
 sky130_fd_sc_hd__a21o_1 _12346_ (.A1(_05566_),
    .A2(_05569_),
    .B1(_05575_),
    .X(_05576_));
 sky130_fd_sc_hd__nand3_1 _12347_ (.A(_05566_),
    .B(_05569_),
    .C(_05575_),
    .Y(_05577_));
 sky130_fd_sc_hd__and2_4 _12348_ (.A(_05576_),
    .B(_05577_),
    .X(new_PC[4]));
 sky130_fd_sc_hd__mux2_1 _12349_ (.A0(reg1_val[5]),
    .A1(curr_PC[5]),
    .S(net260),
    .X(_05578_));
 sky130_fd_sc_hd__nand2_1 _12350_ (.A(_05591_),
    .B(_05578_),
    .Y(_05579_));
 sky130_fd_sc_hd__or2_1 _12351_ (.A(_05591_),
    .B(_05578_),
    .X(_05580_));
 sky130_fd_sc_hd__nand2_1 _12352_ (.A(_05579_),
    .B(_05580_),
    .Y(_05581_));
 sky130_fd_sc_hd__a21o_1 _12353_ (.A1(_05573_),
    .A2(_05576_),
    .B1(_05581_),
    .X(_05583_));
 sky130_fd_sc_hd__nand3_1 _12354_ (.A(_05573_),
    .B(_05576_),
    .C(_05581_),
    .Y(_05584_));
 sky130_fd_sc_hd__and2_4 _12355_ (.A(_05583_),
    .B(_05584_),
    .X(new_PC[5]));
 sky130_fd_sc_hd__mux2_1 _12356_ (.A0(reg1_val[6]),
    .A1(curr_PC[6]),
    .S(net259),
    .X(_05585_));
 sky130_fd_sc_hd__nand2_1 _12357_ (.A(_05512_),
    .B(_05585_),
    .Y(_05586_));
 sky130_fd_sc_hd__or2_1 _12358_ (.A(_05512_),
    .B(_05585_),
    .X(_05587_));
 sky130_fd_sc_hd__nand2_1 _12359_ (.A(_05586_),
    .B(_05587_),
    .Y(_05588_));
 sky130_fd_sc_hd__a21o_1 _12360_ (.A1(_05579_),
    .A2(_05583_),
    .B1(_05588_),
    .X(_05589_));
 sky130_fd_sc_hd__nand3_1 _12361_ (.A(_05579_),
    .B(_05583_),
    .C(_05588_),
    .Y(_05590_));
 sky130_fd_sc_hd__and2_4 _12362_ (.A(_05589_),
    .B(_05590_),
    .X(new_PC[6]));
 sky130_fd_sc_hd__mux2_1 _12363_ (.A0(reg1_val[7]),
    .A1(curr_PC[7]),
    .S(net260),
    .X(_05592_));
 sky130_fd_sc_hd__nand2_1 _12364_ (.A(_05436_),
    .B(_05592_),
    .Y(_05593_));
 sky130_fd_sc_hd__or2_1 _12365_ (.A(_05436_),
    .B(_05592_),
    .X(_05594_));
 sky130_fd_sc_hd__nand2_1 _12366_ (.A(_05593_),
    .B(_05594_),
    .Y(_05595_));
 sky130_fd_sc_hd__a21o_1 _12367_ (.A1(_05586_),
    .A2(_05589_),
    .B1(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__nand3_1 _12368_ (.A(_05586_),
    .B(_05589_),
    .C(_05595_),
    .Y(_05597_));
 sky130_fd_sc_hd__and2_4 _12369_ (.A(_05596_),
    .B(_05597_),
    .X(new_PC[7]));
 sky130_fd_sc_hd__mux2_1 _12370_ (.A0(reg1_val[8]),
    .A1(curr_PC[8]),
    .S(net260),
    .X(_05598_));
 sky130_fd_sc_hd__nand2_1 _12371_ (.A(_05350_),
    .B(_05598_),
    .Y(_05599_));
 sky130_fd_sc_hd__or2_1 _12372_ (.A(_05350_),
    .B(_05598_),
    .X(_05600_));
 sky130_fd_sc_hd__nand2_1 _12373_ (.A(_05599_),
    .B(_05600_),
    .Y(_05602_));
 sky130_fd_sc_hd__a21o_1 _12374_ (.A1(_05593_),
    .A2(_05596_),
    .B1(_05602_),
    .X(_05603_));
 sky130_fd_sc_hd__nand3_1 _12375_ (.A(_05593_),
    .B(_05596_),
    .C(_05602_),
    .Y(_05604_));
 sky130_fd_sc_hd__and2_4 _12376_ (.A(_05603_),
    .B(_05604_),
    .X(new_PC[8]));
 sky130_fd_sc_hd__mux2_1 _12377_ (.A0(reg1_val[9]),
    .A1(curr_PC[9]),
    .S(net259),
    .X(_05605_));
 sky130_fd_sc_hd__nand2_1 _12378_ (.A(_05089_),
    .B(_05605_),
    .Y(_05606_));
 sky130_fd_sc_hd__or2_1 _12379_ (.A(_05089_),
    .B(_05605_),
    .X(_05607_));
 sky130_fd_sc_hd__nand2_1 _12380_ (.A(_05606_),
    .B(_05607_),
    .Y(_05608_));
 sky130_fd_sc_hd__a21o_1 _12381_ (.A1(_05599_),
    .A2(_05603_),
    .B1(_05608_),
    .X(_05609_));
 sky130_fd_sc_hd__nand3_1 _12382_ (.A(_05599_),
    .B(_05603_),
    .C(_05608_),
    .Y(_05610_));
 sky130_fd_sc_hd__and2_4 _12383_ (.A(_05609_),
    .B(_05610_),
    .X(new_PC[9]));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(reg1_val[10]),
    .A1(curr_PC[10]),
    .S(net260),
    .X(_05612_));
 sky130_fd_sc_hd__nand2_1 _12385_ (.A(_04959_),
    .B(_05612_),
    .Y(_05613_));
 sky130_fd_sc_hd__or2_1 _12386_ (.A(_04959_),
    .B(_05612_),
    .X(_05614_));
 sky130_fd_sc_hd__nand2_1 _12387_ (.A(_05613_),
    .B(_05614_),
    .Y(_05615_));
 sky130_fd_sc_hd__a21o_1 _12388_ (.A1(_05606_),
    .A2(_05609_),
    .B1(_05615_),
    .X(_05616_));
 sky130_fd_sc_hd__nand3_1 _12389_ (.A(_05606_),
    .B(_05609_),
    .C(_05615_),
    .Y(_05617_));
 sky130_fd_sc_hd__and2_4 _12390_ (.A(_05616_),
    .B(_05617_),
    .X(new_PC[10]));
 sky130_fd_sc_hd__mux2_1 _12391_ (.A0(reg1_val[11]),
    .A1(curr_PC[11]),
    .S(net259),
    .X(_05618_));
 sky130_fd_sc_hd__nand2_1 _12392_ (.A(_04807_),
    .B(_05618_),
    .Y(_05619_));
 sky130_fd_sc_hd__or2_1 _12393_ (.A(_04807_),
    .B(_05618_),
    .X(_05621_));
 sky130_fd_sc_hd__nand2_1 _12394_ (.A(_05619_),
    .B(_05621_),
    .Y(_05622_));
 sky130_fd_sc_hd__a21o_1 _12395_ (.A1(_05613_),
    .A2(_05616_),
    .B1(_05622_),
    .X(_05623_));
 sky130_fd_sc_hd__nand3_1 _12396_ (.A(_05613_),
    .B(_05616_),
    .C(_05622_),
    .Y(_05624_));
 sky130_fd_sc_hd__and2_4 _12397_ (.A(_05623_),
    .B(_05624_),
    .X(new_PC[11]));
 sky130_fd_sc_hd__mux2_1 _12398_ (.A0(reg1_val[12]),
    .A1(curr_PC[12]),
    .S(net259),
    .X(_05625_));
 sky130_fd_sc_hd__nand2_1 _12399_ (.A(_04872_),
    .B(_05625_),
    .Y(_05626_));
 sky130_fd_sc_hd__or2_1 _12400_ (.A(_04872_),
    .B(_05625_),
    .X(_05627_));
 sky130_fd_sc_hd__nand2_1 _12401_ (.A(_05626_),
    .B(_05627_),
    .Y(_05628_));
 sky130_fd_sc_hd__a21o_1 _12402_ (.A1(_05619_),
    .A2(_05623_),
    .B1(_05628_),
    .X(_05629_));
 sky130_fd_sc_hd__nand3_1 _12403_ (.A(_05619_),
    .B(_05623_),
    .C(_05628_),
    .Y(_05631_));
 sky130_fd_sc_hd__and2_4 _12404_ (.A(_05629_),
    .B(_05631_),
    .X(new_PC[12]));
 sky130_fd_sc_hd__mux2_1 _12405_ (.A0(net303),
    .A1(curr_PC[13]),
    .S(net259),
    .X(_05632_));
 sky130_fd_sc_hd__nand2_1 _12406_ (.A(_05241_),
    .B(_05632_),
    .Y(_05633_));
 sky130_fd_sc_hd__or2_1 _12407_ (.A(_05241_),
    .B(_05632_),
    .X(_05634_));
 sky130_fd_sc_hd__nand2_1 _12408_ (.A(_05633_),
    .B(_05634_),
    .Y(_05635_));
 sky130_fd_sc_hd__a21o_1 _12409_ (.A1(_05626_),
    .A2(_05629_),
    .B1(_05635_),
    .X(_05636_));
 sky130_fd_sc_hd__nand3_1 _12410_ (.A(_05626_),
    .B(_05629_),
    .C(_05635_),
    .Y(_05637_));
 sky130_fd_sc_hd__and2_4 _12411_ (.A(_05636_),
    .B(_05637_),
    .X(new_PC[13]));
 sky130_fd_sc_hd__mux2_1 _12412_ (.A0(reg1_val[14]),
    .A1(curr_PC[14]),
    .S(net259),
    .X(_05638_));
 sky130_fd_sc_hd__nand2_1 _12413_ (.A(_05165_),
    .B(_05638_),
    .Y(_05640_));
 sky130_fd_sc_hd__or2_1 _12414_ (.A(_05165_),
    .B(_05638_),
    .X(_05641_));
 sky130_fd_sc_hd__nand2_1 _12415_ (.A(_05640_),
    .B(_05641_),
    .Y(_05642_));
 sky130_fd_sc_hd__a21o_1 _12416_ (.A1(_05633_),
    .A2(_05636_),
    .B1(_05642_),
    .X(_05643_));
 sky130_fd_sc_hd__nand3_1 _12417_ (.A(_05633_),
    .B(_05636_),
    .C(_05642_),
    .Y(_05644_));
 sky130_fd_sc_hd__and2_4 _12418_ (.A(_05643_),
    .B(_05644_),
    .X(new_PC[14]));
 sky130_fd_sc_hd__mux2_1 _12419_ (.A0(reg1_val[15]),
    .A1(curr_PC[15]),
    .S(net259),
    .X(_05645_));
 sky130_fd_sc_hd__nand2_1 _12420_ (.A(_05024_),
    .B(_05645_),
    .Y(_05646_));
 sky130_fd_sc_hd__or2_1 _12421_ (.A(_05024_),
    .B(_05645_),
    .X(_05647_));
 sky130_fd_sc_hd__nand2_1 _12422_ (.A(_05646_),
    .B(_05647_),
    .Y(_05648_));
 sky130_fd_sc_hd__a21o_1 _12423_ (.A1(_05640_),
    .A2(_05643_),
    .B1(_05648_),
    .X(_05650_));
 sky130_fd_sc_hd__nand3_1 _12424_ (.A(_05640_),
    .B(_05643_),
    .C(_05648_),
    .Y(_05651_));
 sky130_fd_sc_hd__and2_4 _12425_ (.A(_05650_),
    .B(_05651_),
    .X(new_PC[15]));
 sky130_fd_sc_hd__mux2_2 _12426_ (.A0(reg1_val[16]),
    .A1(curr_PC[16]),
    .S(net259),
    .X(_05652_));
 sky130_fd_sc_hd__xnor2_1 _12427_ (.A(net277),
    .B(_05652_),
    .Y(_05653_));
 sky130_fd_sc_hd__a21o_1 _12428_ (.A1(_05646_),
    .A2(_05650_),
    .B1(_05653_),
    .X(_05654_));
 sky130_fd_sc_hd__nand3_1 _12429_ (.A(_05646_),
    .B(_05650_),
    .C(_05653_),
    .Y(_05655_));
 sky130_fd_sc_hd__and2_4 _12430_ (.A(_05654_),
    .B(_05655_),
    .X(new_PC[16]));
 sky130_fd_sc_hd__mux2_2 _12431_ (.A0(reg1_val[17]),
    .A1(curr_PC[17]),
    .S(net259),
    .X(_05656_));
 sky130_fd_sc_hd__xnor2_4 _12432_ (.A(net276),
    .B(_05656_),
    .Y(_05657_));
 sky130_fd_sc_hd__a21bo_1 _12433_ (.A1(net276),
    .A2(_05652_),
    .B1_N(_05654_),
    .X(_05659_));
 sky130_fd_sc_hd__xnor2_4 _12434_ (.A(_05657_),
    .B(_05659_),
    .Y(new_PC[17]));
 sky130_fd_sc_hd__mux2_1 _12435_ (.A0(reg1_val[18]),
    .A1(curr_PC[18]),
    .S(net259),
    .X(_05660_));
 sky130_fd_sc_hd__nand2_1 _12436_ (.A(net276),
    .B(_05660_),
    .Y(_05661_));
 sky130_fd_sc_hd__or2_1 _12437_ (.A(net276),
    .B(_05660_),
    .X(_05662_));
 sky130_fd_sc_hd__nand2_1 _12438_ (.A(_05661_),
    .B(_05662_),
    .Y(_05663_));
 sky130_fd_sc_hd__or2_1 _12439_ (.A(_05654_),
    .B(_05657_),
    .X(_05664_));
 sky130_fd_sc_hd__o21ai_1 _12440_ (.A1(_05652_),
    .A2(_05656_),
    .B1(net276),
    .Y(_05665_));
 sky130_fd_sc_hd__a21o_1 _12441_ (.A1(_05664_),
    .A2(_05665_),
    .B1(_05663_),
    .X(_05666_));
 sky130_fd_sc_hd__nand3_1 _12442_ (.A(_05663_),
    .B(_05664_),
    .C(_05665_),
    .Y(_05667_));
 sky130_fd_sc_hd__and2_4 _12443_ (.A(_05666_),
    .B(_05667_),
    .X(new_PC[18]));
 sky130_fd_sc_hd__mux2_1 _12444_ (.A0(reg1_val[19]),
    .A1(curr_PC[19]),
    .S(net259),
    .X(_05669_));
 sky130_fd_sc_hd__nand2_1 _12445_ (.A(net276),
    .B(_05669_),
    .Y(_05670_));
 sky130_fd_sc_hd__or2_1 _12446_ (.A(net276),
    .B(_05669_),
    .X(_05671_));
 sky130_fd_sc_hd__nand2_2 _12447_ (.A(_05670_),
    .B(_05671_),
    .Y(_05672_));
 sky130_fd_sc_hd__nand2_2 _12448_ (.A(_05661_),
    .B(_05666_),
    .Y(_05673_));
 sky130_fd_sc_hd__xnor2_4 _12449_ (.A(_05672_),
    .B(_05673_),
    .Y(new_PC[19]));
 sky130_fd_sc_hd__mux2_2 _12450_ (.A0(reg1_val[20]),
    .A1(curr_PC[20]),
    .S(net260),
    .X(_05674_));
 sky130_fd_sc_hd__nand2_1 _12451_ (.A(net276),
    .B(_05674_),
    .Y(_05675_));
 sky130_fd_sc_hd__or2_1 _12452_ (.A(net276),
    .B(_05674_),
    .X(_05676_));
 sky130_fd_sc_hd__nand2_2 _12453_ (.A(_05675_),
    .B(_05676_),
    .Y(_05678_));
 sky130_fd_sc_hd__or3_1 _12454_ (.A(_05663_),
    .B(_05664_),
    .C(_05672_),
    .X(_05679_));
 sky130_fd_sc_hd__and3_1 _12455_ (.A(_05661_),
    .B(_05665_),
    .C(_05670_),
    .X(_05680_));
 sky130_fd_sc_hd__nand2_2 _12456_ (.A(_05679_),
    .B(_05680_),
    .Y(_05681_));
 sky130_fd_sc_hd__inv_2 _12457_ (.A(_05681_),
    .Y(_05682_));
 sky130_fd_sc_hd__xnor2_4 _12458_ (.A(_05678_),
    .B(_05681_),
    .Y(new_PC[20]));
 sky130_fd_sc_hd__mux2_2 _12459_ (.A0(reg1_val[21]),
    .A1(curr_PC[21]),
    .S(net260),
    .X(_05683_));
 sky130_fd_sc_hd__xnor2_4 _12460_ (.A(net276),
    .B(_05683_),
    .Y(_05684_));
 sky130_fd_sc_hd__o21ai_2 _12461_ (.A1(_05678_),
    .A2(_05682_),
    .B1(_05675_),
    .Y(_05685_));
 sky130_fd_sc_hd__xnor2_4 _12462_ (.A(_05684_),
    .B(_05685_),
    .Y(new_PC[21]));
 sky130_fd_sc_hd__mux2_1 _12463_ (.A0(reg1_val[22]),
    .A1(curr_PC[22]),
    .S(net260),
    .X(_05687_));
 sky130_fd_sc_hd__and2_1 _12464_ (.A(net276),
    .B(_05687_),
    .X(_05688_));
 sky130_fd_sc_hd__or2_1 _12465_ (.A(net276),
    .B(_05687_),
    .X(_05689_));
 sky130_fd_sc_hd__nand2b_2 _12466_ (.A_N(_05688_),
    .B(_05689_),
    .Y(_05690_));
 sky130_fd_sc_hd__o21ai_2 _12467_ (.A1(_05674_),
    .A2(_05683_),
    .B1(net277),
    .Y(_05691_));
 sky130_fd_sc_hd__nor2_1 _12468_ (.A(_05678_),
    .B(_05684_),
    .Y(_05692_));
 sky130_fd_sc_hd__inv_2 _12469_ (.A(_05692_),
    .Y(_05693_));
 sky130_fd_sc_hd__o21ai_4 _12470_ (.A1(_05682_),
    .A2(_05693_),
    .B1(_05691_),
    .Y(_05694_));
 sky130_fd_sc_hd__xnor2_4 _12471_ (.A(_05690_),
    .B(_05694_),
    .Y(new_PC[22]));
 sky130_fd_sc_hd__mux2_2 _12472_ (.A0(reg1_val[23]),
    .A1(curr_PC[23]),
    .S(net260),
    .X(_05695_));
 sky130_fd_sc_hd__xnor2_4 _12473_ (.A(net276),
    .B(_05695_),
    .Y(_05697_));
 sky130_fd_sc_hd__a21o_1 _12474_ (.A1(_05689_),
    .A2(_05694_),
    .B1(_05688_),
    .X(_05698_));
 sky130_fd_sc_hd__xnor2_4 _12475_ (.A(_05697_),
    .B(_05698_),
    .Y(new_PC[23]));
 sky130_fd_sc_hd__mux2_2 _12476_ (.A0(reg1_val[24]),
    .A1(curr_PC[24]),
    .S(net260),
    .X(_05699_));
 sky130_fd_sc_hd__xnor2_4 _12477_ (.A(net277),
    .B(_05699_),
    .Y(_05700_));
 sky130_fd_sc_hd__or4_1 _12478_ (.A(_05679_),
    .B(_05690_),
    .C(_05693_),
    .D(_05697_),
    .X(_05701_));
 sky130_fd_sc_hd__o21ai_1 _12479_ (.A1(_05687_),
    .A2(_05695_),
    .B1(net277),
    .Y(_05702_));
 sky130_fd_sc_hd__and4_2 _12480_ (.A(_05680_),
    .B(_05691_),
    .C(_05701_),
    .D(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__xor2_4 _12481_ (.A(_05700_),
    .B(_05703_),
    .X(new_PC[24]));
 sky130_fd_sc_hd__mux2_1 _12482_ (.A0(reg1_val[25]),
    .A1(curr_PC[25]),
    .S(net260),
    .X(_05704_));
 sky130_fd_sc_hd__and2_1 _12483_ (.A(net277),
    .B(_05704_),
    .X(_05706_));
 sky130_fd_sc_hd__nor2_1 _12484_ (.A(net277),
    .B(_05704_),
    .Y(_05707_));
 sky130_fd_sc_hd__nor2_2 _12485_ (.A(_05706_),
    .B(_05707_),
    .Y(_05708_));
 sky130_fd_sc_hd__o2bb2a_2 _12486_ (.A1_N(net277),
    .A2_N(_05699_),
    .B1(_05700_),
    .B2(_05703_),
    .X(_05709_));
 sky130_fd_sc_hd__xnor2_4 _12487_ (.A(_05708_),
    .B(_05709_),
    .Y(new_PC[25]));
 sky130_fd_sc_hd__mux2_1 _12488_ (.A0(reg1_val[26]),
    .A1(curr_PC[26]),
    .S(net260),
    .X(_05710_));
 sky130_fd_sc_hd__and2_1 _12489_ (.A(net276),
    .B(_05710_),
    .X(_05711_));
 sky130_fd_sc_hd__nor2_1 _12490_ (.A(net276),
    .B(_05710_),
    .Y(_05712_));
 sky130_fd_sc_hd__nor2_2 _12491_ (.A(_05711_),
    .B(_05712_),
    .Y(_05713_));
 sky130_fd_sc_hd__o21ba_2 _12492_ (.A1(_05707_),
    .A2(_05709_),
    .B1_N(_05706_),
    .X(_05714_));
 sky130_fd_sc_hd__xnor2_4 _12493_ (.A(_05713_),
    .B(_05714_),
    .Y(new_PC[26]));
 sky130_fd_sc_hd__o21ba_1 _12494_ (.A1(_05712_),
    .A2(_05714_),
    .B1_N(_05711_),
    .X(_05716_));
 sky130_fd_sc_hd__mux2_1 _12495_ (.A0(reg1_val[27]),
    .A1(curr_PC[27]),
    .S(net260),
    .X(_05717_));
 sky130_fd_sc_hd__xor2_2 _12496_ (.A(net276),
    .B(_05717_),
    .X(_05718_));
 sky130_fd_sc_hd__xnor2_4 _12497_ (.A(_05716_),
    .B(_05718_),
    .Y(new_PC[27]));
 sky130_fd_sc_hd__and3_4 _12498_ (.A(reg1_val[0]),
    .B(instruction[25]),
    .C(net282),
    .X(_05719_));
 sky130_fd_sc_hd__nor2_2 _12499_ (.A(net304),
    .B(_04654_),
    .Y(_05720_));
 sky130_fd_sc_hd__nor2_8 _12500_ (.A(_05719_),
    .B(_05720_),
    .Y(loadstore_address[0]));
 sky130_fd_sc_hd__nor2_1 _12501_ (.A(_04438_),
    .B(_05899_),
    .Y(_05721_));
 sky130_fd_sc_hd__or2_2 _12502_ (.A(reg1_val[1]),
    .B(_05893_),
    .X(_05722_));
 sky130_fd_sc_hd__nand2b_2 _12503_ (.A_N(_05721_),
    .B(_05722_),
    .Y(_05724_));
 sky130_fd_sc_hd__xnor2_4 _12504_ (.A(_05719_),
    .B(_05724_),
    .Y(loadstore_address[1]));
 sky130_fd_sc_hd__a21oi_4 _12505_ (.A1(_05719_),
    .A2(_05722_),
    .B1(_05721_),
    .Y(_05725_));
 sky130_fd_sc_hd__nor2_1 _12506_ (.A(reg1_val[2]),
    .B(_05823_),
    .Y(_05726_));
 sky130_fd_sc_hd__nand2_1 _12507_ (.A(reg1_val[2]),
    .B(_05823_),
    .Y(_05727_));
 sky130_fd_sc_hd__nand2b_2 _12508_ (.A_N(_05726_),
    .B(_05727_),
    .Y(_05728_));
 sky130_fd_sc_hd__xor2_4 _12509_ (.A(_05725_),
    .B(_05728_),
    .X(loadstore_address[2]));
 sky130_fd_sc_hd__o21a_2 _12510_ (.A1(_05725_),
    .A2(_05726_),
    .B1(_05727_),
    .X(_05729_));
 sky130_fd_sc_hd__nor2_1 _12511_ (.A(reg1_val[3]),
    .B(_05750_),
    .Y(_05730_));
 sky130_fd_sc_hd__nand2_1 _12512_ (.A(reg1_val[3]),
    .B(_05750_),
    .Y(_05731_));
 sky130_fd_sc_hd__nand2b_2 _12513_ (.A_N(_05730_),
    .B(_05731_),
    .Y(_05733_));
 sky130_fd_sc_hd__xor2_4 _12514_ (.A(_05729_),
    .B(_05733_),
    .X(loadstore_address[3]));
 sky130_fd_sc_hd__o21a_2 _12515_ (.A1(_05729_),
    .A2(_05730_),
    .B1(_05731_),
    .X(_05734_));
 sky130_fd_sc_hd__nor2_1 _12516_ (.A(reg1_val[4]),
    .B(_05677_),
    .Y(_05735_));
 sky130_fd_sc_hd__nand2_1 _12517_ (.A(reg1_val[4]),
    .B(_05677_),
    .Y(_05736_));
 sky130_fd_sc_hd__nand2b_2 _12518_ (.A_N(_05735_),
    .B(_05736_),
    .Y(_05737_));
 sky130_fd_sc_hd__xor2_4 _12519_ (.A(_05734_),
    .B(_05737_),
    .X(loadstore_address[4]));
 sky130_fd_sc_hd__o21a_2 _12520_ (.A1(_05734_),
    .A2(_05735_),
    .B1(_05736_),
    .X(_05738_));
 sky130_fd_sc_hd__nor2_1 _12521_ (.A(reg1_val[5]),
    .B(_05591_),
    .Y(_05739_));
 sky130_fd_sc_hd__nand2_1 _12522_ (.A(reg1_val[5]),
    .B(_05591_),
    .Y(_05740_));
 sky130_fd_sc_hd__nand2b_2 _12523_ (.A_N(_05739_),
    .B(_05740_),
    .Y(_05742_));
 sky130_fd_sc_hd__xor2_4 _12524_ (.A(_05738_),
    .B(_05742_),
    .X(loadstore_address[5]));
 sky130_fd_sc_hd__o21a_2 _12525_ (.A1(_05738_),
    .A2(_05739_),
    .B1(_05740_),
    .X(_05743_));
 sky130_fd_sc_hd__nor2_1 _12526_ (.A(reg1_val[6]),
    .B(_05512_),
    .Y(_05744_));
 sky130_fd_sc_hd__nand2_1 _12527_ (.A(reg1_val[6]),
    .B(_05512_),
    .Y(_05745_));
 sky130_fd_sc_hd__and2b_1 _12528_ (.A_N(_05744_),
    .B(_05745_),
    .X(_05746_));
 sky130_fd_sc_hd__xnor2_4 _12529_ (.A(_05743_),
    .B(_05746_),
    .Y(loadstore_address[6]));
 sky130_fd_sc_hd__o21a_2 _12530_ (.A1(_05743_),
    .A2(_05744_),
    .B1(_05745_),
    .X(_05747_));
 sky130_fd_sc_hd__nor2_1 _12531_ (.A(reg1_val[7]),
    .B(_05436_),
    .Y(_05748_));
 sky130_fd_sc_hd__nand2_1 _12532_ (.A(reg1_val[7]),
    .B(_05436_),
    .Y(_05749_));
 sky130_fd_sc_hd__nand2b_2 _12533_ (.A_N(_05748_),
    .B(_05749_),
    .Y(_05751_));
 sky130_fd_sc_hd__xor2_4 _12534_ (.A(_05747_),
    .B(_05751_),
    .X(loadstore_address[7]));
 sky130_fd_sc_hd__o21a_2 _12535_ (.A1(_05747_),
    .A2(_05748_),
    .B1(_05749_),
    .X(_05752_));
 sky130_fd_sc_hd__nor2_1 _12536_ (.A(reg1_val[8]),
    .B(_05350_),
    .Y(_05753_));
 sky130_fd_sc_hd__nand2_1 _12537_ (.A(reg1_val[8]),
    .B(_05350_),
    .Y(_05754_));
 sky130_fd_sc_hd__nand2b_2 _12538_ (.A_N(_05753_),
    .B(_05754_),
    .Y(_05755_));
 sky130_fd_sc_hd__xor2_4 _12539_ (.A(_05752_),
    .B(_05755_),
    .X(loadstore_address[8]));
 sky130_fd_sc_hd__o21a_2 _12540_ (.A1(_05752_),
    .A2(_05753_),
    .B1(_05754_),
    .X(_05756_));
 sky130_fd_sc_hd__or2_1 _12541_ (.A(reg1_val[9]),
    .B(_05089_),
    .X(_05757_));
 sky130_fd_sc_hd__nand2_1 _12542_ (.A(reg1_val[9]),
    .B(_05089_),
    .Y(_05758_));
 sky130_fd_sc_hd__nand2_2 _12543_ (.A(_05757_),
    .B(_05758_),
    .Y(_05760_));
 sky130_fd_sc_hd__xor2_4 _12544_ (.A(_05756_),
    .B(_05760_),
    .X(loadstore_address[9]));
 sky130_fd_sc_hd__or2_1 _12545_ (.A(reg1_val[10]),
    .B(_04959_),
    .X(_05761_));
 sky130_fd_sc_hd__nand2_1 _12546_ (.A(reg1_val[10]),
    .B(_04959_),
    .Y(_05762_));
 sky130_fd_sc_hd__nand2_1 _12547_ (.A(_05761_),
    .B(_05762_),
    .Y(_05763_));
 sky130_fd_sc_hd__nand2b_1 _12548_ (.A_N(_05756_),
    .B(_05757_),
    .Y(_05764_));
 sky130_fd_sc_hd__a21o_1 _12549_ (.A1(_05758_),
    .A2(_05764_),
    .B1(_05763_),
    .X(_05765_));
 sky130_fd_sc_hd__nand3_1 _12550_ (.A(_05758_),
    .B(_05763_),
    .C(_05764_),
    .Y(_05766_));
 sky130_fd_sc_hd__and2_4 _12551_ (.A(_05765_),
    .B(_05766_),
    .X(loadstore_address[10]));
 sky130_fd_sc_hd__or2_1 _12552_ (.A(reg1_val[11]),
    .B(_04807_),
    .X(_05767_));
 sky130_fd_sc_hd__nand2_1 _12553_ (.A(reg1_val[11]),
    .B(_04807_),
    .Y(_05769_));
 sky130_fd_sc_hd__nand2_1 _12554_ (.A(_05767_),
    .B(_05769_),
    .Y(_05770_));
 sky130_fd_sc_hd__a21o_1 _12555_ (.A1(_05762_),
    .A2(_05765_),
    .B1(_05770_),
    .X(_05771_));
 sky130_fd_sc_hd__nand3_1 _12556_ (.A(_05762_),
    .B(_05765_),
    .C(_05770_),
    .Y(_05772_));
 sky130_fd_sc_hd__and2_4 _12557_ (.A(_05771_),
    .B(_05772_),
    .X(loadstore_address[11]));
 sky130_fd_sc_hd__or2_1 _12558_ (.A(reg1_val[12]),
    .B(_04872_),
    .X(_05773_));
 sky130_fd_sc_hd__nand2_1 _12559_ (.A(reg1_val[12]),
    .B(_04872_),
    .Y(_05774_));
 sky130_fd_sc_hd__nand2_1 _12560_ (.A(_05773_),
    .B(_05774_),
    .Y(_05775_));
 sky130_fd_sc_hd__a21o_1 _12561_ (.A1(_05769_),
    .A2(_05771_),
    .B1(_05775_),
    .X(_05776_));
 sky130_fd_sc_hd__nand3_1 _12562_ (.A(_05769_),
    .B(_05771_),
    .C(_05775_),
    .Y(_05777_));
 sky130_fd_sc_hd__and2_4 _12563_ (.A(_05776_),
    .B(_05777_),
    .X(loadstore_address[12]));
 sky130_fd_sc_hd__or2_1 _12564_ (.A(reg1_val[13]),
    .B(_05241_),
    .X(_05779_));
 sky130_fd_sc_hd__nand2_1 _12565_ (.A(reg1_val[13]),
    .B(_05241_),
    .Y(_05780_));
 sky130_fd_sc_hd__nand2_1 _12566_ (.A(_05779_),
    .B(_05780_),
    .Y(_05781_));
 sky130_fd_sc_hd__a21o_1 _12567_ (.A1(_05774_),
    .A2(_05776_),
    .B1(_05781_),
    .X(_05782_));
 sky130_fd_sc_hd__nand3_1 _12568_ (.A(_05774_),
    .B(_05776_),
    .C(_05781_),
    .Y(_05783_));
 sky130_fd_sc_hd__and2_4 _12569_ (.A(_05782_),
    .B(_05783_),
    .X(loadstore_address[13]));
 sky130_fd_sc_hd__or2_1 _12570_ (.A(reg1_val[14]),
    .B(_05165_),
    .X(_05784_));
 sky130_fd_sc_hd__nand2_1 _12571_ (.A(reg1_val[14]),
    .B(_05165_),
    .Y(_05785_));
 sky130_fd_sc_hd__nand2_1 _12572_ (.A(_05784_),
    .B(_05785_),
    .Y(_05786_));
 sky130_fd_sc_hd__a21o_1 _12573_ (.A1(_05780_),
    .A2(_05782_),
    .B1(_05786_),
    .X(_05788_));
 sky130_fd_sc_hd__nand3_1 _12574_ (.A(_05780_),
    .B(_05782_),
    .C(_05786_),
    .Y(_05789_));
 sky130_fd_sc_hd__and2_4 _12575_ (.A(_05788_),
    .B(_05789_),
    .X(loadstore_address[14]));
 sky130_fd_sc_hd__xnor2_2 _12576_ (.A(reg1_val[15]),
    .B(_05024_),
    .Y(_05790_));
 sky130_fd_sc_hd__a21oi_4 _12577_ (.A1(_05785_),
    .A2(_05788_),
    .B1(_05790_),
    .Y(_05791_));
 sky130_fd_sc_hd__and3_2 _12578_ (.A(_05785_),
    .B(_05788_),
    .C(_05790_),
    .X(_05792_));
 sky130_fd_sc_hd__nor2_8 _12579_ (.A(_05791_),
    .B(_05792_),
    .Y(loadstore_address[15]));
 sky130_fd_sc_hd__nor2_1 _12580_ (.A(reg1_val[16]),
    .B(net278),
    .Y(_05793_));
 sky130_fd_sc_hd__and2_1 _12581_ (.A(reg1_val[16]),
    .B(net278),
    .X(_05794_));
 sky130_fd_sc_hd__nor2_2 _12582_ (.A(_05793_),
    .B(_05794_),
    .Y(_05795_));
 sky130_fd_sc_hd__a21oi_4 _12583_ (.A1(reg1_val[15]),
    .A2(_05024_),
    .B1(_05791_),
    .Y(_05797_));
 sky130_fd_sc_hd__or3_1 _12584_ (.A(_05793_),
    .B(_05794_),
    .C(_05797_),
    .X(_05798_));
 sky130_fd_sc_hd__xnor2_4 _12585_ (.A(_05795_),
    .B(_05797_),
    .Y(loadstore_address[16]));
 sky130_fd_sc_hd__nand2b_2 _12586_ (.A_N(_05794_),
    .B(_05798_),
    .Y(_05799_));
 sky130_fd_sc_hd__xnor2_2 _12587_ (.A(reg1_val[17]),
    .B(net278),
    .Y(_05800_));
 sky130_fd_sc_hd__xnor2_4 _12588_ (.A(_05799_),
    .B(_05800_),
    .Y(loadstore_address[17]));
 sky130_fd_sc_hd__or2_1 _12589_ (.A(reg1_val[18]),
    .B(net278),
    .X(_05801_));
 sky130_fd_sc_hd__nand2_1 _12590_ (.A(reg1_val[18]),
    .B(net278),
    .Y(_05802_));
 sky130_fd_sc_hd__nand2_2 _12591_ (.A(_05801_),
    .B(_05802_),
    .Y(_05803_));
 sky130_fd_sc_hd__or2_1 _12592_ (.A(_05798_),
    .B(_05800_),
    .X(_05804_));
 sky130_fd_sc_hd__a21bo_2 _12593_ (.A1(net278),
    .A2(_00239_),
    .B1_N(_05804_),
    .X(_05806_));
 sky130_fd_sc_hd__xnor2_4 _12594_ (.A(_05803_),
    .B(_05806_),
    .Y(loadstore_address[18]));
 sky130_fd_sc_hd__a21bo_1 _12595_ (.A1(_05801_),
    .A2(_05806_),
    .B1_N(_05802_),
    .X(_05807_));
 sky130_fd_sc_hd__xnor2_4 _12596_ (.A(reg1_val[19]),
    .B(net278),
    .Y(_05808_));
 sky130_fd_sc_hd__xnor2_4 _12597_ (.A(_05807_),
    .B(_05808_),
    .Y(loadstore_address[19]));
 sky130_fd_sc_hd__xnor2_2 _12598_ (.A(reg1_val[20]),
    .B(net278),
    .Y(_05809_));
 sky130_fd_sc_hd__or3_2 _12599_ (.A(_05803_),
    .B(_05804_),
    .C(_05808_),
    .X(_05810_));
 sky130_fd_sc_hd__nand2_1 _12600_ (.A(net278),
    .B(_00241_),
    .Y(_05811_));
 sky130_fd_sc_hd__a21oi_4 _12601_ (.A1(_05810_),
    .A2(_05811_),
    .B1(_05809_),
    .Y(_05812_));
 sky130_fd_sc_hd__and3_2 _12602_ (.A(_05809_),
    .B(_05810_),
    .C(_05811_),
    .X(_05813_));
 sky130_fd_sc_hd__nor2_8 _12603_ (.A(_05812_),
    .B(_05813_),
    .Y(loadstore_address[20]));
 sky130_fd_sc_hd__nor2_1 _12604_ (.A(reg1_val[21]),
    .B(net278),
    .Y(_05815_));
 sky130_fd_sc_hd__nand2_2 _12605_ (.A(reg1_val[21]),
    .B(net278),
    .Y(_05816_));
 sky130_fd_sc_hd__nand2b_2 _12606_ (.A_N(_05815_),
    .B(_05816_),
    .Y(_05817_));
 sky130_fd_sc_hd__a21oi_4 _12607_ (.A1(reg1_val[20]),
    .A2(net278),
    .B1(_05812_),
    .Y(_05818_));
 sky130_fd_sc_hd__xor2_4 _12608_ (.A(_05817_),
    .B(_05818_),
    .X(loadstore_address[21]));
 sky130_fd_sc_hd__or2_1 _12609_ (.A(reg1_val[22]),
    .B(net278),
    .X(_05819_));
 sky130_fd_sc_hd__nand2_1 _12610_ (.A(reg1_val[22]),
    .B(net278),
    .Y(_05820_));
 sky130_fd_sc_hd__nand2_2 _12611_ (.A(_05819_),
    .B(_05820_),
    .Y(_05821_));
 sky130_fd_sc_hd__o21ai_4 _12612_ (.A1(_05815_),
    .A2(_05818_),
    .B1(_05816_),
    .Y(_05822_));
 sky130_fd_sc_hd__xnor2_4 _12613_ (.A(_05821_),
    .B(_05822_),
    .Y(loadstore_address[22]));
 sky130_fd_sc_hd__a21bo_1 _12614_ (.A1(_05819_),
    .A2(_05822_),
    .B1_N(_05820_),
    .X(_05824_));
 sky130_fd_sc_hd__xnor2_2 _12615_ (.A(reg1_val[23]),
    .B(net278),
    .Y(_05825_));
 sky130_fd_sc_hd__xnor2_4 _12616_ (.A(_05824_),
    .B(_05825_),
    .Y(loadstore_address[23]));
 sky130_fd_sc_hd__or2_1 _12617_ (.A(reg1_val[24]),
    .B(net279),
    .X(_05826_));
 sky130_fd_sc_hd__nand2_1 _12618_ (.A(reg1_val[24]),
    .B(net279),
    .Y(_05827_));
 sky130_fd_sc_hd__nand2_2 _12619_ (.A(_05826_),
    .B(_05827_),
    .Y(_05828_));
 sky130_fd_sc_hd__or4_1 _12620_ (.A(_05809_),
    .B(_05817_),
    .C(_05821_),
    .D(_05825_),
    .X(_05829_));
 sky130_fd_sc_hd__a2bb2o_2 _12621_ (.A1_N(_05810_),
    .A2_N(_05829_),
    .B1(net278),
    .B2(_00243_),
    .X(_05830_));
 sky130_fd_sc_hd__nand2b_1 _12622_ (.A_N(_05828_),
    .B(_05830_),
    .Y(_05831_));
 sky130_fd_sc_hd__xnor2_4 _12623_ (.A(_05828_),
    .B(_05830_),
    .Y(loadstore_address[24]));
 sky130_fd_sc_hd__nand2_2 _12624_ (.A(_05827_),
    .B(_05831_),
    .Y(_05833_));
 sky130_fd_sc_hd__xnor2_2 _12625_ (.A(reg1_val[25]),
    .B(net279),
    .Y(_05834_));
 sky130_fd_sc_hd__xnor2_4 _12626_ (.A(_05833_),
    .B(_05834_),
    .Y(loadstore_address[25]));
 sky130_fd_sc_hd__or2_1 _12627_ (.A(reg1_val[26]),
    .B(net279),
    .X(_05835_));
 sky130_fd_sc_hd__nand2_1 _12628_ (.A(reg1_val[26]),
    .B(net279),
    .Y(_05836_));
 sky130_fd_sc_hd__nand2_2 _12629_ (.A(_05835_),
    .B(_05836_),
    .Y(_05837_));
 sky130_fd_sc_hd__or2_1 _12630_ (.A(_05831_),
    .B(_05834_),
    .X(_05838_));
 sky130_fd_sc_hd__a21bo_2 _12631_ (.A1(net279),
    .A2(_00245_),
    .B1_N(_05838_),
    .X(_05839_));
 sky130_fd_sc_hd__xnor2_4 _12632_ (.A(_05837_),
    .B(_05839_),
    .Y(loadstore_address[26]));
 sky130_fd_sc_hd__a21bo_1 _12633_ (.A1(_05835_),
    .A2(_05839_),
    .B1_N(_05836_),
    .X(_05841_));
 sky130_fd_sc_hd__xnor2_4 _12634_ (.A(reg1_val[27]),
    .B(net279),
    .Y(_05842_));
 sky130_fd_sc_hd__xnor2_4 _12635_ (.A(_05841_),
    .B(_05842_),
    .Y(loadstore_address[27]));
 sky130_fd_sc_hd__nor2_1 _12636_ (.A(reg1_val[28]),
    .B(net279),
    .Y(_05843_));
 sky130_fd_sc_hd__and2_1 _12637_ (.A(reg1_val[28]),
    .B(net279),
    .X(_05844_));
 sky130_fd_sc_hd__or2_1 _12638_ (.A(_05843_),
    .B(_05844_),
    .X(_05845_));
 sky130_fd_sc_hd__nand2_1 _12639_ (.A(net279),
    .B(_00329_),
    .Y(_05846_));
 sky130_fd_sc_hd__or3_2 _12640_ (.A(_05837_),
    .B(_05838_),
    .C(_05842_),
    .X(_05847_));
 sky130_fd_sc_hd__a21oi_4 _12641_ (.A1(_05846_),
    .A2(_05847_),
    .B1(_05845_),
    .Y(_05848_));
 sky130_fd_sc_hd__and3_2 _12642_ (.A(_05845_),
    .B(_05846_),
    .C(_05847_),
    .X(_05849_));
 sky130_fd_sc_hd__nor2_8 _12643_ (.A(_05848_),
    .B(_05849_),
    .Y(loadstore_address[28]));
 sky130_fd_sc_hd__nand2_1 _12644_ (.A(reg1_val[29]),
    .B(net279),
    .Y(_05851_));
 sky130_fd_sc_hd__or2_1 _12645_ (.A(reg1_val[29]),
    .B(net279),
    .X(_05852_));
 sky130_fd_sc_hd__nand2_2 _12646_ (.A(_05851_),
    .B(_05852_),
    .Y(_05853_));
 sky130_fd_sc_hd__or2_2 _12647_ (.A(_05844_),
    .B(_05848_),
    .X(_05854_));
 sky130_fd_sc_hd__xnor2_4 _12648_ (.A(_05853_),
    .B(_05854_),
    .Y(loadstore_address[29]));
 sky130_fd_sc_hd__or2_1 _12649_ (.A(reg1_val[30]),
    .B(net279),
    .X(_05855_));
 sky130_fd_sc_hd__nand2_1 _12650_ (.A(reg1_val[30]),
    .B(net279),
    .Y(_05856_));
 sky130_fd_sc_hd__nand2_2 _12651_ (.A(_05855_),
    .B(_05856_),
    .Y(_05857_));
 sky130_fd_sc_hd__a21bo_2 _12652_ (.A1(_05852_),
    .A2(_05854_),
    .B1_N(_05851_),
    .X(_05858_));
 sky130_fd_sc_hd__xnor2_4 _12653_ (.A(_05857_),
    .B(_05858_),
    .Y(loadstore_address[30]));
 sky130_fd_sc_hd__a21bo_1 _12654_ (.A1(_05855_),
    .A2(_05858_),
    .B1_N(_05856_),
    .X(_05860_));
 sky130_fd_sc_hd__xnor2_2 _12655_ (.A(reg1_val[31]),
    .B(_05860_),
    .Y(_05861_));
 sky130_fd_sc_hd__xnor2_4 _12656_ (.A(net279),
    .B(_05861_),
    .Y(loadstore_address[31]));
 sky130_fd_sc_hd__nand2_1 _12657_ (.A(net472),
    .B(net408),
    .Y(_05862_));
 sky130_fd_sc_hd__nand3_1 _12658_ (.A(net469),
    .B(net472),
    .C(net408),
    .Y(_05863_));
 sky130_fd_sc_hd__and4_1 _12659_ (.A(net441),
    .B(net469),
    .C(\div_counter[1] ),
    .D(net408),
    .X(_05864_));
 sky130_fd_sc_hd__inv_2 _12660_ (.A(_05864_),
    .Y(_05865_));
 sky130_fd_sc_hd__nand2_1 _12661_ (.A(net331),
    .B(net470),
    .Y(_05866_));
 sky130_fd_sc_hd__nor2_1 _12662_ (.A(net268),
    .B(net471),
    .Y(_05867_));
 sky130_fd_sc_hd__nor3_1 _12663_ (.A(rst),
    .B(net221),
    .C(_05867_),
    .Y(_00000_));
 sky130_fd_sc_hd__nor2_1 _12664_ (.A(net272),
    .B(_06397_),
    .Y(_05869_));
 sky130_fd_sc_hd__nand2_1 _12665_ (.A(net267),
    .B(_06396_),
    .Y(_05870_));
 sky130_fd_sc_hd__or2_1 _12666_ (.A(net341),
    .B(net201),
    .X(_05871_));
 sky130_fd_sc_hd__o211a_1 _12667_ (.A1(_00728_),
    .A2(net196),
    .B1(net342),
    .C1(net296),
    .X(_00001_));
 sky130_fd_sc_hd__nand2_1 _12668_ (.A(net226),
    .B(net201),
    .Y(_05872_));
 sky130_fd_sc_hd__o211a_1 _12669_ (.A1(net343),
    .A2(net201),
    .B1(_05872_),
    .C1(net294),
    .X(_00002_));
 sky130_fd_sc_hd__or2_1 _12670_ (.A(net361),
    .B(net201),
    .X(_05873_));
 sky130_fd_sc_hd__o211a_1 _12671_ (.A1(_00338_),
    .A2(net195),
    .B1(net362),
    .C1(net294),
    .X(_00003_));
 sky130_fd_sc_hd__or2_1 _12672_ (.A(net384),
    .B(net201),
    .X(_05874_));
 sky130_fd_sc_hd__o211a_1 _12673_ (.A1(_00424_),
    .A2(net195),
    .B1(net385),
    .C1(net294),
    .X(_00004_));
 sky130_fd_sc_hd__or2_1 _12674_ (.A(net380),
    .B(net201),
    .X(_05876_));
 sky130_fd_sc_hd__o211a_1 _12675_ (.A1(_00252_),
    .A2(net197),
    .B1(net381),
    .C1(net293),
    .X(_00005_));
 sky130_fd_sc_hd__or2_1 _12676_ (.A(net353),
    .B(net199),
    .X(_05877_));
 sky130_fd_sc_hd__o211a_1 _12677_ (.A1(_00263_),
    .A2(net197),
    .B1(net354),
    .C1(net293),
    .X(_00006_));
 sky130_fd_sc_hd__or2_1 _12678_ (.A(net359),
    .B(net201),
    .X(_05878_));
 sky130_fd_sc_hd__o211a_1 _12679_ (.A1(_00300_),
    .A2(net197),
    .B1(net360),
    .C1(net292),
    .X(_00007_));
 sky130_fd_sc_hd__or2_1 _12680_ (.A(net376),
    .B(net201),
    .X(_05879_));
 sky130_fd_sc_hd__o211a_1 _12681_ (.A1(_00310_),
    .A2(net196),
    .B1(net377),
    .C1(net294),
    .X(_00008_));
 sky130_fd_sc_hd__or2_1 _12682_ (.A(net382),
    .B(net200),
    .X(_05880_));
 sky130_fd_sc_hd__o211a_1 _12683_ (.A1(_00276_),
    .A2(net196),
    .B1(net383),
    .C1(net294),
    .X(_00009_));
 sky130_fd_sc_hd__nand2_1 _12684_ (.A(net144),
    .B(net200),
    .Y(_05882_));
 sky130_fd_sc_hd__o211a_1 _12685_ (.A1(net335),
    .A2(net200),
    .B1(_05882_),
    .C1(net296),
    .X(_00010_));
 sky130_fd_sc_hd__nand2_1 _12686_ (.A(net134),
    .B(net200),
    .Y(_05883_));
 sky130_fd_sc_hd__o211a_1 _12687_ (.A1(net333),
    .A2(net200),
    .B1(_05883_),
    .C1(net297),
    .X(_00011_));
 sky130_fd_sc_hd__nand2_1 _12688_ (.A(net91),
    .B(net201),
    .Y(_05884_));
 sky130_fd_sc_hd__o211a_1 _12689_ (.A1(net319),
    .A2(net201),
    .B1(_05884_),
    .C1(net296),
    .X(_00012_));
 sky130_fd_sc_hd__nand2_1 _12690_ (.A(net88),
    .B(net201),
    .Y(_05885_));
 sky130_fd_sc_hd__o211a_1 _12691_ (.A1(net323),
    .A2(net201),
    .B1(_05885_),
    .C1(net296),
    .X(_00013_));
 sky130_fd_sc_hd__or2_1 _12692_ (.A(net378),
    .B(net201),
    .X(_05886_));
 sky130_fd_sc_hd__o211a_1 _12693_ (.A1(_00430_),
    .A2(net197),
    .B1(net379),
    .C1(net292),
    .X(_00014_));
 sky130_fd_sc_hd__nand2_1 _12694_ (.A(net127),
    .B(net199),
    .Y(_05888_));
 sky130_fd_sc_hd__o211a_1 _12695_ (.A1(net317),
    .A2(net199),
    .B1(_05888_),
    .C1(net292),
    .X(_00015_));
 sky130_fd_sc_hd__or2_1 _12696_ (.A(net370),
    .B(net199),
    .X(_05889_));
 sky130_fd_sc_hd__o211a_1 _12697_ (.A1(_06483_),
    .A2(net197),
    .B1(net371),
    .C1(net292),
    .X(_00016_));
 sky130_fd_sc_hd__or2_1 _12698_ (.A(net355),
    .B(net199),
    .X(_05890_));
 sky130_fd_sc_hd__o211a_1 _12699_ (.A1(_06459_),
    .A2(net197),
    .B1(net356),
    .C1(net292),
    .X(_00017_));
 sky130_fd_sc_hd__or2_1 _12700_ (.A(net374),
    .B(net199),
    .X(_05891_));
 sky130_fd_sc_hd__o211a_1 _12701_ (.A1(_06467_),
    .A2(net197),
    .B1(net375),
    .C1(net291),
    .X(_00018_));
 sky130_fd_sc_hd__nand2_1 _12702_ (.A(net101),
    .B(net199),
    .Y(_05892_));
 sky130_fd_sc_hd__o211a_1 _12703_ (.A1(net313),
    .A2(net199),
    .B1(_05892_),
    .C1(net290),
    .X(_00019_));
 sky130_fd_sc_hd__nand2_1 _12704_ (.A(net120),
    .B(net198),
    .Y(_05894_));
 sky130_fd_sc_hd__o211a_1 _12705_ (.A1(net311),
    .A2(net198),
    .B1(_05894_),
    .C1(net290),
    .X(_00020_));
 sky130_fd_sc_hd__nand2_1 _12706_ (.A(net72),
    .B(net198),
    .Y(_05895_));
 sky130_fd_sc_hd__o211a_1 _12707_ (.A1(net309),
    .A2(net198),
    .B1(_05895_),
    .C1(net290),
    .X(_00021_));
 sky130_fd_sc_hd__or2_1 _12708_ (.A(net474),
    .B(net199),
    .X(_05896_));
 sky130_fd_sc_hd__o211a_1 _12709_ (.A1(_06503_),
    .A2(net197),
    .B1(net475),
    .C1(net292),
    .X(_00022_));
 sky130_fd_sc_hd__nand2_1 _12710_ (.A(net75),
    .B(net198),
    .Y(_05897_));
 sky130_fd_sc_hd__o211a_1 _12711_ (.A1(net321),
    .A2(net198),
    .B1(_05897_),
    .C1(net290),
    .X(_00023_));
 sky130_fd_sc_hd__nand2_1 _12712_ (.A(net69),
    .B(net198),
    .Y(_05898_));
 sky130_fd_sc_hd__o211a_1 _12713_ (.A1(net329),
    .A2(net198),
    .B1(_05898_),
    .C1(net290),
    .X(_00024_));
 sky130_fd_sc_hd__nand2_1 _12714_ (.A(net66),
    .B(net198),
    .Y(_05900_));
 sky130_fd_sc_hd__o211a_1 _12715_ (.A1(net325),
    .A2(net198),
    .B1(_05900_),
    .C1(net290),
    .X(_00025_));
 sky130_fd_sc_hd__nand2_1 _12716_ (.A(net59),
    .B(net198),
    .Y(_05901_));
 sky130_fd_sc_hd__o211a_1 _12717_ (.A1(net337),
    .A2(net198),
    .B1(_05901_),
    .C1(net290),
    .X(_00026_));
 sky130_fd_sc_hd__nand2_1 _12718_ (.A(net56),
    .B(net198),
    .Y(_05902_));
 sky130_fd_sc_hd__o211a_1 _12719_ (.A1(net327),
    .A2(net198),
    .B1(_05902_),
    .C1(net290),
    .X(_00027_));
 sky130_fd_sc_hd__nand2_1 _12720_ (.A(_00185_),
    .B(net198),
    .Y(_05903_));
 sky130_fd_sc_hd__o211a_1 _12721_ (.A1(net339),
    .A2(net198),
    .B1(_05903_),
    .C1(net290),
    .X(_00028_));
 sky130_fd_sc_hd__or2_1 _12722_ (.A(net403),
    .B(net199),
    .X(_05904_));
 sky130_fd_sc_hd__o211a_1 _12723_ (.A1(_00197_),
    .A2(net197),
    .B1(net404),
    .C1(net292),
    .X(_00029_));
 sky130_fd_sc_hd__or2_1 _12724_ (.A(net357),
    .B(net199),
    .X(_05906_));
 sky130_fd_sc_hd__o211a_1 _12725_ (.A1(_00222_),
    .A2(net197),
    .B1(net358),
    .C1(net292),
    .X(_00030_));
 sky130_fd_sc_hd__or2_1 _12726_ (.A(net389),
    .B(net199),
    .X(_05907_));
 sky130_fd_sc_hd__o211a_1 _12727_ (.A1(_00228_),
    .A2(net197),
    .B1(net390),
    .C1(net292),
    .X(_00031_));
 sky130_fd_sc_hd__nand2_1 _12728_ (.A(_00408_),
    .B(net199),
    .Y(_05908_));
 sky130_fd_sc_hd__o211a_1 _12729_ (.A1(net315),
    .A2(net199),
    .B1(_05908_),
    .C1(net293),
    .X(_00032_));
 sky130_fd_sc_hd__or2_1 _12730_ (.A(net372),
    .B(net199),
    .X(_05909_));
 sky130_fd_sc_hd__o211a_1 _12731_ (.A1(_00756_),
    .A2(net197),
    .B1(net373),
    .C1(net293),
    .X(_00033_));
 sky130_fd_sc_hd__or2_1 _12732_ (.A(_04351_),
    .B(net315),
    .X(_05910_));
 sky130_fd_sc_hd__nand2_1 _12733_ (.A(_04351_),
    .B(net315),
    .Y(_05912_));
 sky130_fd_sc_hd__nand2_1 _12734_ (.A(_05910_),
    .B(_05912_),
    .Y(_05913_));
 sky130_fd_sc_hd__and2b_1 _12735_ (.A_N(net389),
    .B(net601),
    .X(_05914_));
 sky130_fd_sc_hd__nand2b_1 _12736_ (.A_N(net601),
    .B(net389),
    .Y(_05915_));
 sky130_fd_sc_hd__and2b_1 _12737_ (.A_N(net357),
    .B(net583),
    .X(_05916_));
 sky130_fd_sc_hd__and2b_1 _12738_ (.A_N(net403),
    .B(net573),
    .X(_05917_));
 sky130_fd_sc_hd__nand2b_1 _12739_ (.A_N(net573),
    .B(net403),
    .Y(_05918_));
 sky130_fd_sc_hd__and2b_1 _12740_ (.A_N(net339),
    .B(net589),
    .X(_05919_));
 sky130_fd_sc_hd__nand2b_1 _12741_ (.A_N(net607),
    .B(net339),
    .Y(_05920_));
 sky130_fd_sc_hd__nand2b_1 _12742_ (.A_N(_05919_),
    .B(_05920_),
    .Y(_05921_));
 sky130_fd_sc_hd__and2b_1 _12743_ (.A_N(net327),
    .B(net579),
    .X(_05923_));
 sky130_fd_sc_hd__nand2b_1 _12744_ (.A_N(net579),
    .B(net327),
    .Y(_05924_));
 sky130_fd_sc_hd__and2b_1 _12745_ (.A_N(net337),
    .B(\div_shifter[55] ),
    .X(_05925_));
 sky130_fd_sc_hd__and2b_1 _12746_ (.A_N(net325),
    .B(net599),
    .X(_05926_));
 sky130_fd_sc_hd__nand2b_1 _12747_ (.A_N(net599),
    .B(net325),
    .Y(_05927_));
 sky130_fd_sc_hd__and2b_1 _12748_ (.A_N(net329),
    .B(net577),
    .X(_05928_));
 sky130_fd_sc_hd__and2b_1 _12749_ (.A_N(net321),
    .B(net571),
    .X(_05929_));
 sky130_fd_sc_hd__nand2b_1 _12750_ (.A_N(net571),
    .B(net321),
    .Y(_05930_));
 sky130_fd_sc_hd__and2b_1 _12751_ (.A_N(net474),
    .B(\div_shifter[51] ),
    .X(_05931_));
 sky130_fd_sc_hd__and2b_1 _12752_ (.A_N(net309),
    .B(\div_shifter[50] ),
    .X(_05932_));
 sky130_fd_sc_hd__nand2b_1 _12753_ (.A_N(\div_shifter[50] ),
    .B(net309),
    .Y(_05934_));
 sky130_fd_sc_hd__nand2b_1 _12754_ (.A_N(\div_shifter[49] ),
    .B(net311),
    .Y(_05935_));
 sky130_fd_sc_hd__and2b_1 _12755_ (.A_N(net313),
    .B(net561),
    .X(_05936_));
 sky130_fd_sc_hd__nand2b_1 _12756_ (.A_N(net561),
    .B(net313),
    .Y(_05937_));
 sky130_fd_sc_hd__and2b_1 _12757_ (.A_N(net374),
    .B(net575),
    .X(_05938_));
 sky130_fd_sc_hd__nand2b_1 _12758_ (.A_N(net575),
    .B(net374),
    .Y(_05939_));
 sky130_fd_sc_hd__and2b_1 _12759_ (.A_N(net355),
    .B(\div_shifter[46] ),
    .X(_05940_));
 sky130_fd_sc_hd__nand2b_1 _12760_ (.A_N(\div_shifter[46] ),
    .B(net355),
    .Y(_05941_));
 sky130_fd_sc_hd__and2b_1 _12761_ (.A_N(net370),
    .B(\div_shifter[45] ),
    .X(_05942_));
 sky130_fd_sc_hd__nand2b_1 _12762_ (.A_N(\div_shifter[45] ),
    .B(net370),
    .Y(_05943_));
 sky130_fd_sc_hd__and2b_1 _12763_ (.A_N(net317),
    .B(net567),
    .X(_05945_));
 sky130_fd_sc_hd__nand2b_1 _12764_ (.A_N(net567),
    .B(net317),
    .Y(_05946_));
 sky130_fd_sc_hd__and2b_1 _12765_ (.A_N(net378),
    .B(net569),
    .X(_05947_));
 sky130_fd_sc_hd__nand2b_1 _12766_ (.A_N(net569),
    .B(net378),
    .Y(_05948_));
 sky130_fd_sc_hd__and2b_1 _12767_ (.A_N(net323),
    .B(\div_shifter[42] ),
    .X(_05949_));
 sky130_fd_sc_hd__nand2b_1 _12768_ (.A_N(\div_shifter[42] ),
    .B(net323),
    .Y(_05950_));
 sky130_fd_sc_hd__and2b_1 _12769_ (.A_N(net319),
    .B(net563),
    .X(_05951_));
 sky130_fd_sc_hd__nand2b_1 _12770_ (.A_N(net563),
    .B(net319),
    .Y(_05952_));
 sky130_fd_sc_hd__and2b_1 _12771_ (.A_N(net333),
    .B(\div_shifter[40] ),
    .X(_05953_));
 sky130_fd_sc_hd__nand2b_1 _12772_ (.A_N(\div_shifter[40] ),
    .B(net333),
    .Y(_05954_));
 sky130_fd_sc_hd__and2b_1 _12773_ (.A_N(net335),
    .B(\div_shifter[39] ),
    .X(_05956_));
 sky130_fd_sc_hd__nand2b_1 _12774_ (.A_N(\div_shifter[39] ),
    .B(net335),
    .Y(_05957_));
 sky130_fd_sc_hd__and2b_1 _12775_ (.A_N(net382),
    .B(net597),
    .X(_05958_));
 sky130_fd_sc_hd__nand2b_1 _12776_ (.A_N(net597),
    .B(net382),
    .Y(_05959_));
 sky130_fd_sc_hd__and2b_1 _12777_ (.A_N(net376),
    .B(net593),
    .X(_05960_));
 sky130_fd_sc_hd__nand2b_1 _12778_ (.A_N(net593),
    .B(net376),
    .Y(_05961_));
 sky130_fd_sc_hd__and2b_1 _12779_ (.A_N(net359),
    .B(\div_shifter[36] ),
    .X(_05962_));
 sky130_fd_sc_hd__nand2b_1 _12780_ (.A_N(\div_shifter[36] ),
    .B(net359),
    .Y(_05963_));
 sky130_fd_sc_hd__nand2b_1 _12781_ (.A_N(_05962_),
    .B(_05963_),
    .Y(_05964_));
 sky130_fd_sc_hd__and2b_1 _12782_ (.A_N(net353),
    .B(net565),
    .X(_05965_));
 sky130_fd_sc_hd__nand2b_1 _12783_ (.A_N(net565),
    .B(net353),
    .Y(_05967_));
 sky130_fd_sc_hd__nand2b_1 _12784_ (.A_N(_05965_),
    .B(_05967_),
    .Y(_05968_));
 sky130_fd_sc_hd__and2b_1 _12785_ (.A_N(net380),
    .B(\div_shifter[34] ),
    .X(_05969_));
 sky130_fd_sc_hd__nand2b_1 _12786_ (.A_N(\div_shifter[34] ),
    .B(net380),
    .Y(_05970_));
 sky130_fd_sc_hd__and2b_1 _12787_ (.A_N(net384),
    .B(net551),
    .X(_05971_));
 sky130_fd_sc_hd__nand2b_1 _12788_ (.A_N(net551),
    .B(net384),
    .Y(_05972_));
 sky130_fd_sc_hd__and2b_1 _12789_ (.A_N(net361),
    .B(net557),
    .X(_05973_));
 sky130_fd_sc_hd__and2b_1 _12790_ (.A_N(\div_shifter[32] ),
    .B(net361),
    .X(_05974_));
 sky130_fd_sc_hd__nor2_1 _12791_ (.A(_05973_),
    .B(_05974_),
    .Y(_05975_));
 sky130_fd_sc_hd__nand2b_1 _12792_ (.A_N(net345),
    .B(net343),
    .Y(_05976_));
 sky130_fd_sc_hd__a21o_1 _12793_ (.A1(_05975_),
    .A2(_05976_),
    .B1(_05973_),
    .X(_05978_));
 sky130_fd_sc_hd__a21o_1 _12794_ (.A1(_05972_),
    .A2(_05978_),
    .B1(_05971_),
    .X(_05979_));
 sky130_fd_sc_hd__a21o_1 _12795_ (.A1(_05970_),
    .A2(_05979_),
    .B1(_05969_),
    .X(_05980_));
 sky130_fd_sc_hd__a21o_1 _12796_ (.A1(_05967_),
    .A2(_05980_),
    .B1(_05965_),
    .X(_05981_));
 sky130_fd_sc_hd__a21o_1 _12797_ (.A1(_05963_),
    .A2(_05981_),
    .B1(_05962_),
    .X(_05982_));
 sky130_fd_sc_hd__a21o_1 _12798_ (.A1(_05961_),
    .A2(_05982_),
    .B1(_05960_),
    .X(_05983_));
 sky130_fd_sc_hd__a21o_1 _12799_ (.A1(_05959_),
    .A2(_05983_),
    .B1(_05958_),
    .X(_05984_));
 sky130_fd_sc_hd__a21o_1 _12800_ (.A1(_05957_),
    .A2(_05984_),
    .B1(_05956_),
    .X(_05985_));
 sky130_fd_sc_hd__a21o_1 _12801_ (.A1(_05954_),
    .A2(_05985_),
    .B1(_05953_),
    .X(_05986_));
 sky130_fd_sc_hd__a21o_1 _12802_ (.A1(_05952_),
    .A2(_05986_),
    .B1(_05951_),
    .X(_05987_));
 sky130_fd_sc_hd__a21o_1 _12803_ (.A1(_05950_),
    .A2(_05987_),
    .B1(_05949_),
    .X(_05989_));
 sky130_fd_sc_hd__a21o_1 _12804_ (.A1(_05948_),
    .A2(_05989_),
    .B1(_05947_),
    .X(_05990_));
 sky130_fd_sc_hd__a21o_1 _12805_ (.A1(_05946_),
    .A2(_05990_),
    .B1(_05945_),
    .X(_05991_));
 sky130_fd_sc_hd__a21o_1 _12806_ (.A1(_05943_),
    .A2(_05991_),
    .B1(_05942_),
    .X(_05992_));
 sky130_fd_sc_hd__a21o_1 _12807_ (.A1(_05941_),
    .A2(_05992_),
    .B1(_05940_),
    .X(_05993_));
 sky130_fd_sc_hd__a21o_1 _12808_ (.A1(_05939_),
    .A2(_05993_),
    .B1(_05938_),
    .X(_05994_));
 sky130_fd_sc_hd__a21o_1 _12809_ (.A1(_05937_),
    .A2(_05994_),
    .B1(_05936_),
    .X(_05995_));
 sky130_fd_sc_hd__nand2b_1 _12810_ (.A_N(net311),
    .B(\div_shifter[49] ),
    .Y(_05996_));
 sky130_fd_sc_hd__a21bo_1 _12811_ (.A1(_05935_),
    .A2(_05995_),
    .B1_N(_05996_),
    .X(_05997_));
 sky130_fd_sc_hd__a21o_1 _12812_ (.A1(_05934_),
    .A2(_05997_),
    .B1(_05932_),
    .X(_05998_));
 sky130_fd_sc_hd__nand2b_1 _12813_ (.A_N(\div_shifter[51] ),
    .B(net474),
    .Y(_06000_));
 sky130_fd_sc_hd__nand2b_1 _12814_ (.A_N(_05931_),
    .B(_06000_),
    .Y(_06001_));
 sky130_fd_sc_hd__a21o_1 _12815_ (.A1(_05998_),
    .A2(_06000_),
    .B1(_05931_),
    .X(_06002_));
 sky130_fd_sc_hd__a21o_1 _12816_ (.A1(_05930_),
    .A2(_06002_),
    .B1(_05929_),
    .X(_06003_));
 sky130_fd_sc_hd__nand2b_1 _12817_ (.A_N(net577),
    .B(net329),
    .Y(_06004_));
 sky130_fd_sc_hd__nand2b_1 _12818_ (.A_N(_05928_),
    .B(_06004_),
    .Y(_06005_));
 sky130_fd_sc_hd__a21o_1 _12819_ (.A1(_06003_),
    .A2(_06004_),
    .B1(_05928_),
    .X(_06006_));
 sky130_fd_sc_hd__a21o_1 _12820_ (.A1(_05927_),
    .A2(_06006_),
    .B1(_05926_),
    .X(_06007_));
 sky130_fd_sc_hd__nand2b_1 _12821_ (.A_N(\div_shifter[55] ),
    .B(net337),
    .Y(_06008_));
 sky130_fd_sc_hd__nand2b_1 _12822_ (.A_N(_05925_),
    .B(_06008_),
    .Y(_06009_));
 sky130_fd_sc_hd__a21o_1 _12823_ (.A1(_06007_),
    .A2(_06008_),
    .B1(_05925_),
    .X(_06011_));
 sky130_fd_sc_hd__a21o_1 _12824_ (.A1(_05924_),
    .A2(_06011_),
    .B1(_05923_),
    .X(_06012_));
 sky130_fd_sc_hd__a21o_1 _12825_ (.A1(_05920_),
    .A2(_06012_),
    .B1(_05919_),
    .X(_06013_));
 sky130_fd_sc_hd__a21oi_1 _12826_ (.A1(_05918_),
    .A2(_06013_),
    .B1(_05917_),
    .Y(_06014_));
 sky130_fd_sc_hd__and2b_1 _12827_ (.A_N(net583),
    .B(net357),
    .X(_06015_));
 sky130_fd_sc_hd__nor2_1 _12828_ (.A(_05916_),
    .B(_06015_),
    .Y(_06016_));
 sky130_fd_sc_hd__o21bai_2 _12829_ (.A1(_06014_),
    .A2(_06015_),
    .B1_N(_05916_),
    .Y(_06017_));
 sky130_fd_sc_hd__a21oi_1 _12830_ (.A1(_05915_),
    .A2(_06017_),
    .B1(_05914_),
    .Y(_06018_));
 sky130_fd_sc_hd__or2_1 _12831_ (.A(_05913_),
    .B(_06018_),
    .X(_06019_));
 sky130_fd_sc_hd__and3_1 _12832_ (.A(net372),
    .B(_05910_),
    .C(_06019_),
    .X(_06020_));
 sky130_fd_sc_hd__a21oi_1 _12833_ (.A1(_05910_),
    .A2(_06019_),
    .B1(net372),
    .Y(_06022_));
 sky130_fd_sc_hd__o21bai_1 _12834_ (.A1(_04340_),
    .A2(_06020_),
    .B1_N(_06022_),
    .Y(_06023_));
 sky130_fd_sc_hd__a22o_1 _12835_ (.A1(net497),
    .A2(net220),
    .B1(net2),
    .B2(net271),
    .X(_06024_));
 sky130_fd_sc_hd__and2_1 _12836_ (.A(net291),
    .B(_06024_),
    .X(_00034_));
 sky130_fd_sc_hd__a22o_1 _12837_ (.A1(net497),
    .A2(net485),
    .B1(net220),
    .B2(\div_res[1] ),
    .X(_06025_));
 sky130_fd_sc_hd__and2_1 _12838_ (.A(net291),
    .B(net498),
    .X(_00035_));
 sky130_fd_sc_hd__a22o_1 _12839_ (.A1(\div_res[1] ),
    .A2(net269),
    .B1(net218),
    .B2(net555),
    .X(_06026_));
 sky130_fd_sc_hd__and2_1 _12840_ (.A(net288),
    .B(net556),
    .X(_00036_));
 sky130_fd_sc_hd__a22o_1 _12841_ (.A1(\div_res[2] ),
    .A2(net269),
    .B1(net218),
    .B2(net502),
    .X(_06027_));
 sky130_fd_sc_hd__and2_1 _12842_ (.A(net288),
    .B(net503),
    .X(_00037_));
 sky130_fd_sc_hd__a22o_1 _12843_ (.A1(net502),
    .A2(net269),
    .B1(net218),
    .B2(net547),
    .X(_06029_));
 sky130_fd_sc_hd__and2_1 _12844_ (.A(net288),
    .B(net548),
    .X(_00038_));
 sky130_fd_sc_hd__a22o_1 _12845_ (.A1(\div_res[4] ),
    .A2(net269),
    .B1(net218),
    .B2(net530),
    .X(_06030_));
 sky130_fd_sc_hd__and2_1 _12846_ (.A(net288),
    .B(net531),
    .X(_00039_));
 sky130_fd_sc_hd__a22o_1 _12847_ (.A1(\div_res[5] ),
    .A2(net269),
    .B1(net218),
    .B2(net521),
    .X(_06031_));
 sky130_fd_sc_hd__and2_1 _12848_ (.A(net288),
    .B(net522),
    .X(_00040_));
 sky130_fd_sc_hd__a22o_1 _12849_ (.A1(net521),
    .A2(net269),
    .B1(net218),
    .B2(net549),
    .X(_06032_));
 sky130_fd_sc_hd__and2_1 _12850_ (.A(net288),
    .B(net550),
    .X(_00041_));
 sky130_fd_sc_hd__a22o_1 _12851_ (.A1(\div_res[7] ),
    .A2(net269),
    .B1(net218),
    .B2(net508),
    .X(_06033_));
 sky130_fd_sc_hd__and2_1 _12852_ (.A(net288),
    .B(net509),
    .X(_00042_));
 sky130_fd_sc_hd__a22o_1 _12853_ (.A1(\div_res[8] ),
    .A2(net269),
    .B1(net218),
    .B2(net505),
    .X(_06035_));
 sky130_fd_sc_hd__and2_1 _12854_ (.A(net288),
    .B(net506),
    .X(_00043_));
 sky130_fd_sc_hd__a22o_1 _12855_ (.A1(net505),
    .A2(net269),
    .B1(net218),
    .B2(net494),
    .X(_06036_));
 sky130_fd_sc_hd__and2_1 _12856_ (.A(net288),
    .B(net512),
    .X(_00044_));
 sky130_fd_sc_hd__a22o_1 _12857_ (.A1(net494),
    .A2(net269),
    .B1(net218),
    .B2(\div_res[11] ),
    .X(_06037_));
 sky130_fd_sc_hd__and2_1 _12858_ (.A(net288),
    .B(net495),
    .X(_00045_));
 sky130_fd_sc_hd__a22o_1 _12859_ (.A1(\div_res[11] ),
    .A2(net269),
    .B1(net218),
    .B2(net515),
    .X(_06038_));
 sky130_fd_sc_hd__and2_1 _12860_ (.A(net289),
    .B(net516),
    .X(_00046_));
 sky130_fd_sc_hd__a22o_1 _12861_ (.A1(net515),
    .A2(net269),
    .B1(net218),
    .B2(net513),
    .X(_06039_));
 sky130_fd_sc_hd__and2_1 _12862_ (.A(net289),
    .B(net525),
    .X(_00047_));
 sky130_fd_sc_hd__a22o_1 _12863_ (.A1(net513),
    .A2(net270),
    .B1(net219),
    .B2(net479),
    .X(_06041_));
 sky130_fd_sc_hd__and2_1 _12864_ (.A(net289),
    .B(net514),
    .X(_00048_));
 sky130_fd_sc_hd__a22o_1 _12865_ (.A1(net479),
    .A2(net270),
    .B1(net219),
    .B2(\div_res[15] ),
    .X(_06042_));
 sky130_fd_sc_hd__and2_1 _12866_ (.A(net289),
    .B(net480),
    .X(_00049_));
 sky130_fd_sc_hd__a22o_1 _12867_ (.A1(net526),
    .A2(net270),
    .B1(net219),
    .B2(net492),
    .X(_06043_));
 sky130_fd_sc_hd__and2_1 _12868_ (.A(net289),
    .B(net527),
    .X(_00050_));
 sky130_fd_sc_hd__a22o_1 _12869_ (.A1(net492),
    .A2(net270),
    .B1(net219),
    .B2(net487),
    .X(_06044_));
 sky130_fd_sc_hd__and2_1 _12870_ (.A(net289),
    .B(net493),
    .X(_00051_));
 sky130_fd_sc_hd__a22o_1 _12871_ (.A1(net487),
    .A2(net270),
    .B1(net219),
    .B2(\div_res[18] ),
    .X(_06045_));
 sky130_fd_sc_hd__and2_1 _12872_ (.A(net289),
    .B(net488),
    .X(_00052_));
 sky130_fd_sc_hd__a22o_1 _12873_ (.A1(net490),
    .A2(net270),
    .B1(net219),
    .B2(net476),
    .X(_06047_));
 sky130_fd_sc_hd__and2_1 _12874_ (.A(net288),
    .B(net491),
    .X(_00053_));
 sky130_fd_sc_hd__a22o_1 _12875_ (.A1(net476),
    .A2(net269),
    .B1(net218),
    .B2(\div_res[20] ),
    .X(_06048_));
 sky130_fd_sc_hd__and2_1 _12876_ (.A(net289),
    .B(net477),
    .X(_00054_));
 sky130_fd_sc_hd__a22o_1 _12877_ (.A1(net518),
    .A2(net269),
    .B1(net218),
    .B2(\div_res[21] ),
    .X(_06049_));
 sky130_fd_sc_hd__and2_1 _12878_ (.A(net289),
    .B(net519),
    .X(_00055_));
 sky130_fd_sc_hd__a22o_1 _12879_ (.A1(\div_res[21] ),
    .A2(net269),
    .B1(net218),
    .B2(net499),
    .X(_06050_));
 sky130_fd_sc_hd__and2_1 _12880_ (.A(net288),
    .B(net500),
    .X(_00056_));
 sky130_fd_sc_hd__a22o_1 _12881_ (.A1(net499),
    .A2(net270),
    .B1(net219),
    .B2(net528),
    .X(_06051_));
 sky130_fd_sc_hd__and2_1 _12882_ (.A(net288),
    .B(net529),
    .X(_00057_));
 sky130_fd_sc_hd__a22o_1 _12883_ (.A1(net528),
    .A2(net270),
    .B1(net219),
    .B2(net539),
    .X(_06053_));
 sky130_fd_sc_hd__and2_1 _12884_ (.A(net289),
    .B(net540),
    .X(_00058_));
 sky130_fd_sc_hd__a22o_1 _12885_ (.A1(\div_res[24] ),
    .A2(net269),
    .B1(net218),
    .B2(net536),
    .X(_06054_));
 sky130_fd_sc_hd__and2_1 _12886_ (.A(net288),
    .B(net537),
    .X(_00059_));
 sky130_fd_sc_hd__a22o_1 _12887_ (.A1(net536),
    .A2(net271),
    .B1(net219),
    .B2(net543),
    .X(_06055_));
 sky130_fd_sc_hd__and2_1 _12888_ (.A(net290),
    .B(net544),
    .X(_00060_));
 sky130_fd_sc_hd__a22o_1 _12889_ (.A1(\div_res[26] ),
    .A2(net271),
    .B1(net220),
    .B2(net533),
    .X(_06056_));
 sky130_fd_sc_hd__and2_1 _12890_ (.A(net290),
    .B(net534),
    .X(_00061_));
 sky130_fd_sc_hd__a22o_1 _12891_ (.A1(net533),
    .A2(net271),
    .B1(net220),
    .B2(net541),
    .X(_06057_));
 sky130_fd_sc_hd__and2_1 _12892_ (.A(net291),
    .B(net546),
    .X(_00062_));
 sky130_fd_sc_hd__a22o_1 _12893_ (.A1(net541),
    .A2(net271),
    .B1(net220),
    .B2(net482),
    .X(_06059_));
 sky130_fd_sc_hd__and2_1 _12894_ (.A(net291),
    .B(net542),
    .X(_00063_));
 sky130_fd_sc_hd__a22o_1 _12895_ (.A1(net482),
    .A2(net271),
    .B1(net220),
    .B2(\div_res[30] ),
    .X(_06060_));
 sky130_fd_sc_hd__and2_1 _12896_ (.A(net291),
    .B(net483),
    .X(_00064_));
 sky130_fd_sc_hd__a22o_1 _12897_ (.A1(\div_res[30] ),
    .A2(net271),
    .B1(net220),
    .B2(net436),
    .X(_06061_));
 sky130_fd_sc_hd__and2_1 _12898_ (.A(net291),
    .B(net437),
    .X(_00065_));
 sky130_fd_sc_hd__a22o_1 _12899_ (.A1(net398),
    .A2(net221),
    .B1(net200),
    .B2(net304),
    .X(_06062_));
 sky130_fd_sc_hd__and2_1 _12900_ (.A(net296),
    .B(net399),
    .X(_00066_));
 sky130_fd_sc_hd__o221a_1 _12901_ (.A1(net398),
    .A2(net268),
    .B1(net217),
    .B2(net432),
    .C1(net296),
    .X(_06063_));
 sky130_fd_sc_hd__o21a_1 _12902_ (.A1(_00187_),
    .A2(net196),
    .B1(net433),
    .X(_00067_));
 sky130_fd_sc_hd__o221a_1 _12903_ (.A1(net432),
    .A2(net268),
    .B1(net217),
    .B2(net460),
    .C1(net296),
    .X(_06065_));
 sky130_fd_sc_hd__a21boi_1 _12904_ (.A1(_00190_),
    .A2(_05869_),
    .B1_N(net461),
    .Y(_00068_));
 sky130_fd_sc_hd__o221a_1 _12905_ (.A1(\div_shifter[2] ),
    .A2(net268),
    .B1(net217),
    .B2(net418),
    .C1(net296),
    .X(_06066_));
 sky130_fd_sc_hd__o21a_1 _12906_ (.A1(_00180_),
    .A2(net196),
    .B1(net419),
    .X(_00069_));
 sky130_fd_sc_hd__o221a_1 _12907_ (.A1(net418),
    .A2(net268),
    .B1(net217),
    .B2(net439),
    .C1(net296),
    .X(_06067_));
 sky130_fd_sc_hd__a21boi_1 _12908_ (.A1(_00204_),
    .A2(net200),
    .B1_N(net440),
    .Y(_00070_));
 sky130_fd_sc_hd__o221a_1 _12909_ (.A1(net439),
    .A2(net268),
    .B1(net217),
    .B2(net454),
    .C1(net297),
    .X(_06068_));
 sky130_fd_sc_hd__a21boi_1 _12910_ (.A1(net211),
    .A2(net200),
    .B1_N(net455),
    .Y(_00071_));
 sky130_fd_sc_hd__o221a_1 _12911_ (.A1(net454),
    .A2(net268),
    .B1(net217),
    .B2(net452),
    .C1(net296),
    .X(_06069_));
 sky130_fd_sc_hd__a21boi_1 _12912_ (.A1(_00161_),
    .A2(net200),
    .B1_N(net457),
    .Y(_00072_));
 sky130_fd_sc_hd__o221a_1 _12913_ (.A1(net452),
    .A2(net268),
    .B1(net217),
    .B2(net427),
    .C1(net297),
    .X(_06071_));
 sky130_fd_sc_hd__a21boi_1 _12914_ (.A1(net190),
    .A2(net201),
    .B1_N(net453),
    .Y(_00073_));
 sky130_fd_sc_hd__o221a_1 _12915_ (.A1(net427),
    .A2(net268),
    .B1(net217),
    .B2(\div_shifter[8] ),
    .C1(net295),
    .X(_06072_));
 sky130_fd_sc_hd__a21boi_1 _12916_ (.A1(_06494_),
    .A2(net200),
    .B1_N(net428),
    .Y(_00074_));
 sky130_fd_sc_hd__o221a_1 _12917_ (.A1(\div_shifter[8] ),
    .A2(net268),
    .B1(net217),
    .B2(net405),
    .C1(net295),
    .X(_06073_));
 sky130_fd_sc_hd__o21a_1 _12918_ (.A1(_06490_),
    .A2(net196),
    .B1(net406),
    .X(_00075_));
 sky130_fd_sc_hd__o221a_1 _12919_ (.A1(net405),
    .A2(net268),
    .B1(net217),
    .B2(net458),
    .C1(net295),
    .X(_06074_));
 sky130_fd_sc_hd__a21boi_1 _12920_ (.A1(_00147_),
    .A2(net200),
    .B1_N(net466),
    .Y(_00076_));
 sky130_fd_sc_hd__o221a_1 _12921_ (.A1(net458),
    .A2(net267),
    .B1(net217),
    .B2(net444),
    .C1(net295),
    .X(_06075_));
 sky130_fd_sc_hd__a21boi_1 _12922_ (.A1(net180),
    .A2(net200),
    .B1_N(net459),
    .Y(_00077_));
 sky130_fd_sc_hd__o221a_1 _12923_ (.A1(net444),
    .A2(net267),
    .B1(net216),
    .B2(net350),
    .C1(net294),
    .X(_06077_));
 sky130_fd_sc_hd__a21boi_1 _12924_ (.A1(_06440_),
    .A2(net200),
    .B1_N(net445),
    .Y(_00078_));
 sky130_fd_sc_hd__o221a_1 _12925_ (.A1(net350),
    .A2(net267),
    .B1(net216),
    .B2(\div_shifter[13] ),
    .C1(net294),
    .X(_06078_));
 sky130_fd_sc_hd__o21a_1 _12926_ (.A1(_06435_),
    .A2(net196),
    .B1(net351),
    .X(_00079_));
 sky130_fd_sc_hd__o221a_1 _12927_ (.A1(\div_shifter[13] ),
    .A2(net267),
    .B1(net216),
    .B2(net449),
    .C1(net294),
    .X(_06079_));
 sky130_fd_sc_hd__a21boi_1 _12928_ (.A1(_06474_),
    .A2(net201),
    .B1_N(net450),
    .Y(_00080_));
 sky130_fd_sc_hd__o221a_1 _12929_ (.A1(\div_shifter[14] ),
    .A2(net267),
    .B1(net216),
    .B2(net393),
    .C1(net294),
    .X(_06080_));
 sky130_fd_sc_hd__o21a_1 _12930_ (.A1(net155),
    .A2(net195),
    .B1(net394),
    .X(_00081_));
 sky130_fd_sc_hd__o221a_1 _12931_ (.A1(net393),
    .A2(net267),
    .B1(net216),
    .B2(net391),
    .C1(net294),
    .X(_06081_));
 sky130_fd_sc_hd__o21a_1 _12932_ (.A1(_00386_),
    .A2(net195),
    .B1(net397),
    .X(_00082_));
 sky130_fd_sc_hd__o221a_1 _12933_ (.A1(net391),
    .A2(net267),
    .B1(net216),
    .B2(net347),
    .C1(net294),
    .X(_06083_));
 sky130_fd_sc_hd__o21a_1 _12934_ (.A1(net138),
    .A2(net195),
    .B1(net392),
    .X(_00083_));
 sky130_fd_sc_hd__o221a_1 _12935_ (.A1(net347),
    .A2(net267),
    .B1(net216),
    .B2(\div_shifter[18] ),
    .C1(net294),
    .X(_06084_));
 sky130_fd_sc_hd__o21a_1 _12936_ (.A1(_00451_),
    .A2(net195),
    .B1(net348),
    .X(_00084_));
 sky130_fd_sc_hd__o221a_1 _12937_ (.A1(\div_shifter[18] ),
    .A2(net267),
    .B1(net216),
    .B2(net424),
    .C1(net294),
    .X(_06085_));
 sky130_fd_sc_hd__o21a_1 _12938_ (.A1(net136),
    .A2(net195),
    .B1(net425),
    .X(_00085_));
 sky130_fd_sc_hd__o221a_1 _12939_ (.A1(net424),
    .A2(net267),
    .B1(net216),
    .B2(net463),
    .C1(net294),
    .X(_06086_));
 sky130_fd_sc_hd__a21boi_1 _12940_ (.A1(_00437_),
    .A2(net200),
    .B1_N(net464),
    .Y(_00086_));
 sky130_fd_sc_hd__o221a_1 _12941_ (.A1(\div_shifter[20] ),
    .A2(net267),
    .B1(net216),
    .B2(net411),
    .C1(net295),
    .X(_06087_));
 sky130_fd_sc_hd__o21a_1 _12942_ (.A1(net103),
    .A2(net195),
    .B1(net412),
    .X(_00087_));
 sky130_fd_sc_hd__o221a_1 _12943_ (.A1(net411),
    .A2(net268),
    .B1(net217),
    .B2(net430),
    .C1(net295),
    .X(_06089_));
 sky130_fd_sc_hd__o21a_1 _12944_ (.A1(_00284_),
    .A2(net195),
    .B1(net431),
    .X(_00088_));
 sky130_fd_sc_hd__o221a_1 _12945_ (.A1(\div_shifter[22] ),
    .A2(net268),
    .B1(net216),
    .B2(net421),
    .C1(net295),
    .X(_06090_));
 sky130_fd_sc_hd__o21a_1 _12946_ (.A1(net107),
    .A2(net195),
    .B1(net422),
    .X(_00089_));
 sky130_fd_sc_hd__o221a_1 _12947_ (.A1(\div_shifter[23] ),
    .A2(net267),
    .B1(net216),
    .B2(net400),
    .C1(net295),
    .X(_06091_));
 sky130_fd_sc_hd__o21a_1 _12948_ (.A1(_00301_),
    .A2(net195),
    .B1(net401),
    .X(_00090_));
 sky130_fd_sc_hd__o221a_1 _12949_ (.A1(net400),
    .A2(net267),
    .B1(net216),
    .B2(net414),
    .C1(net295),
    .X(_06092_));
 sky130_fd_sc_hd__o21a_1 _12950_ (.A1(net110),
    .A2(net195),
    .B1(net417),
    .X(_00091_));
 sky130_fd_sc_hd__o221a_1 _12951_ (.A1(net414),
    .A2(net268),
    .B1(net216),
    .B2(net386),
    .C1(net295),
    .X(_06093_));
 sky130_fd_sc_hd__o21a_1 _12952_ (.A1(_00256_),
    .A2(net195),
    .B1(net415),
    .X(_00092_));
 sky130_fd_sc_hd__o221a_1 _12953_ (.A1(net386),
    .A2(net267),
    .B1(net216),
    .B2(\div_shifter[27] ),
    .C1(net295),
    .X(_06095_));
 sky130_fd_sc_hd__o21a_1 _12954_ (.A1(net113),
    .A2(net195),
    .B1(net387),
    .X(_00093_));
 sky130_fd_sc_hd__o221a_1 _12955_ (.A1(net446),
    .A2(net268),
    .B1(net216),
    .B2(\div_shifter[28] ),
    .C1(net295),
    .X(_06096_));
 sky130_fd_sc_hd__o21a_1 _12956_ (.A1(_00333_),
    .A2(net195),
    .B1(net447),
    .X(_00094_));
 sky130_fd_sc_hd__a221o_1 _12957_ (.A1(_04384_),
    .A2(net272),
    .B1(net221),
    .B2(net364),
    .C1(rst),
    .X(_06097_));
 sky130_fd_sc_hd__a21oi_1 _12958_ (.A1(net98),
    .A2(net200),
    .B1(net365),
    .Y(_00095_));
 sky130_fd_sc_hd__a221o_1 _12959_ (.A1(net364),
    .A2(net272),
    .B1(net221),
    .B2(net368),
    .C1(rst),
    .X(_06098_));
 sky130_fd_sc_hd__a21oi_1 _12960_ (.A1(_00418_),
    .A2(net200),
    .B1(net369),
    .Y(_00096_));
 sky130_fd_sc_hd__a21oi_1 _12961_ (.A1(_04362_),
    .A2(net272),
    .B1(rst),
    .Y(_06099_));
 sky130_fd_sc_hd__o221a_1 _12962_ (.A1(net345),
    .A2(net217),
    .B1(_00728_),
    .B2(net195),
    .C1(_06099_),
    .X(_00097_));
 sky130_fd_sc_hd__nand3_1 _12963_ (.A(net345),
    .B(net343),
    .C(net1),
    .Y(_06101_));
 sky130_fd_sc_hd__a21o_1 _12964_ (.A1(net343),
    .A2(net1),
    .B1(net345),
    .X(_06102_));
 sky130_fd_sc_hd__a32o_1 _12965_ (.A1(net272),
    .A2(_06101_),
    .A3(_06102_),
    .B1(net221),
    .B2(net557),
    .X(_06103_));
 sky130_fd_sc_hd__and2_1 _12966_ (.A(net294),
    .B(net558),
    .X(_00098_));
 sky130_fd_sc_hd__xor2_1 _12967_ (.A(_05975_),
    .B(_05976_),
    .X(_06104_));
 sky130_fd_sc_hd__mux2_1 _12968_ (.A0(\div_shifter[32] ),
    .A1(_06104_),
    .S(net1),
    .X(_06105_));
 sky130_fd_sc_hd__a22o_1 _12969_ (.A1(net551),
    .A2(net221),
    .B1(_06105_),
    .B2(net272),
    .X(_06106_));
 sky130_fd_sc_hd__and2_1 _12970_ (.A(net294),
    .B(net552),
    .X(_00099_));
 sky130_fd_sc_hd__nand2b_1 _12971_ (.A_N(_05971_),
    .B(_05972_),
    .Y(_06107_));
 sky130_fd_sc_hd__xnor2_1 _12972_ (.A(_05978_),
    .B(_06107_),
    .Y(_06108_));
 sky130_fd_sc_hd__mux2_1 _12973_ (.A0(net551),
    .A1(_06108_),
    .S(net1),
    .X(_06110_));
 sky130_fd_sc_hd__a22o_1 _12974_ (.A1(net604),
    .A2(net221),
    .B1(_06110_),
    .B2(net272),
    .X(_06111_));
 sky130_fd_sc_hd__and2_1 _12975_ (.A(net293),
    .B(_06111_),
    .X(_00100_));
 sky130_fd_sc_hd__nand2b_1 _12976_ (.A_N(_05969_),
    .B(_05970_),
    .Y(_06112_));
 sky130_fd_sc_hd__xnor2_1 _12977_ (.A(_05979_),
    .B(_06112_),
    .Y(_06113_));
 sky130_fd_sc_hd__mux2_1 _12978_ (.A0(\div_shifter[34] ),
    .A1(_06113_),
    .S(net1),
    .X(_06114_));
 sky130_fd_sc_hd__a22o_1 _12979_ (.A1(net565),
    .A2(net222),
    .B1(_06114_),
    .B2(net273),
    .X(_06115_));
 sky130_fd_sc_hd__and2_1 _12980_ (.A(net293),
    .B(net566),
    .X(_00101_));
 sky130_fd_sc_hd__xnor2_1 _12981_ (.A(_05968_),
    .B(_05980_),
    .Y(_06116_));
 sky130_fd_sc_hd__mux2_1 _12982_ (.A0(net565),
    .A1(_06116_),
    .S(net1),
    .X(_06117_));
 sky130_fd_sc_hd__a22o_1 _12983_ (.A1(net602),
    .A2(net222),
    .B1(_06117_),
    .B2(net273),
    .X(_06119_));
 sky130_fd_sc_hd__and2_1 _12984_ (.A(net293),
    .B(net603),
    .X(_00102_));
 sky130_fd_sc_hd__xnor2_1 _12985_ (.A(_05964_),
    .B(_05981_),
    .Y(_06120_));
 sky130_fd_sc_hd__mux2_1 _12986_ (.A0(\div_shifter[36] ),
    .A1(_06120_),
    .S(net1),
    .X(_06121_));
 sky130_fd_sc_hd__a22o_1 _12987_ (.A1(net593),
    .A2(net222),
    .B1(_06121_),
    .B2(net273),
    .X(_06122_));
 sky130_fd_sc_hd__and2_1 _12988_ (.A(net292),
    .B(net594),
    .X(_00103_));
 sky130_fd_sc_hd__nand2b_1 _12989_ (.A_N(_05960_),
    .B(_05961_),
    .Y(_06123_));
 sky130_fd_sc_hd__xnor2_1 _12990_ (.A(_05982_),
    .B(_06123_),
    .Y(_06124_));
 sky130_fd_sc_hd__mux2_1 _12991_ (.A0(net593),
    .A1(_06124_),
    .S(net554),
    .X(_06125_));
 sky130_fd_sc_hd__a22o_1 _12992_ (.A1(net597),
    .A2(net221),
    .B1(_06125_),
    .B2(net272),
    .X(_06126_));
 sky130_fd_sc_hd__and2_1 _12993_ (.A(net296),
    .B(net598),
    .X(_00104_));
 sky130_fd_sc_hd__nand2b_1 _12994_ (.A_N(_05958_),
    .B(_05959_),
    .Y(_06128_));
 sky130_fd_sc_hd__xnor2_1 _12995_ (.A(_05983_),
    .B(_06128_),
    .Y(_06129_));
 sky130_fd_sc_hd__mux2_1 _12996_ (.A0(net597),
    .A1(_06129_),
    .S(net554),
    .X(_06130_));
 sky130_fd_sc_hd__a22o_1 _12997_ (.A1(net608),
    .A2(net221),
    .B1(_06130_),
    .B2(net272),
    .X(_06131_));
 sky130_fd_sc_hd__and2_1 _12998_ (.A(net296),
    .B(_06131_),
    .X(_00105_));
 sky130_fd_sc_hd__nand2b_1 _12999_ (.A_N(_05956_),
    .B(_05957_),
    .Y(_06132_));
 sky130_fd_sc_hd__xnor2_1 _13000_ (.A(_05984_),
    .B(_06132_),
    .Y(_06133_));
 sky130_fd_sc_hd__mux2_1 _13001_ (.A0(\div_shifter[39] ),
    .A1(_06133_),
    .S(net1),
    .X(_06134_));
 sky130_fd_sc_hd__a22o_1 _13002_ (.A1(net587),
    .A2(net221),
    .B1(_06134_),
    .B2(net273),
    .X(_06135_));
 sky130_fd_sc_hd__and2_1 _13003_ (.A(net296),
    .B(net588),
    .X(_00106_));
 sky130_fd_sc_hd__nand2b_1 _13004_ (.A_N(_05953_),
    .B(_05954_),
    .Y(_06137_));
 sky130_fd_sc_hd__xnor2_1 _13005_ (.A(_05985_),
    .B(_06137_),
    .Y(_06138_));
 sky130_fd_sc_hd__mux2_1 _13006_ (.A0(\div_shifter[40] ),
    .A1(_06138_),
    .S(net1),
    .X(_06139_));
 sky130_fd_sc_hd__a22o_1 _13007_ (.A1(net563),
    .A2(net221),
    .B1(_06139_),
    .B2(net485),
    .X(_06140_));
 sky130_fd_sc_hd__and2_1 _13008_ (.A(net296),
    .B(net564),
    .X(_00107_));
 sky130_fd_sc_hd__nand2b_1 _13009_ (.A_N(_05951_),
    .B(_05952_),
    .Y(_06141_));
 sky130_fd_sc_hd__xnor2_1 _13010_ (.A(_05986_),
    .B(_06141_),
    .Y(_06142_));
 sky130_fd_sc_hd__mux2_1 _13011_ (.A0(net563),
    .A1(_06142_),
    .S(net1),
    .X(_06143_));
 sky130_fd_sc_hd__a22o_1 _13012_ (.A1(net585),
    .A2(net221),
    .B1(_06143_),
    .B2(net273),
    .X(_06144_));
 sky130_fd_sc_hd__and2_1 _13013_ (.A(net296),
    .B(net586),
    .X(_00108_));
 sky130_fd_sc_hd__nand2b_1 _13014_ (.A_N(_05949_),
    .B(_05950_),
    .Y(_06146_));
 sky130_fd_sc_hd__xnor2_1 _13015_ (.A(_05987_),
    .B(_06146_),
    .Y(_06147_));
 sky130_fd_sc_hd__mux2_1 _13016_ (.A0(\div_shifter[42] ),
    .A1(_06147_),
    .S(net1),
    .X(_06148_));
 sky130_fd_sc_hd__a22o_1 _13017_ (.A1(net569),
    .A2(net222),
    .B1(_06148_),
    .B2(net273),
    .X(_06149_));
 sky130_fd_sc_hd__and2_1 _13018_ (.A(net292),
    .B(net570),
    .X(_00109_));
 sky130_fd_sc_hd__nand2b_1 _13019_ (.A_N(_05947_),
    .B(_05948_),
    .Y(_06150_));
 sky130_fd_sc_hd__xnor2_1 _13020_ (.A(_05989_),
    .B(_06150_),
    .Y(_06151_));
 sky130_fd_sc_hd__mux2_1 _13021_ (.A0(\div_shifter[43] ),
    .A1(_06151_),
    .S(net554),
    .X(_06152_));
 sky130_fd_sc_hd__a22o_1 _13022_ (.A1(net567),
    .A2(net222),
    .B1(_06152_),
    .B2(net273),
    .X(_06153_));
 sky130_fd_sc_hd__and2_1 _13023_ (.A(net293),
    .B(net568),
    .X(_00110_));
 sky130_fd_sc_hd__nand2b_1 _13024_ (.A_N(_05945_),
    .B(_05946_),
    .Y(_06155_));
 sky130_fd_sc_hd__xnor2_1 _13025_ (.A(_05990_),
    .B(_06155_),
    .Y(_06156_));
 sky130_fd_sc_hd__mux2_1 _13026_ (.A0(net567),
    .A1(_06156_),
    .S(net1),
    .X(_06157_));
 sky130_fd_sc_hd__a22o_1 _13027_ (.A1(net605),
    .A2(net222),
    .B1(_06157_),
    .B2(net273),
    .X(_06158_));
 sky130_fd_sc_hd__and2_1 _13028_ (.A(net292),
    .B(_06158_),
    .X(_00111_));
 sky130_fd_sc_hd__nand2b_1 _13029_ (.A_N(_05942_),
    .B(_05943_),
    .Y(_06159_));
 sky130_fd_sc_hd__xnor2_1 _13030_ (.A(_05991_),
    .B(_06159_),
    .Y(_06160_));
 sky130_fd_sc_hd__mux2_1 _13031_ (.A0(\div_shifter[45] ),
    .A1(_06160_),
    .S(net2),
    .X(_06161_));
 sky130_fd_sc_hd__a22o_1 _13032_ (.A1(net581),
    .A2(net222),
    .B1(_06161_),
    .B2(net273),
    .X(_06162_));
 sky130_fd_sc_hd__and2_1 _13033_ (.A(net290),
    .B(net582),
    .X(_00112_));
 sky130_fd_sc_hd__nand2b_1 _13034_ (.A_N(_05940_),
    .B(_05941_),
    .Y(_06164_));
 sky130_fd_sc_hd__xnor2_1 _13035_ (.A(_05992_),
    .B(_06164_),
    .Y(_06165_));
 sky130_fd_sc_hd__mux2_1 _13036_ (.A0(\div_shifter[46] ),
    .A1(_06165_),
    .S(net2),
    .X(_06166_));
 sky130_fd_sc_hd__a22o_1 _13037_ (.A1(net575),
    .A2(net220),
    .B1(_06166_),
    .B2(net271),
    .X(_06167_));
 sky130_fd_sc_hd__and2_1 _13038_ (.A(net291),
    .B(net576),
    .X(_00113_));
 sky130_fd_sc_hd__nand2b_1 _13039_ (.A_N(_05938_),
    .B(_05939_),
    .Y(_06168_));
 sky130_fd_sc_hd__xnor2_1 _13040_ (.A(_05993_),
    .B(_06168_),
    .Y(_06169_));
 sky130_fd_sc_hd__mux2_1 _13041_ (.A0(\div_shifter[47] ),
    .A1(_06169_),
    .S(net2),
    .X(_06170_));
 sky130_fd_sc_hd__a22o_1 _13042_ (.A1(net561),
    .A2(net220),
    .B1(_06170_),
    .B2(net271),
    .X(_06171_));
 sky130_fd_sc_hd__and2_1 _13043_ (.A(net291),
    .B(net562),
    .X(_00114_));
 sky130_fd_sc_hd__nand2b_1 _13044_ (.A_N(_05936_),
    .B(_05937_),
    .Y(_06173_));
 sky130_fd_sc_hd__xnor2_1 _13045_ (.A(_05994_),
    .B(_06173_),
    .Y(_06174_));
 sky130_fd_sc_hd__mux2_1 _13046_ (.A0(net561),
    .A1(_06174_),
    .S(net2),
    .X(_06175_));
 sky130_fd_sc_hd__a22o_1 _13047_ (.A1(net606),
    .A2(net220),
    .B1(_06175_),
    .B2(net271),
    .X(_06176_));
 sky130_fd_sc_hd__and2_1 _13048_ (.A(net291),
    .B(_06176_),
    .X(_00115_));
 sky130_fd_sc_hd__nand2_1 _13049_ (.A(_05935_),
    .B(_05996_),
    .Y(_06177_));
 sky130_fd_sc_hd__xnor2_1 _13050_ (.A(_05995_),
    .B(_06177_),
    .Y(_06178_));
 sky130_fd_sc_hd__mux2_1 _13051_ (.A0(\div_shifter[49] ),
    .A1(_06178_),
    .S(net2),
    .X(_06179_));
 sky130_fd_sc_hd__a22o_1 _13052_ (.A1(net595),
    .A2(net220),
    .B1(_06179_),
    .B2(net271),
    .X(_06180_));
 sky130_fd_sc_hd__and2_1 _13053_ (.A(net290),
    .B(net596),
    .X(_00116_));
 sky130_fd_sc_hd__nand2b_1 _13054_ (.A_N(_05932_),
    .B(_05934_),
    .Y(_06182_));
 sky130_fd_sc_hd__xnor2_1 _13055_ (.A(_05997_),
    .B(_06182_),
    .Y(_06183_));
 sky130_fd_sc_hd__mux2_1 _13056_ (.A0(\div_shifter[50] ),
    .A1(_06183_),
    .S(net2),
    .X(_06184_));
 sky130_fd_sc_hd__a22o_1 _13057_ (.A1(net591),
    .A2(net220),
    .B1(_06184_),
    .B2(net271),
    .X(_06185_));
 sky130_fd_sc_hd__and2_1 _13058_ (.A(net290),
    .B(net592),
    .X(_00117_));
 sky130_fd_sc_hd__xnor2_1 _13059_ (.A(_05998_),
    .B(_06001_),
    .Y(_06186_));
 sky130_fd_sc_hd__mux2_1 _13060_ (.A0(\div_shifter[51] ),
    .A1(_06186_),
    .S(net2),
    .X(_06187_));
 sky130_fd_sc_hd__a22o_1 _13061_ (.A1(net571),
    .A2(net219),
    .B1(_06187_),
    .B2(net270),
    .X(_06188_));
 sky130_fd_sc_hd__and2_1 _13062_ (.A(net289),
    .B(net572),
    .X(_00118_));
 sky130_fd_sc_hd__nand2b_1 _13063_ (.A_N(_05929_),
    .B(_05930_),
    .Y(_06190_));
 sky130_fd_sc_hd__xnor2_1 _13064_ (.A(_06002_),
    .B(_06190_),
    .Y(_06191_));
 sky130_fd_sc_hd__mux2_1 _13065_ (.A0(net571),
    .A1(_06191_),
    .S(net2),
    .X(_06192_));
 sky130_fd_sc_hd__a22o_1 _13066_ (.A1(net577),
    .A2(net219),
    .B1(_06192_),
    .B2(net270),
    .X(_06193_));
 sky130_fd_sc_hd__and2_1 _13067_ (.A(net288),
    .B(net578),
    .X(_00119_));
 sky130_fd_sc_hd__xnor2_1 _13068_ (.A(_06003_),
    .B(_06005_),
    .Y(_06194_));
 sky130_fd_sc_hd__mux2_1 _13069_ (.A0(net577),
    .A1(_06194_),
    .S(net2),
    .X(_06195_));
 sky130_fd_sc_hd__a22o_1 _13070_ (.A1(net599),
    .A2(net219),
    .B1(_06195_),
    .B2(net270),
    .X(_06196_));
 sky130_fd_sc_hd__and2_1 _13071_ (.A(net288),
    .B(_06196_),
    .X(_00120_));
 sky130_fd_sc_hd__nand2b_1 _13072_ (.A_N(_05926_),
    .B(_05927_),
    .Y(_06197_));
 sky130_fd_sc_hd__xnor2_1 _13073_ (.A(_06006_),
    .B(_06197_),
    .Y(_06199_));
 sky130_fd_sc_hd__mux2_1 _13074_ (.A0(net599),
    .A1(_06199_),
    .S(net2),
    .X(_06200_));
 sky130_fd_sc_hd__a22o_1 _13075_ (.A1(net600),
    .A2(net220),
    .B1(_06200_),
    .B2(net271),
    .X(_06201_));
 sky130_fd_sc_hd__and2_1 _13076_ (.A(net290),
    .B(_06201_),
    .X(_00121_));
 sky130_fd_sc_hd__xnor2_1 _13077_ (.A(_06007_),
    .B(_06009_),
    .Y(_06202_));
 sky130_fd_sc_hd__mux2_1 _13078_ (.A0(\div_shifter[55] ),
    .A1(_06202_),
    .S(net2),
    .X(_06203_));
 sky130_fd_sc_hd__a22o_1 _13079_ (.A1(net579),
    .A2(net220),
    .B1(_06203_),
    .B2(net271),
    .X(_06204_));
 sky130_fd_sc_hd__and2_1 _13080_ (.A(net290),
    .B(net580),
    .X(_00122_));
 sky130_fd_sc_hd__nand2b_1 _13081_ (.A_N(_05923_),
    .B(_05924_),
    .Y(_06205_));
 sky130_fd_sc_hd__xnor2_1 _13082_ (.A(_06011_),
    .B(_06205_),
    .Y(_06206_));
 sky130_fd_sc_hd__mux2_1 _13083_ (.A0(net579),
    .A1(_06206_),
    .S(net2),
    .X(_06208_));
 sky130_fd_sc_hd__a22o_1 _13084_ (.A1(net589),
    .A2(net220),
    .B1(_06208_),
    .B2(net271),
    .X(_06209_));
 sky130_fd_sc_hd__and2_1 _13085_ (.A(net291),
    .B(net590),
    .X(_00123_));
 sky130_fd_sc_hd__xnor2_1 _13086_ (.A(_05921_),
    .B(_06012_),
    .Y(_06210_));
 sky130_fd_sc_hd__mux2_1 _13087_ (.A0(\div_shifter[57] ),
    .A1(_06210_),
    .S(net2),
    .X(_06211_));
 sky130_fd_sc_hd__a22o_1 _13088_ (.A1(net573),
    .A2(net222),
    .B1(_06211_),
    .B2(net273),
    .X(_06212_));
 sky130_fd_sc_hd__and2_1 _13089_ (.A(net292),
    .B(net574),
    .X(_00124_));
 sky130_fd_sc_hd__nand2b_1 _13090_ (.A_N(_05917_),
    .B(_05918_),
    .Y(_06213_));
 sky130_fd_sc_hd__xnor2_1 _13091_ (.A(_06013_),
    .B(_06213_),
    .Y(_06214_));
 sky130_fd_sc_hd__mux2_1 _13092_ (.A0(net573),
    .A1(_06214_),
    .S(net2),
    .X(_06215_));
 sky130_fd_sc_hd__a22o_1 _13093_ (.A1(net583),
    .A2(net222),
    .B1(_06215_),
    .B2(net273),
    .X(_06217_));
 sky130_fd_sc_hd__and2_1 _13094_ (.A(net292),
    .B(net584),
    .X(_00125_));
 sky130_fd_sc_hd__xnor2_1 _13095_ (.A(_06014_),
    .B(_06016_),
    .Y(_06218_));
 sky130_fd_sc_hd__mux2_1 _13096_ (.A0(net583),
    .A1(_06218_),
    .S(net1),
    .X(_06219_));
 sky130_fd_sc_hd__a22o_1 _13097_ (.A1(net601),
    .A2(net222),
    .B1(_06219_),
    .B2(net273),
    .X(_06220_));
 sky130_fd_sc_hd__and2_1 _13098_ (.A(net292),
    .B(_06220_),
    .X(_00126_));
 sky130_fd_sc_hd__nand2b_1 _13099_ (.A_N(_05914_),
    .B(_05915_),
    .Y(_06221_));
 sky130_fd_sc_hd__xnor2_1 _13100_ (.A(_06017_),
    .B(_06221_),
    .Y(_06222_));
 sky130_fd_sc_hd__mux2_1 _13101_ (.A0(\div_shifter[60] ),
    .A1(_06222_),
    .S(net1),
    .X(_06223_));
 sky130_fd_sc_hd__a22o_1 _13102_ (.A1(net559),
    .A2(net222),
    .B1(_06223_),
    .B2(net273),
    .X(_06224_));
 sky130_fd_sc_hd__and2_1 _13103_ (.A(net292),
    .B(net560),
    .X(_00127_));
 sky130_fd_sc_hd__nand2_1 _13104_ (.A(_05913_),
    .B(_06018_),
    .Y(_06226_));
 sky130_fd_sc_hd__nor2_1 _13105_ (.A(_04351_),
    .B(net1),
    .Y(_06227_));
 sky130_fd_sc_hd__a31o_1 _13106_ (.A1(_06019_),
    .A2(net1),
    .A3(_06226_),
    .B1(_06227_),
    .X(_06228_));
 sky130_fd_sc_hd__a22o_1 _13107_ (.A1(net553),
    .A2(net222),
    .B1(_06228_),
    .B2(net273),
    .X(_06229_));
 sky130_fd_sc_hd__and2_1 _13108_ (.A(net293),
    .B(_06229_),
    .X(_00128_));
 sky130_fd_sc_hd__or3_1 _13109_ (.A(_04340_),
    .B(_06020_),
    .C(_06022_),
    .X(_06230_));
 sky130_fd_sc_hd__a32o_1 _13110_ (.A1(net609),
    .A2(net273),
    .A3(_06230_),
    .B1(net222),
    .B2(net434),
    .X(_06231_));
 sky130_fd_sc_hd__and2_1 _13111_ (.A(net293),
    .B(net435),
    .X(_00129_));
 sky130_fd_sc_hd__nand2_1 _13112_ (.A(net408),
    .B(net217),
    .Y(_06232_));
 sky130_fd_sc_hd__o211a_1 _13113_ (.A1(net408),
    .A2(net272),
    .B1(net296),
    .C1(net409),
    .X(_00130_));
 sky130_fd_sc_hd__a22o_1 _13114_ (.A1(net472),
    .A2(net221),
    .B1(_05862_),
    .B2(net272),
    .X(_06234_));
 sky130_fd_sc_hd__o211a_1 _13115_ (.A1(net472),
    .A2(net408),
    .B1(net297),
    .C1(_06234_),
    .X(_00131_));
 sky130_fd_sc_hd__a22o_1 _13116_ (.A1(net469),
    .A2(net221),
    .B1(_05863_),
    .B2(net272),
    .X(_06235_));
 sky130_fd_sc_hd__a21o_1 _13117_ (.A1(net472),
    .A2(net408),
    .B1(net469),
    .X(_06236_));
 sky130_fd_sc_hd__and3_1 _13118_ (.A(net297),
    .B(_06235_),
    .C(_06236_),
    .X(_00132_));
 sky130_fd_sc_hd__a22o_1 _13119_ (.A1(net441),
    .A2(net221),
    .B1(_05865_),
    .B2(net272),
    .X(_06237_));
 sky130_fd_sc_hd__a31o_1 _13120_ (.A1(\div_counter[2] ),
    .A2(\div_counter[1] ),
    .A3(net408),
    .B1(net441),
    .X(_06238_));
 sky130_fd_sc_hd__and3_1 _13121_ (.A(net297),
    .B(_06237_),
    .C(net442),
    .X(_00133_));
 sky130_fd_sc_hd__a22o_1 _13122_ (.A1(net331),
    .A2(net221),
    .B1(_05866_),
    .B2(net272),
    .X(_06239_));
 sky130_fd_sc_hd__o211a_1 _13123_ (.A1(net331),
    .A2(_05864_),
    .B1(_06239_),
    .C1(net297),
    .X(_00134_));
 sky130_fd_sc_hd__o21a_1 _13124_ (.A1(net467),
    .A2(_05867_),
    .B1(net297),
    .X(_00135_));
 sky130_fd_sc_hd__dfxtp_1 _13125_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00000_),
    .Q(busy_l));
 sky130_fd_sc_hd__dfxtp_1 _13126_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00001_),
    .Q(divi1_sign));
 sky130_fd_sc_hd__dfxtp_1 _13127_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(net344),
    .Q(\divi2_l[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13128_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00003_),
    .Q(\divi2_l[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13129_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00004_),
    .Q(\divi2_l[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13130_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00005_),
    .Q(\divi2_l[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13131_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00006_),
    .Q(\divi2_l[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13132_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00007_),
    .Q(\divi2_l[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13133_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00008_),
    .Q(\divi2_l[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13134_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00009_),
    .Q(\divi2_l[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13135_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net336),
    .Q(\divi2_l[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13136_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net334),
    .Q(\divi2_l[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13137_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net320),
    .Q(\divi2_l[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13138_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(net324),
    .Q(\divi2_l[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13139_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00014_),
    .Q(\divi2_l[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13140_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(net318),
    .Q(\divi2_l[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13141_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00016_),
    .Q(\divi2_l[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13142_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00017_),
    .Q(\divi2_l[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13143_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00018_),
    .Q(\divi2_l[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13144_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net314),
    .Q(\divi2_l[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13145_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net312),
    .Q(\divi2_l[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13146_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net310),
    .Q(\divi2_l[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13147_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00022_),
    .Q(\divi2_l[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13148_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(net322),
    .Q(\divi2_l[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13149_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net330),
    .Q(\divi2_l[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13150_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net326),
    .Q(\divi2_l[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13151_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net338),
    .Q(\divi2_l[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13152_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net328),
    .Q(\divi2_l[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13153_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(net340),
    .Q(\divi2_l[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13154_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00029_),
    .Q(\divi2_l[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13155_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00030_),
    .Q(\divi2_l[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13156_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00031_),
    .Q(\divi2_l[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13157_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net316),
    .Q(\divi2_l[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13158_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00033_),
    .Q(\divi2_l[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13159_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00034_),
    .Q(\div_res[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13160_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00035_),
    .Q(\div_res[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13161_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00036_),
    .Q(\div_res[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13162_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net504),
    .Q(\div_res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13163_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00038_),
    .Q(\div_res[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13164_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net532),
    .Q(\div_res[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13165_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net523),
    .Q(\div_res[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13166_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00041_),
    .Q(\div_res[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13167_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net510),
    .Q(\div_res[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13168_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(net507),
    .Q(\div_res[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13169_ (.CLK(clknet_4_0_0_wb_clk_i),
    .D(_00044_),
    .Q(\div_res[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13170_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net496),
    .Q(\div_res[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13171_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net517),
    .Q(\div_res[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13172_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00047_),
    .Q(\div_res[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13173_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00048_),
    .Q(\div_res[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13174_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net481),
    .Q(\div_res[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13175_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00050_),
    .Q(\div_res[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13176_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00051_),
    .Q(\div_res[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13177_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(net489),
    .Q(\div_res[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13178_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00053_),
    .Q(\div_res[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13179_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net478),
    .Q(\div_res[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13180_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net520),
    .Q(\div_res[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13181_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net501),
    .Q(\div_res[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13182_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00057_),
    .Q(\div_res[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13183_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00058_),
    .Q(\div_res[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13184_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(net538),
    .Q(\div_res[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13185_ (.CLK(clknet_4_1_0_wb_clk_i),
    .D(_00060_),
    .Q(\div_res[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13186_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(net535),
    .Q(\div_res[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13187_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00062_),
    .Q(\div_res[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13188_ (.CLK(clknet_4_3_0_wb_clk_i),
    .D(_00063_),
    .Q(\div_res[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13189_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net484),
    .Q(\div_res[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13190_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(net438),
    .Q(\div_res[31] ));
 sky130_fd_sc_hd__dfxtp_1 _13191_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00066_),
    .Q(\div_shifter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13192_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00067_),
    .Q(\div_shifter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13193_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net462),
    .Q(\div_shifter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13194_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(net420),
    .Q(\div_shifter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13195_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00070_),
    .Q(\div_shifter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13196_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00071_),
    .Q(\div_shifter[5] ));
 sky130_fd_sc_hd__dfxtp_1 _13197_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00072_),
    .Q(\div_shifter[6] ));
 sky130_fd_sc_hd__dfxtp_1 _13198_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00073_),
    .Q(\div_shifter[7] ));
 sky130_fd_sc_hd__dfxtp_1 _13199_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net429),
    .Q(\div_shifter[8] ));
 sky130_fd_sc_hd__dfxtp_1 _13200_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net407),
    .Q(\div_shifter[9] ));
 sky130_fd_sc_hd__dfxtp_1 _13201_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00076_),
    .Q(\div_shifter[10] ));
 sky130_fd_sc_hd__dfxtp_1 _13202_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00077_),
    .Q(\div_shifter[11] ));
 sky130_fd_sc_hd__dfxtp_1 _13203_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00078_),
    .Q(\div_shifter[12] ));
 sky130_fd_sc_hd__dfxtp_1 _13204_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net352),
    .Q(\div_shifter[13] ));
 sky130_fd_sc_hd__dfxtp_1 _13205_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net451),
    .Q(\div_shifter[14] ));
 sky130_fd_sc_hd__dfxtp_1 _13206_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(net395),
    .Q(\div_shifter[15] ));
 sky130_fd_sc_hd__dfxtp_1 _13207_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00082_),
    .Q(\div_shifter[16] ));
 sky130_fd_sc_hd__dfxtp_1 _13208_ (.CLK(clknet_4_8_0_wb_clk_i),
    .D(_00083_),
    .Q(\div_shifter[17] ));
 sky130_fd_sc_hd__dfxtp_1 _13209_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net349),
    .Q(\div_shifter[18] ));
 sky130_fd_sc_hd__dfxtp_1 _13210_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net426),
    .Q(\div_shifter[19] ));
 sky130_fd_sc_hd__dfxtp_1 _13211_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00086_),
    .Q(\div_shifter[20] ));
 sky130_fd_sc_hd__dfxtp_1 _13212_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net413),
    .Q(\div_shifter[21] ));
 sky130_fd_sc_hd__dfxtp_1 _13213_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00088_),
    .Q(\div_shifter[22] ));
 sky130_fd_sc_hd__dfxtp_1 _13214_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net423),
    .Q(\div_shifter[23] ));
 sky130_fd_sc_hd__dfxtp_1 _13215_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(net402),
    .Q(\div_shifter[24] ));
 sky130_fd_sc_hd__dfxtp_1 _13216_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00091_),
    .Q(\div_shifter[25] ));
 sky130_fd_sc_hd__dfxtp_1 _13217_ (.CLK(clknet_4_10_0_wb_clk_i),
    .D(_00092_),
    .Q(\div_shifter[26] ));
 sky130_fd_sc_hd__dfxtp_1 _13218_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net388),
    .Q(\div_shifter[27] ));
 sky130_fd_sc_hd__dfxtp_1 _13219_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net448),
    .Q(\div_shifter[28] ));
 sky130_fd_sc_hd__dfxtp_1 _13220_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net366),
    .Q(\div_shifter[29] ));
 sky130_fd_sc_hd__dfxtp_1 _13221_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(_00096_),
    .Q(\div_shifter[30] ));
 sky130_fd_sc_hd__dfxtp_1 _13222_ (.CLK(clknet_4_11_0_wb_clk_i),
    .D(net346),
    .Q(\div_shifter[31] ));
 sky130_fd_sc_hd__dfxtp_2 _13223_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00098_),
    .Q(\div_shifter[32] ));
 sky130_fd_sc_hd__dfxtp_1 _13224_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00099_),
    .Q(\div_shifter[33] ));
 sky130_fd_sc_hd__dfxtp_1 _13225_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00100_),
    .Q(\div_shifter[34] ));
 sky130_fd_sc_hd__dfxtp_1 _13226_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00101_),
    .Q(\div_shifter[35] ));
 sky130_fd_sc_hd__dfxtp_1 _13227_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00102_),
    .Q(\div_shifter[36] ));
 sky130_fd_sc_hd__dfxtp_1 _13228_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00103_),
    .Q(\div_shifter[37] ));
 sky130_fd_sc_hd__dfxtp_1 _13229_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00104_),
    .Q(\div_shifter[38] ));
 sky130_fd_sc_hd__dfxtp_1 _13230_ (.CLK(clknet_4_14_0_wb_clk_i),
    .D(_00105_),
    .Q(\div_shifter[39] ));
 sky130_fd_sc_hd__dfxtp_1 _13231_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00106_),
    .Q(\div_shifter[40] ));
 sky130_fd_sc_hd__dfxtp_1 _13232_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00107_),
    .Q(\div_shifter[41] ));
 sky130_fd_sc_hd__dfxtp_1 _13233_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(_00108_),
    .Q(\div_shifter[42] ));
 sky130_fd_sc_hd__dfxtp_1 _13234_ (.CLK(clknet_4_13_0_wb_clk_i),
    .D(_00109_),
    .Q(\div_shifter[43] ));
 sky130_fd_sc_hd__dfxtp_1 _13235_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00110_),
    .Q(\div_shifter[44] ));
 sky130_fd_sc_hd__dfxtp_1 _13236_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00111_),
    .Q(\div_shifter[45] ));
 sky130_fd_sc_hd__dfxtp_1 _13237_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00112_),
    .Q(\div_shifter[46] ));
 sky130_fd_sc_hd__dfxtp_1 _13238_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00113_),
    .Q(\div_shifter[47] ));
 sky130_fd_sc_hd__dfxtp_1 _13239_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00114_),
    .Q(\div_shifter[48] ));
 sky130_fd_sc_hd__dfxtp_1 _13240_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00115_),
    .Q(\div_shifter[49] ));
 sky130_fd_sc_hd__dfxtp_1 _13241_ (.CLK(clknet_4_6_0_wb_clk_i),
    .D(_00116_),
    .Q(\div_shifter[50] ));
 sky130_fd_sc_hd__dfxtp_1 _13242_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00117_),
    .Q(\div_shifter[51] ));
 sky130_fd_sc_hd__dfxtp_1 _13243_ (.CLK(clknet_4_4_0_wb_clk_i),
    .D(_00118_),
    .Q(\div_shifter[52] ));
 sky130_fd_sc_hd__dfxtp_1 _13244_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00119_),
    .Q(\div_shifter[53] ));
 sky130_fd_sc_hd__dfxtp_1 _13245_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00120_),
    .Q(\div_shifter[54] ));
 sky130_fd_sc_hd__dfxtp_1 _13246_ (.CLK(clknet_4_5_0_wb_clk_i),
    .D(_00121_),
    .Q(\div_shifter[55] ));
 sky130_fd_sc_hd__dfxtp_1 _13247_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00122_),
    .Q(\div_shifter[56] ));
 sky130_fd_sc_hd__dfxtp_1 _13248_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00123_),
    .Q(\div_shifter[57] ));
 sky130_fd_sc_hd__dfxtp_1 _13249_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00124_),
    .Q(\div_shifter[58] ));
 sky130_fd_sc_hd__dfxtp_1 _13250_ (.CLK(clknet_4_7_0_wb_clk_i),
    .D(_00125_),
    .Q(\div_shifter[59] ));
 sky130_fd_sc_hd__dfxtp_1 _13251_ (.CLK(clknet_4_12_0_wb_clk_i),
    .D(_00126_),
    .Q(\div_shifter[60] ));
 sky130_fd_sc_hd__dfxtp_1 _13252_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00127_),
    .Q(\div_shifter[61] ));
 sky130_fd_sc_hd__dfxtp_1 _13253_ (.CLK(clknet_4_9_0_wb_clk_i),
    .D(_00128_),
    .Q(\div_shifter[62] ));
 sky130_fd_sc_hd__dfxtp_1 _13254_ (.CLK(clknet_4_2_0_wb_clk_i),
    .D(_00129_),
    .Q(\div_shifter[63] ));
 sky130_fd_sc_hd__dfxtp_1 _13255_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net410),
    .Q(\div_counter[0] ));
 sky130_fd_sc_hd__dfxtp_1 _13256_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net473),
    .Q(\div_counter[1] ));
 sky130_fd_sc_hd__dfxtp_1 _13257_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net486),
    .Q(\div_counter[2] ));
 sky130_fd_sc_hd__dfxtp_1 _13258_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net443),
    .Q(\div_counter[3] ));
 sky130_fd_sc_hd__dfxtp_1 _13259_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net332),
    .Q(\div_counter[4] ));
 sky130_fd_sc_hd__dfxtp_1 _13260_ (.CLK(clknet_4_15_0_wb_clk_i),
    .D(net468),
    .Q(div_complete));
 sky130_fd_sc_hd__buf_12 _13261_ (.A(instruction[11]),
    .X(loadstore_dest[0]));
 sky130_fd_sc_hd__buf_12 _13262_ (.A(instruction[12]),
    .X(loadstore_dest[1]));
 sky130_fd_sc_hd__buf_12 _13263_ (.A(instruction[13]),
    .X(loadstore_dest[2]));
 sky130_fd_sc_hd__buf_12 _13264_ (.A(instruction[14]),
    .X(loadstore_dest[3]));
 sky130_fd_sc_hd__buf_12 _13265_ (.A(instruction[15]),
    .X(loadstore_dest[4]));
 sky130_fd_sc_hd__buf_12 _13266_ (.A(instruction[5]),
    .X(loadstore_size[0]));
 sky130_fd_sc_hd__buf_12 _13267_ (.A(instruction[6]),
    .X(loadstore_size[1]));
 sky130_fd_sc_hd__buf_12 _13268_ (.A(instruction[8]),
    .X(pred_idx[0]));
 sky130_fd_sc_hd__buf_12 _13269_ (.A(instruction[9]),
    .X(pred_idx[1]));
 sky130_fd_sc_hd__buf_12 _13270_ (.A(instruction[10]),
    .X(pred_idx[2]));
 sky130_fd_sc_hd__buf_12 _13271_ (.A(instruction[4]),
    .X(sign_extend));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_0_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_10_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_11_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_12_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_13_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_14_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_15_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_1_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_2_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_3_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_4_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_5_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_6_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_7_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_8_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_4_9_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 fanout1 (.A(net2),
    .X(net1));
 sky130_fd_sc_hd__buf_6 fanout10 (.A(_00408_),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_4 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__buf_8 fanout101 (.A(_00318_),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_16 fanout102 (.A(net104),
    .X(net102));
 sky130_fd_sc_hd__buf_6 fanout103 (.A(net104),
    .X(net103));
 sky130_fd_sc_hd__buf_8 fanout104 (.A(_00280_),
    .X(net104));
 sky130_fd_sc_hd__buf_8 fanout105 (.A(net107),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_8 fanout106 (.A(net107),
    .X(net106));
 sky130_fd_sc_hd__buf_8 fanout107 (.A(_00272_),
    .X(net107));
 sky130_fd_sc_hd__buf_12 fanout108 (.A(net110),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_8 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_8 fanout11 (.A(net12),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_16 fanout110 (.A(_00255_),
    .X(net110));
 sky130_fd_sc_hd__buf_8 fanout111 (.A(_00248_),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_8 fanout112 (.A(_00248_),
    .X(net112));
 sky130_fd_sc_hd__buf_8 fanout113 (.A(_00248_),
    .X(net113));
 sky130_fd_sc_hd__buf_6 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__buf_8 fanout115 (.A(_00152_),
    .X(net115));
 sky130_fd_sc_hd__buf_6 fanout116 (.A(net117),
    .X(net116));
 sky130_fd_sc_hd__buf_8 fanout117 (.A(_00150_),
    .X(net117));
 sky130_fd_sc_hd__buf_6 fanout118 (.A(net120),
    .X(net118));
 sky130_fd_sc_hd__buf_4 fanout119 (.A(net120),
    .X(net119));
 sky130_fd_sc_hd__buf_6 fanout12 (.A(_00336_),
    .X(net12));
 sky130_fd_sc_hd__buf_6 fanout120 (.A(_00145_),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_8 fanout121 (.A(net122),
    .X(net121));
 sky130_fd_sc_hd__buf_8 fanout122 (.A(_06484_),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_8 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__buf_8 fanout124 (.A(_06482_),
    .X(net124));
 sky130_fd_sc_hd__buf_8 fanout125 (.A(net127),
    .X(net125));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net127),
    .X(net126));
 sky130_fd_sc_hd__buf_6 fanout127 (.A(_06481_),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_8 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__buf_6 fanout129 (.A(_06468_),
    .X(net129));
 sky130_fd_sc_hd__buf_8 fanout13 (.A(_00306_),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_8 fanout130 (.A(net131),
    .X(net130));
 sky130_fd_sc_hd__buf_8 fanout131 (.A(_06460_),
    .X(net131));
 sky130_fd_sc_hd__buf_8 fanout132 (.A(net134),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_8 fanout134 (.A(_00443_),
    .X(net134));
 sky130_fd_sc_hd__buf_12 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__buf_12 fanout136 (.A(_00435_),
    .X(net136));
 sky130_fd_sc_hd__buf_6 fanout137 (.A(net138),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_16 fanout138 (.A(net139),
    .X(net138));
 sky130_fd_sc_hd__buf_8 fanout139 (.A(_00385_),
    .X(net139));
 sky130_fd_sc_hd__buf_8 fanout14 (.A(net15),
    .X(net14));
 sky130_fd_sc_hd__buf_6 fanout140 (.A(net141),
    .X(net140));
 sky130_fd_sc_hd__buf_8 fanout141 (.A(_00311_),
    .X(net141));
 sky130_fd_sc_hd__buf_6 fanout142 (.A(net143),
    .X(net142));
 sky130_fd_sc_hd__buf_8 fanout143 (.A(_00299_),
    .X(net143));
 sky130_fd_sc_hd__buf_8 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__buf_8 fanout145 (.A(_00290_),
    .X(net145));
 sky130_fd_sc_hd__buf_6 fanout146 (.A(_00275_),
    .X(net146));
 sky130_fd_sc_hd__buf_6 fanout147 (.A(_00275_),
    .X(net147));
 sky130_fd_sc_hd__buf_6 fanout148 (.A(net149),
    .X(net148));
 sky130_fd_sc_hd__buf_8 fanout149 (.A(_00264_),
    .X(net149));
 sky130_fd_sc_hd__buf_6 fanout15 (.A(_00259_),
    .X(net15));
 sky130_fd_sc_hd__buf_6 fanout150 (.A(net151),
    .X(net150));
 sky130_fd_sc_hd__buf_8 fanout151 (.A(_00137_),
    .X(net151));
 sky130_fd_sc_hd__buf_6 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__buf_8 fanout153 (.A(_06497_),
    .X(net153));
 sky130_fd_sc_hd__buf_8 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_12 fanout155 (.A(net156),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_16 fanout156 (.A(_06473_),
    .X(net156));
 sky130_fd_sc_hd__buf_8 fanout157 (.A(net159),
    .X(net157));
 sky130_fd_sc_hd__buf_4 fanout158 (.A(net159),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_16 fanout159 (.A(_06436_),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_8 fanout16 (.A(_00227_),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_8 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__buf_8 fanout161 (.A(_00423_),
    .X(net161));
 sky130_fd_sc_hd__buf_6 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__buf_8 fanout163 (.A(_00339_),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_8 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__buf_8 fanout165 (.A(_00251_),
    .X(net165));
 sky130_fd_sc_hd__buf_6 fanout166 (.A(net167),
    .X(net166));
 sky130_fd_sc_hd__buf_8 fanout167 (.A(_00209_),
    .X(net167));
 sky130_fd_sc_hd__buf_6 fanout168 (.A(net169),
    .X(net168));
 sky130_fd_sc_hd__buf_8 fanout169 (.A(_00207_),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 fanout17 (.A(_00227_),
    .X(net17));
 sky130_fd_sc_hd__buf_6 fanout170 (.A(net171),
    .X(net170));
 sky130_fd_sc_hd__buf_8 fanout171 (.A(_00194_),
    .X(net171));
 sky130_fd_sc_hd__buf_6 fanout172 (.A(net173),
    .X(net172));
 sky130_fd_sc_hd__buf_8 fanout173 (.A(_00193_),
    .X(net173));
 sky130_fd_sc_hd__buf_6 fanout174 (.A(net175),
    .X(net174));
 sky130_fd_sc_hd__buf_8 fanout175 (.A(_00168_),
    .X(net175));
 sky130_fd_sc_hd__buf_6 fanout176 (.A(_00164_),
    .X(net176));
 sky130_fd_sc_hd__buf_6 fanout177 (.A(_00164_),
    .X(net177));
 sky130_fd_sc_hd__buf_12 fanout179 (.A(net181),
    .X(net179));
 sky130_fd_sc_hd__buf_6 fanout18 (.A(_00223_),
    .X(net18));
 sky130_fd_sc_hd__buf_6 fanout180 (.A(net181),
    .X(net180));
 sky130_fd_sc_hd__buf_12 fanout181 (.A(_06438_),
    .X(net181));
 sky130_fd_sc_hd__buf_4 fanout182 (.A(_02289_),
    .X(net182));
 sky130_fd_sc_hd__buf_2 fanout183 (.A(_02289_),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_8 fanout184 (.A(net186),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_4 fanout185 (.A(net186),
    .X(net185));
 sky130_fd_sc_hd__buf_4 fanout186 (.A(_02218_),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_8 fanout187 (.A(_02217_),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_16 fanout188 (.A(net190),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_16 fanout189 (.A(net190),
    .X(net189));
 sky130_fd_sc_hd__buf_4 fanout19 (.A(net27),
    .X(net19));
 sky130_fd_sc_hd__buf_8 fanout190 (.A(_06492_),
    .X(net190));
 sky130_fd_sc_hd__buf_12 fanout191 (.A(net192),
    .X(net191));
 sky130_fd_sc_hd__buf_12 fanout192 (.A(_06489_),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_8 fanout193 (.A(_06446_),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_4 fanout194 (.A(_06446_),
    .X(net194));
 sky130_fd_sc_hd__buf_4 fanout195 (.A(net196),
    .X(net195));
 sky130_fd_sc_hd__buf_2 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__buf_4 fanout197 (.A(_05870_),
    .X(net197));
 sky130_fd_sc_hd__buf_4 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(_05869_),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_8 fanout2 (.A(_06023_),
    .X(net2));
 sky130_fd_sc_hd__buf_4 fanout20 (.A(net22),
    .X(net20));
 sky130_fd_sc_hd__buf_4 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__buf_4 fanout201 (.A(_05869_),
    .X(net201));
 sky130_fd_sc_hd__buf_4 fanout202 (.A(net203),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_4 fanout203 (.A(_02306_),
    .X(net203));
 sky130_fd_sc_hd__buf_4 fanout204 (.A(_02301_),
    .X(net204));
 sky130_fd_sc_hd__buf_4 fanout205 (.A(_02290_),
    .X(net205));
 sky130_fd_sc_hd__buf_4 fanout206 (.A(_02213_),
    .X(net206));
 sky130_fd_sc_hd__buf_12 fanout207 (.A(net208),
    .X(net207));
 sky130_fd_sc_hd__buf_12 fanout208 (.A(_00179_),
    .X(net208));
 sky130_fd_sc_hd__buf_12 fanout209 (.A(net211),
    .X(net209));
 sky130_fd_sc_hd__buf_2 fanout21 (.A(net22),
    .X(net21));
 sky130_fd_sc_hd__buf_12 fanout210 (.A(net211),
    .X(net210));
 sky130_fd_sc_hd__buf_8 fanout211 (.A(_00159_),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_8 fanout212 (.A(_06425_),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_4 fanout213 (.A(_06425_),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_8 fanout214 (.A(_06413_),
    .X(net214));
 sky130_fd_sc_hd__buf_4 fanout216 (.A(net217),
    .X(net216));
 sky130_fd_sc_hd__buf_4 fanout217 (.A(_06399_),
    .X(net217));
 sky130_fd_sc_hd__buf_4 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__buf_4 fanout219 (.A(net220),
    .X(net219));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(net27),
    .X(net22));
 sky130_fd_sc_hd__buf_4 fanout220 (.A(_06398_),
    .X(net220));
 sky130_fd_sc_hd__buf_4 fanout221 (.A(net222),
    .X(net221));
 sky130_fd_sc_hd__buf_6 fanout222 (.A(_06398_),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_8 fanout223 (.A(net226),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_8 fanout224 (.A(net225),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_8 fanout225 (.A(net226),
    .X(net225));
 sky130_fd_sc_hd__buf_8 fanout226 (.A(_06309_),
    .X(net226));
 sky130_fd_sc_hd__buf_8 fanout227 (.A(_06308_),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_8 fanout228 (.A(net229),
    .X(net228));
 sky130_fd_sc_hd__buf_4 fanout229 (.A(_06300_),
    .X(net229));
 sky130_fd_sc_hd__buf_4 fanout23 (.A(net24),
    .X(net23));
 sky130_fd_sc_hd__buf_4 fanout231 (.A(net233),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_8 fanout232 (.A(net233),
    .X(net232));
 sky130_fd_sc_hd__buf_6 fanout233 (.A(_06293_),
    .X(net233));
 sky130_fd_sc_hd__buf_4 fanout234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__buf_4 fanout235 (.A(net236),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_4 fanout236 (.A(_06287_),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_8 fanout237 (.A(_06281_),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_8 fanout238 (.A(net240),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__buf_4 fanout24 (.A(net25),
    .X(net24));
 sky130_fd_sc_hd__buf_4 fanout240 (.A(_06280_),
    .X(net240));
 sky130_fd_sc_hd__buf_4 fanout241 (.A(net242),
    .X(net241));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(_06271_),
    .X(net242));
 sky130_fd_sc_hd__buf_8 fanout243 (.A(_04719_),
    .X(net243));
 sky130_fd_sc_hd__buf_4 fanout244 (.A(_02494_),
    .X(net244));
 sky130_fd_sc_hd__buf_2 fanout245 (.A(_02494_),
    .X(net245));
 sky130_fd_sc_hd__buf_4 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__buf_4 fanout247 (.A(_02494_),
    .X(net247));
 sky130_fd_sc_hd__buf_4 fanout248 (.A(_02304_),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 fanout249 (.A(_02304_),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_4 fanout25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_8 fanout250 (.A(_02299_),
    .X(net250));
 sky130_fd_sc_hd__buf_4 fanout251 (.A(_02292_),
    .X(net251));
 sky130_fd_sc_hd__buf_6 fanout252 (.A(net253),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_8 fanout253 (.A(_00216_),
    .X(net253));
 sky130_fd_sc_hd__buf_12 fanout254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__buf_12 fanout255 (.A(_00188_),
    .X(net255));
 sky130_fd_sc_hd__buf_8 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__buf_4 fanout258 (.A(_06391_),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_8 fanout259 (.A(net261),
    .X(net259));
 sky130_fd_sc_hd__buf_4 fanout26 (.A(net27),
    .X(net26));
 sky130_fd_sc_hd__buf_4 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_16 fanout261 (.A(_06391_),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_16 fanout262 (.A(_06390_),
    .X(net262));
 sky130_fd_sc_hd__buf_4 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_4 fanout264 (.A(_06270_),
    .X(net264));
 sky130_fd_sc_hd__buf_6 fanout265 (.A(net266),
    .X(net265));
 sky130_fd_sc_hd__buf_4 fanout266 (.A(_04698_),
    .X(net266));
 sky130_fd_sc_hd__buf_4 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__buf_4 fanout268 (.A(_04395_),
    .X(net268));
 sky130_fd_sc_hd__buf_4 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_4 fanout27 (.A(_02136_),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout270 (.A(net271),
    .X(net270));
 sky130_fd_sc_hd__buf_4 fanout271 (.A(net485),
    .X(net271));
 sky130_fd_sc_hd__buf_4 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__clkbuf_8 fanout273 (.A(net485),
    .X(net273));
 sky130_fd_sc_hd__buf_4 fanout274 (.A(net275),
    .X(net274));
 sky130_fd_sc_hd__buf_4 fanout275 (.A(_06429_),
    .X(net275));
 sky130_fd_sc_hd__buf_8 fanout276 (.A(net277),
    .X(net276));
 sky130_fd_sc_hd__buf_4 fanout277 (.A(net280),
    .X(net277));
 sky130_fd_sc_hd__buf_6 fanout278 (.A(net280),
    .X(net278));
 sky130_fd_sc_hd__buf_6 fanout279 (.A(net280),
    .X(net279));
 sky130_fd_sc_hd__clkbuf_8 fanout28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__buf_6 fanout280 (.A(_04621_),
    .X(net280));
 sky130_fd_sc_hd__buf_4 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__buf_4 fanout282 (.A(_04611_),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_4 fanout283 (.A(net284),
    .X(net283));
 sky130_fd_sc_hd__buf_6 fanout284 (.A(net285),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_8 fanout285 (.A(_04589_),
    .X(net285));
 sky130_fd_sc_hd__buf_6 fanout286 (.A(net287),
    .X(net286));
 sky130_fd_sc_hd__buf_4 fanout287 (.A(_04578_),
    .X(net287));
 sky130_fd_sc_hd__clkbuf_4 fanout288 (.A(net298),
    .X(net288));
 sky130_fd_sc_hd__buf_2 fanout289 (.A(net298),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_4 fanout29 (.A(net32),
    .X(net29));
 sky130_fd_sc_hd__buf_4 fanout290 (.A(net291),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_4 fanout291 (.A(net298),
    .X(net291));
 sky130_fd_sc_hd__buf_4 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_4 fanout293 (.A(net298),
    .X(net293));
 sky130_fd_sc_hd__buf_4 fanout294 (.A(net298),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_4 fanout295 (.A(net298),
    .X(net295));
 sky130_fd_sc_hd__buf_4 fanout296 (.A(net298),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_4 fanout298 (.A(_04525_),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_8 fanout299 (.A(net300),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_8 fanout3 (.A(net4),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_8 fanout30 (.A(net32),
    .X(net30));
 sky130_fd_sc_hd__buf_4 fanout300 (.A(_04504_),
    .X(net300));
 sky130_fd_sc_hd__buf_6 fanout301 (.A(net302),
    .X(net301));
 sky130_fd_sc_hd__buf_8 fanout302 (.A(_04416_),
    .X(net302));
 sky130_fd_sc_hd__buf_8 fanout303 (.A(reg1_val[13]),
    .X(net303));
 sky130_fd_sc_hd__buf_8 fanout304 (.A(reg1_val[0]),
    .X(net304));
 sky130_fd_sc_hd__buf_4 fanout305 (.A(instruction[7]),
    .X(net305));
 sky130_fd_sc_hd__buf_4 fanout306 (.A(instruction[7]),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_8 fanout307 (.A(instruction[7]),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_8 fanout308 (.A(instruction[2]),
    .X(net308));
 sky130_fd_sc_hd__buf_8 fanout31 (.A(net32),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_8 fanout32 (.A(_00729_),
    .X(net32));
 sky130_fd_sc_hd__buf_8 fanout33 (.A(_00728_),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_8 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__buf_8 fanout35 (.A(_00458_),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_8 fanout36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__buf_8 fanout37 (.A(_00455_),
    .X(net37));
 sky130_fd_sc_hd__buf_6 fanout38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__buf_8 fanout39 (.A(_00444_),
    .X(net39));
 sky130_fd_sc_hd__buf_6 fanout4 (.A(_00757_),
    .X(net4));
 sky130_fd_sc_hd__buf_6 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__buf_8 fanout41 (.A(_00440_),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_8 fanout42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__buf_8 fanout43 (.A(_00389_),
    .X(net43));
 sky130_fd_sc_hd__buf_6 fanout44 (.A(net46),
    .X(net44));
 sky130_fd_sc_hd__buf_4 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__buf_4 fanout46 (.A(_00340_),
    .X(net46));
 sky130_fd_sc_hd__buf_6 fanout47 (.A(_00309_),
    .X(net47));
 sky130_fd_sc_hd__buf_6 fanout48 (.A(net49),
    .X(net48));
 sky130_fd_sc_hd__buf_8 fanout49 (.A(_00291_),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_8 fanout5 (.A(net6),
    .X(net5));
 sky130_fd_sc_hd__buf_6 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__buf_8 fanout51 (.A(_00288_),
    .X(net51));
 sky130_fd_sc_hd__buf_6 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__buf_6 fanout53 (.A(_00265_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_8 fanout54 (.A(net56),
    .X(net54));
 sky130_fd_sc_hd__buf_4 fanout55 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__buf_4 fanout56 (.A(_00212_),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_8 fanout57 (.A(net59),
    .X(net57));
 sky130_fd_sc_hd__buf_4 fanout58 (.A(net59),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_8 fanout59 (.A(_00202_),
    .X(net59));
 sky130_fd_sc_hd__buf_8 fanout6 (.A(_00730_),
    .X(net6));
 sky130_fd_sc_hd__buf_6 fanout60 (.A(net61),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_8 fanout61 (.A(_00196_),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_8 fanout62 (.A(_00185_),
    .X(net62));
 sky130_fd_sc_hd__buf_4 fanout63 (.A(_00185_),
    .X(net63));
 sky130_fd_sc_hd__buf_6 fanout64 (.A(net66),
    .X(net64));
 sky130_fd_sc_hd__buf_4 fanout65 (.A(net66),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_8 fanout66 (.A(_00170_),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_8 fanout67 (.A(net69),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 fanout68 (.A(net69),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_8 fanout69 (.A(_00167_),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_8 fanout7 (.A(net8),
    .X(net7));
 sky130_fd_sc_hd__buf_6 fanout70 (.A(net72),
    .X(net70));
 sky130_fd_sc_hd__buf_4 fanout71 (.A(net72),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_8 fanout72 (.A(_00155_),
    .X(net72));
 sky130_fd_sc_hd__buf_6 fanout73 (.A(net75),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_4 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_8 fanout75 (.A(_00140_),
    .X(net75));
 sky130_fd_sc_hd__buf_6 fanout76 (.A(net77),
    .X(net76));
 sky130_fd_sc_hd__buf_8 fanout77 (.A(_00136_),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_8 fanout78 (.A(net79),
    .X(net78));
 sky130_fd_sc_hd__buf_8 fanout79 (.A(_06478_),
    .X(net79));
 sky130_fd_sc_hd__buf_6 fanout8 (.A(_00421_),
    .X(net8));
 sky130_fd_sc_hd__buf_6 fanout80 (.A(net81),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_8 fanout81 (.A(_06458_),
    .X(net81));
 sky130_fd_sc_hd__buf_6 fanout82 (.A(net83),
    .X(net82));
 sky130_fd_sc_hd__buf_6 fanout83 (.A(_06444_),
    .X(net83));
 sky130_fd_sc_hd__buf_4 fanout84 (.A(_02137_),
    .X(net84));
 sky130_fd_sc_hd__buf_4 fanout85 (.A(net86),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_4 fanout86 (.A(_02137_),
    .X(net86));
 sky130_fd_sc_hd__buf_8 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_16 fanout88 (.A(_00457_),
    .X(net88));
 sky130_fd_sc_hd__buf_8 fanout89 (.A(net91),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_8 fanout9 (.A(net10),
    .X(net9));
 sky130_fd_sc_hd__buf_4 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__buf_8 fanout91 (.A(_00449_),
    .X(net91));
 sky130_fd_sc_hd__buf_6 fanout92 (.A(net93),
    .X(net92));
 sky130_fd_sc_hd__buf_8 fanout93 (.A(_00431_),
    .X(net93));
 sky130_fd_sc_hd__buf_6 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__buf_8 fanout95 (.A(_00391_),
    .X(net95));
 sky130_fd_sc_hd__buf_8 fanout96 (.A(net98),
    .X(net96));
 sky130_fd_sc_hd__buf_8 fanout97 (.A(net98),
    .X(net97));
 sky130_fd_sc_hd__buf_8 fanout98 (.A(_00331_),
    .X(net98));
 sky130_fd_sc_hd__buf_6 fanout99 (.A(net101),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\divi2_l[19] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(_00015_),
    .X(net318));
 sky130_fd_sc_hd__clkbuf_2 hold100 (.A(\div_counter[0] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(_06232_),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(_00130_),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\div_shifter[21] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(_06087_),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(_00087_),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net416),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(_06093_),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\div_shifter[25] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_06092_),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\divi2_l[10] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\div_shifter[3] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(_06066_),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(_00069_),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\div_shifter[23] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(_06090_),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(_00089_),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\div_shifter[19] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(_06085_),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(_00085_),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\div_shifter[7] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_00012_),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(_06072_),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(_00074_),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\div_shifter[22] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(_06089_),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\div_shifter[1] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(_06063_),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\div_shifter[63] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(_06231_),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\div_res[31] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(_06061_),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\divi2_l[21] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_00065_),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\div_shifter[4] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(_06067_),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\div_counter[3] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(_06238_),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(_00133_),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\div_shifter[11] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(_06077_),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\div_shifter[27] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(_06096_),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_00023_),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(_00094_),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\div_shifter[14] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_06079_),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(_00080_),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(net456),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(_06071_),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\div_shifter[5] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(_06068_),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\div_shifter[6] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_06069_),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\divi2_l[11] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\div_shifter[10] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(_06075_),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\div_shifter[2] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(_06065_),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(_00068_),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\div_shifter[20] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(_06086_),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\div_shifter[9] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(_06074_),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(div_complete),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_00013_),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(_00135_),
    .X(net468));
 sky130_fd_sc_hd__buf_1 hold161 (.A(\div_counter[2] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(_05864_),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(_05866_),
    .X(net471));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold164 (.A(\div_counter[1] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(_00131_),
    .X(net473));
 sky130_fd_sc_hd__buf_1 hold166 (.A(\divi2_l[20] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(_05896_),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\div_res[19] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(_06048_),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\divi2_l[23] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(_00054_),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\div_res[14] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(_06042_),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(_00049_),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\div_res[29] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(_06060_),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(_00064_),
    .X(net484));
 sky130_fd_sc_hd__buf_2 hold177 (.A(busy_l),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(_00132_),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\div_res[17] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_00025_),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(_06045_),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(_00052_),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\div_res[18] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(_06047_),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\div_res[16] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(_06044_),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(net511),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(_06037_),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(_00045_),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\div_res[0] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\divi2_l[25] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(_06025_),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\div_res[22] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(_06050_),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(_00056_),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\div_res[3] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(_06027_),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(_00037_),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\div_res[9] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(_06035_),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(_00043_),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_00021_),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(_00027_),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\div_res[8] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(_06033_),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(_00042_),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\div_res[10] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(_06036_),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(net524),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(_06041_),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\div_res[12] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(_06038_),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(_00046_),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\divi2_l[22] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\div_res[20] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(_06049_),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(_00055_),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\div_res[6] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(_06031_),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(_00040_),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\div_res[13] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(_06039_),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\div_res[15] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(_06043_),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_00024_),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\div_res[23] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(_06051_),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\div_res[5] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(_06030_),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_00039_),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(net545),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(_06056_),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(_00061_),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\div_res[25] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(_06054_),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\div_counter[4] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(_00059_),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\div_res[24] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(_06053_),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\div_res[28] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(_06059_),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\div_res[26] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_06055_),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\div_res[27] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(_06057_),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\div_res[4] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_00134_),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(_06029_),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\div_res[7] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(_06032_),
    .X(net550));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold243 (.A(\div_shifter[33] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(_06106_),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\div_shifter[62] ),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_2 hold246 (.A(_06023_),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\div_res[2] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(_06026_),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\div_shifter[32] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\divi2_l[9] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(_06103_),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\div_shifter[61] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(_06224_),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\div_shifter[48] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(_06171_),
    .X(net562));
 sky130_fd_sc_hd__buf_1 hold255 (.A(\div_shifter[41] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(_06140_),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\div_shifter[35] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(_06115_),
    .X(net566));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold259 (.A(\div_shifter[44] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(_00011_),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(_06153_),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\div_shifter[43] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(_06149_),
    .X(net570));
 sky130_fd_sc_hd__buf_1 hold263 (.A(\div_shifter[52] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(_06188_),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\div_shifter[58] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(_06212_),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\div_shifter[47] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(_06167_),
    .X(net576));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold269 (.A(\div_shifter[53] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\divi2_l[8] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(_06193_),
    .X(net578));
 sky130_fd_sc_hd__buf_1 hold271 (.A(\div_shifter[56] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(_06204_),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\div_shifter[46] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(_06162_),
    .X(net582));
 sky130_fd_sc_hd__buf_1 hold275 (.A(net610),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(_06217_),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\div_shifter[42] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(_06144_),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\div_shifter[40] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_00010_),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_06135_),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\div_shifter[57] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(_06209_),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\div_shifter[51] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(_06185_),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\div_shifter[37] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_06122_),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\div_shifter[50] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(_06180_),
    .X(net596));
 sky130_fd_sc_hd__buf_1 hold289 (.A(\div_shifter[38] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\divi2_l[24] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(_06126_),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\div_shifter[54] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\div_shifter[55] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\div_shifter[60] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\div_shifter[36] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(_06119_),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\div_shifter[34] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\div_shifter[45] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\div_shifter[49] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\div_shifter[57] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\divi2_l[18] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_00026_),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\div_shifter[39] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\div_shifter[62] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\div_shifter[59] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\divi2_l[26] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_00028_),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(divi1_sign),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(_05871_),
    .X(net342));
 sky130_fd_sc_hd__buf_1 hold35 (.A(\divi2_l[0] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_00002_),
    .X(net344));
 sky130_fd_sc_hd__buf_1 hold37 (.A(\div_shifter[31] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_00097_),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\div_shifter[17] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_00020_),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_06084_),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(_00084_),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\div_shifter[12] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(_06078_),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(_00079_),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\divi2_l[4] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_05877_),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\divi2_l[15] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_05890_),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\divi2_l[28] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\divi2_l[17] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(_05906_),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\divi2_l[5] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(_05878_),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\divi2_l[1] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_05873_),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\div_shifter[29] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(_04373_),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_06097_),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(_00095_),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\div_shifter[30] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_00019_),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_04362_),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(_06098_),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\divi2_l[14] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_05889_),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\divi2_l[31] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(_05909_),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\divi2_l[16] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(_05891_),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\divi2_l[6] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_05879_),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\divi2_l[30] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\divi2_l[12] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(_05886_),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\divi2_l[3] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_05876_),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\divi2_l[7] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_05880_),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\divi2_l[2] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(_05874_),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\div_shifter[26] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(_06095_),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_00032_),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(_00093_),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\divi2_l[29] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_05907_),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net396),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_06083_),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\div_shifter[15] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_06080_),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_00081_),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\div_shifter[16] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(_06081_),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\divi2_l[13] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\div_shifter[0] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(_06062_),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\div_shifter[24] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_06091_),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(_00090_),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\divi2_l[27] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_05904_),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net465),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(_06073_),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(_00075_),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_2 max_cap178 (.A(_06463_),
    .X(net178));
 sky130_fd_sc_hd__buf_4 max_cap215 (.A(_06412_),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_8 max_cap230 (.A(_06299_),
    .X(net230));
 sky130_fd_sc_hd__buf_4 max_cap256 (.A(_00187_),
    .X(net256));
endmodule

